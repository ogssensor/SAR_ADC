VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO power_ring
  CLASS BLOCK ;
  FOREIGN power_ring ;
  ORIGIN 0.000 0.000 ;
  SIZE 122.000 BY 105.000 ;
  OBS
      LAYER met3 ;
        RECT 0.000 103.000 122.000 105.000 ;
        RECT 4.000 99.000 118.000 101.000 ;
        RECT 4.000 4.000 118.000 6.000 ;
        RECT 0.000 0.000 122.000 2.000 ;
      LAYER via3 ;
        RECT 0.200 104.400 0.600 104.800 ;
        RECT 0.800 104.400 1.200 104.800 ;
        RECT 1.400 104.400 1.800 104.800 ;
        RECT 18.200 104.400 18.600 104.800 ;
        RECT 18.800 104.400 19.200 104.800 ;
        RECT 19.400 104.400 19.800 104.800 ;
        RECT 46.200 104.400 46.600 104.800 ;
        RECT 46.800 104.400 47.200 104.800 ;
        RECT 47.400 104.400 47.800 104.800 ;
        RECT 74.200 104.400 74.600 104.800 ;
        RECT 74.800 104.400 75.200 104.800 ;
        RECT 75.400 104.400 75.800 104.800 ;
        RECT 102.200 104.400 102.600 104.800 ;
        RECT 102.800 104.400 103.200 104.800 ;
        RECT 103.400 104.400 103.800 104.800 ;
        RECT 120.200 104.400 120.600 104.800 ;
        RECT 120.800 104.400 121.200 104.800 ;
        RECT 121.400 104.400 121.800 104.800 ;
        RECT 0.200 103.800 0.600 104.200 ;
        RECT 0.800 103.800 1.200 104.200 ;
        RECT 1.400 103.800 1.800 104.200 ;
        RECT 18.200 103.800 18.600 104.200 ;
        RECT 18.800 103.800 19.200 104.200 ;
        RECT 19.400 103.800 19.800 104.200 ;
        RECT 46.200 103.800 46.600 104.200 ;
        RECT 46.800 103.800 47.200 104.200 ;
        RECT 47.400 103.800 47.800 104.200 ;
        RECT 74.200 103.800 74.600 104.200 ;
        RECT 74.800 103.800 75.200 104.200 ;
        RECT 75.400 103.800 75.800 104.200 ;
        RECT 102.200 103.800 102.600 104.200 ;
        RECT 102.800 103.800 103.200 104.200 ;
        RECT 103.400 103.800 103.800 104.200 ;
        RECT 120.200 103.800 120.600 104.200 ;
        RECT 120.800 103.800 121.200 104.200 ;
        RECT 121.400 103.800 121.800 104.200 ;
        RECT 0.200 103.200 0.600 103.600 ;
        RECT 0.800 103.200 1.200 103.600 ;
        RECT 1.400 103.200 1.800 103.600 ;
        RECT 18.200 103.200 18.600 103.600 ;
        RECT 18.800 103.200 19.200 103.600 ;
        RECT 19.400 103.200 19.800 103.600 ;
        RECT 46.200 103.200 46.600 103.600 ;
        RECT 46.800 103.200 47.200 103.600 ;
        RECT 47.400 103.200 47.800 103.600 ;
        RECT 74.200 103.200 74.600 103.600 ;
        RECT 74.800 103.200 75.200 103.600 ;
        RECT 75.400 103.200 75.800 103.600 ;
        RECT 102.200 103.200 102.600 103.600 ;
        RECT 102.800 103.200 103.200 103.600 ;
        RECT 103.400 103.200 103.800 103.600 ;
        RECT 120.200 103.200 120.600 103.600 ;
        RECT 120.800 103.200 121.200 103.600 ;
        RECT 121.400 103.200 121.800 103.600 ;
        RECT 4.200 100.400 4.600 100.800 ;
        RECT 4.800 100.400 5.200 100.800 ;
        RECT 5.400 100.400 5.800 100.800 ;
        RECT 32.200 100.400 32.600 100.800 ;
        RECT 32.800 100.400 33.200 100.800 ;
        RECT 33.400 100.400 33.800 100.800 ;
        RECT 60.200 100.400 60.600 100.800 ;
        RECT 60.800 100.400 61.200 100.800 ;
        RECT 61.400 100.400 61.800 100.800 ;
        RECT 88.200 100.400 88.600 100.800 ;
        RECT 88.800 100.400 89.200 100.800 ;
        RECT 89.400 100.400 89.800 100.800 ;
        RECT 116.200 100.400 116.600 100.800 ;
        RECT 116.800 100.400 117.200 100.800 ;
        RECT 117.400 100.400 117.800 100.800 ;
        RECT 4.200 99.800 4.600 100.200 ;
        RECT 4.800 99.800 5.200 100.200 ;
        RECT 5.400 99.800 5.800 100.200 ;
        RECT 32.200 99.800 32.600 100.200 ;
        RECT 32.800 99.800 33.200 100.200 ;
        RECT 33.400 99.800 33.800 100.200 ;
        RECT 60.200 99.800 60.600 100.200 ;
        RECT 60.800 99.800 61.200 100.200 ;
        RECT 61.400 99.800 61.800 100.200 ;
        RECT 88.200 99.800 88.600 100.200 ;
        RECT 88.800 99.800 89.200 100.200 ;
        RECT 89.400 99.800 89.800 100.200 ;
        RECT 116.200 99.800 116.600 100.200 ;
        RECT 116.800 99.800 117.200 100.200 ;
        RECT 117.400 99.800 117.800 100.200 ;
        RECT 4.200 99.200 4.600 99.600 ;
        RECT 4.800 99.200 5.200 99.600 ;
        RECT 5.400 99.200 5.800 99.600 ;
        RECT 32.200 99.200 32.600 99.600 ;
        RECT 32.800 99.200 33.200 99.600 ;
        RECT 33.400 99.200 33.800 99.600 ;
        RECT 60.200 99.200 60.600 99.600 ;
        RECT 60.800 99.200 61.200 99.600 ;
        RECT 61.400 99.200 61.800 99.600 ;
        RECT 88.200 99.200 88.600 99.600 ;
        RECT 88.800 99.200 89.200 99.600 ;
        RECT 89.400 99.200 89.800 99.600 ;
        RECT 116.200 99.200 116.600 99.600 ;
        RECT 116.800 99.200 117.200 99.600 ;
        RECT 117.400 99.200 117.800 99.600 ;
        RECT 4.200 5.400 4.600 5.800 ;
        RECT 4.800 5.400 5.200 5.800 ;
        RECT 5.400 5.400 5.800 5.800 ;
        RECT 32.200 5.400 32.600 5.800 ;
        RECT 32.800 5.400 33.200 5.800 ;
        RECT 33.400 5.400 33.800 5.800 ;
        RECT 60.200 5.400 60.600 5.800 ;
        RECT 60.800 5.400 61.200 5.800 ;
        RECT 61.400 5.400 61.800 5.800 ;
        RECT 88.200 5.400 88.600 5.800 ;
        RECT 88.800 5.400 89.200 5.800 ;
        RECT 89.400 5.400 89.800 5.800 ;
        RECT 116.200 5.400 116.600 5.800 ;
        RECT 116.800 5.400 117.200 5.800 ;
        RECT 117.400 5.400 117.800 5.800 ;
        RECT 4.200 4.800 4.600 5.200 ;
        RECT 4.800 4.800 5.200 5.200 ;
        RECT 5.400 4.800 5.800 5.200 ;
        RECT 32.200 4.800 32.600 5.200 ;
        RECT 32.800 4.800 33.200 5.200 ;
        RECT 33.400 4.800 33.800 5.200 ;
        RECT 60.200 4.800 60.600 5.200 ;
        RECT 60.800 4.800 61.200 5.200 ;
        RECT 61.400 4.800 61.800 5.200 ;
        RECT 88.200 4.800 88.600 5.200 ;
        RECT 88.800 4.800 89.200 5.200 ;
        RECT 89.400 4.800 89.800 5.200 ;
        RECT 116.200 4.800 116.600 5.200 ;
        RECT 116.800 4.800 117.200 5.200 ;
        RECT 117.400 4.800 117.800 5.200 ;
        RECT 4.200 4.200 4.600 4.600 ;
        RECT 4.800 4.200 5.200 4.600 ;
        RECT 5.400 4.200 5.800 4.600 ;
        RECT 32.200 4.200 32.600 4.600 ;
        RECT 32.800 4.200 33.200 4.600 ;
        RECT 33.400 4.200 33.800 4.600 ;
        RECT 60.200 4.200 60.600 4.600 ;
        RECT 60.800 4.200 61.200 4.600 ;
        RECT 61.400 4.200 61.800 4.600 ;
        RECT 88.200 4.200 88.600 4.600 ;
        RECT 88.800 4.200 89.200 4.600 ;
        RECT 89.400 4.200 89.800 4.600 ;
        RECT 116.200 4.200 116.600 4.600 ;
        RECT 116.800 4.200 117.200 4.600 ;
        RECT 117.400 4.200 117.800 4.600 ;
        RECT 0.200 1.400 0.600 1.800 ;
        RECT 0.800 1.400 1.200 1.800 ;
        RECT 1.400 1.400 1.800 1.800 ;
        RECT 18.200 1.400 18.600 1.800 ;
        RECT 18.800 1.400 19.200 1.800 ;
        RECT 19.400 1.400 19.800 1.800 ;
        RECT 46.200 1.400 46.600 1.800 ;
        RECT 46.800 1.400 47.200 1.800 ;
        RECT 47.400 1.400 47.800 1.800 ;
        RECT 74.200 1.400 74.600 1.800 ;
        RECT 74.800 1.400 75.200 1.800 ;
        RECT 75.400 1.400 75.800 1.800 ;
        RECT 102.200 1.400 102.600 1.800 ;
        RECT 102.800 1.400 103.200 1.800 ;
        RECT 103.400 1.400 103.800 1.800 ;
        RECT 120.200 1.400 120.600 1.800 ;
        RECT 120.800 1.400 121.200 1.800 ;
        RECT 121.400 1.400 121.800 1.800 ;
        RECT 0.200 0.800 0.600 1.200 ;
        RECT 0.800 0.800 1.200 1.200 ;
        RECT 1.400 0.800 1.800 1.200 ;
        RECT 18.200 0.800 18.600 1.200 ;
        RECT 18.800 0.800 19.200 1.200 ;
        RECT 19.400 0.800 19.800 1.200 ;
        RECT 46.200 0.800 46.600 1.200 ;
        RECT 46.800 0.800 47.200 1.200 ;
        RECT 47.400 0.800 47.800 1.200 ;
        RECT 74.200 0.800 74.600 1.200 ;
        RECT 74.800 0.800 75.200 1.200 ;
        RECT 75.400 0.800 75.800 1.200 ;
        RECT 102.200 0.800 102.600 1.200 ;
        RECT 102.800 0.800 103.200 1.200 ;
        RECT 103.400 0.800 103.800 1.200 ;
        RECT 120.200 0.800 120.600 1.200 ;
        RECT 120.800 0.800 121.200 1.200 ;
        RECT 121.400 0.800 121.800 1.200 ;
        RECT 0.200 0.200 0.600 0.600 ;
        RECT 0.800 0.200 1.200 0.600 ;
        RECT 1.400 0.200 1.800 0.600 ;
        RECT 18.200 0.200 18.600 0.600 ;
        RECT 18.800 0.200 19.200 0.600 ;
        RECT 19.400 0.200 19.800 0.600 ;
        RECT 46.200 0.200 46.600 0.600 ;
        RECT 46.800 0.200 47.200 0.600 ;
        RECT 47.400 0.200 47.800 0.600 ;
        RECT 74.200 0.200 74.600 0.600 ;
        RECT 74.800 0.200 75.200 0.600 ;
        RECT 75.400 0.200 75.800 0.600 ;
        RECT 102.200 0.200 102.600 0.600 ;
        RECT 102.800 0.200 103.200 0.600 ;
        RECT 103.400 0.200 103.800 0.600 ;
        RECT 120.200 0.200 120.600 0.600 ;
        RECT 120.800 0.200 121.200 0.600 ;
        RECT 121.400 0.200 121.800 0.600 ;
      LAYER met4 ;
        RECT 0.000 0.000 2.000 105.000 ;
        RECT 4.000 4.000 6.000 101.000 ;
        RECT 18.000 0.000 20.000 105.000 ;
        RECT 32.000 4.000 34.000 101.000 ;
        RECT 46.000 0.000 48.000 105.000 ;
        RECT 60.000 4.000 62.000 101.000 ;
        RECT 74.000 0.000 76.000 105.000 ;
        RECT 88.000 4.000 90.000 101.000 ;
        RECT 102.000 0.000 104.000 105.000 ;
        RECT 116.000 4.000 118.000 101.000 ;
        RECT 120.000 0.000 122.000 105.000 ;
  END
END power_ring
MACRO ring_osc
  CLASS BLOCK ;
  FOREIGN ring_osc ;
  ORIGIN 7.950 1.720 ;
  SIZE 123.550 BY 33.220 ;
  OBS
      LAYER nwell ;
        RECT -1.000 24.105 1.680 25.950 ;
        RECT 2.995 24.105 4.755 25.950 ;
        RECT 8.480 22.965 97.550 29.840 ;
        RECT 19.520 22.960 26.710 22.965 ;
        RECT 37.230 22.960 44.420 22.965 ;
        RECT 54.940 22.960 62.130 22.965 ;
        RECT 72.650 22.960 79.840 22.965 ;
        RECT 90.360 22.960 97.550 22.965 ;
      LAYER pwell ;
        RECT -0.660 22.715 -0.490 22.885 ;
        RECT 3.330 22.715 3.500 22.885 ;
        RECT 8.480 15.470 97.550 22.570 ;
        RECT 100.500 20.000 103.500 25.000 ;
        RECT 100.500 19.000 108.500 20.000 ;
        RECT 102.500 17.000 108.500 19.000 ;
        RECT 0.000 7.270 106.780 14.370 ;
      LAYER nwell ;
        RECT 0.000 6.875 7.190 6.880 ;
        RECT 17.710 6.875 24.900 6.880 ;
        RECT 35.420 6.875 42.610 6.880 ;
        RECT 53.130 6.875 60.320 6.880 ;
        RECT 70.840 6.875 78.030 6.880 ;
        RECT 88.550 6.875 95.740 6.880 ;
        RECT 0.000 0.000 106.780 6.875 ;
      LAYER li1 ;
        RECT 8.660 29.660 10.550 29.690 ;
        RECT 12.340 29.660 16.190 29.690 ;
        RECT 17.850 29.660 21.700 29.690 ;
        RECT 23.540 29.660 24.940 29.690 ;
        RECT 26.370 29.660 28.260 29.690 ;
        RECT 30.050 29.660 33.900 29.690 ;
        RECT 35.560 29.660 39.410 29.690 ;
        RECT 41.250 29.660 42.650 29.690 ;
        RECT 44.080 29.660 45.970 29.690 ;
        RECT 47.760 29.660 51.610 29.690 ;
        RECT 53.270 29.660 57.120 29.690 ;
        RECT 58.960 29.660 60.360 29.690 ;
        RECT 61.790 29.660 63.680 29.690 ;
        RECT 65.470 29.660 69.320 29.690 ;
        RECT 70.980 29.660 74.830 29.690 ;
        RECT 76.670 29.660 78.070 29.690 ;
        RECT 79.500 29.660 81.390 29.690 ;
        RECT 83.180 29.660 87.030 29.690 ;
        RECT 88.690 29.660 92.540 29.690 ;
        RECT 94.380 29.660 95.780 29.690 ;
        RECT 8.660 29.490 97.370 29.660 ;
        RECT 8.660 29.330 10.550 29.490 ;
        RECT 12.340 29.330 16.190 29.490 ;
        RECT 17.850 29.330 21.700 29.490 ;
        RECT 23.540 29.330 24.940 29.490 ;
        RECT 26.370 29.330 28.260 29.490 ;
        RECT 30.050 29.330 33.900 29.490 ;
        RECT 35.560 29.330 39.410 29.490 ;
        RECT 41.250 29.330 42.650 29.490 ;
        RECT 44.080 29.330 45.970 29.490 ;
        RECT 47.760 29.330 51.610 29.490 ;
        RECT 53.270 29.330 57.120 29.490 ;
        RECT 58.960 29.330 60.360 29.490 ;
        RECT 61.790 29.330 63.680 29.490 ;
        RECT 65.470 29.330 69.320 29.490 ;
        RECT 70.980 29.330 74.830 29.490 ;
        RECT 76.670 29.330 78.070 29.490 ;
        RECT 79.500 29.330 81.390 29.490 ;
        RECT 83.180 29.330 87.030 29.490 ;
        RECT 88.690 29.330 92.540 29.490 ;
        RECT 94.380 29.330 95.780 29.490 ;
        RECT -0.810 25.605 0.190 25.770 ;
        RECT 3.185 25.605 4.185 25.770 ;
        RECT -0.810 25.435 1.490 25.605 ;
        RECT 3.185 25.435 4.565 25.605 ;
        RECT -0.725 24.865 -0.465 25.265 ;
        RECT -0.295 25.035 0.640 25.435 ;
        RECT 0.810 24.925 1.405 25.265 ;
        RECT -0.725 24.695 0.640 24.865 ;
        RECT -0.725 24.300 -0.265 24.525 ;
        RECT -7.900 24.000 -0.265 24.300 ;
        RECT -0.725 23.795 -0.265 24.000 ;
        RECT -0.095 23.625 0.640 24.695 ;
        RECT -0.725 23.455 0.640 23.625 ;
        RECT 0.810 23.605 0.985 24.925 ;
        RECT 1.165 24.750 1.405 24.755 ;
        RECT 1.680 24.750 3.005 24.960 ;
        RECT 1.165 24.740 3.005 24.750 ;
        RECT 1.165 24.530 1.900 24.740 ;
        RECT 2.785 24.535 3.005 24.740 ;
        RECT 3.460 24.710 3.790 25.435 ;
        RECT 3.270 24.535 3.790 24.540 ;
        RECT 1.165 23.775 1.405 24.530 ;
        RECT 2.785 24.315 3.790 24.535 ;
        RECT 0.810 23.480 1.405 23.605 ;
        RECT 2.210 23.480 2.510 24.310 ;
        RECT -0.725 23.055 -0.465 23.455 ;
        RECT -0.295 22.885 0.640 23.285 ;
        RECT 0.810 23.180 2.510 23.480 ;
        RECT 0.810 23.055 1.405 23.180 ;
        RECT 3.270 23.055 3.790 24.315 ;
        RECT 3.960 23.715 4.480 25.265 ;
        RECT 8.660 24.460 8.830 29.330 ;
        RECT 9.170 24.040 9.460 29.330 ;
        RECT 3.960 22.885 4.300 23.545 ;
        RECT 10.380 22.950 10.760 23.000 ;
        RECT -0.810 22.715 1.490 22.885 ;
        RECT 3.185 22.715 4.565 22.885 ;
        RECT 9.430 22.590 10.760 22.950 ;
        RECT 10.380 22.540 10.760 22.590 ;
        RECT 9.170 16.090 9.460 21.540 ;
        RECT 11.355 16.500 11.655 29.090 ;
        RECT 13.550 24.040 13.840 29.330 ;
        RECT 14.180 24.460 14.350 29.330 ;
        RECT 14.690 24.040 14.980 29.330 ;
        RECT 12.250 22.950 12.630 23.000 ;
        RECT 15.900 22.950 16.280 23.000 ;
        RECT 12.250 22.590 13.580 22.950 ;
        RECT 14.950 22.590 16.280 22.950 ;
        RECT 12.250 22.540 12.630 22.590 ;
        RECT 15.900 22.540 16.280 22.590 ;
        RECT 13.550 16.090 13.840 21.540 ;
        RECT 14.690 16.090 14.980 21.540 ;
        RECT 16.875 16.500 17.175 29.090 ;
        RECT 19.070 24.040 19.360 29.330 ;
        RECT 19.700 24.460 19.870 29.330 ;
        RECT 20.210 24.030 20.500 29.330 ;
        RECT 17.770 22.950 18.150 23.000 ;
        RECT 21.420 22.950 21.800 23.000 ;
        RECT 17.770 22.590 19.100 22.950 ;
        RECT 20.470 22.590 21.800 22.950 ;
        RECT 17.770 22.540 18.150 22.590 ;
        RECT 21.420 22.540 21.800 22.590 ;
        RECT 19.070 16.090 19.360 21.540 ;
        RECT 20.210 16.090 20.500 21.540 ;
        RECT 22.400 16.500 22.700 29.090 ;
        RECT 23.540 24.030 23.830 29.330 ;
        RECT 24.750 22.950 25.130 23.000 ;
        RECT 23.800 22.590 25.130 22.950 ;
        RECT 24.750 22.540 25.130 22.590 ;
        RECT 23.540 16.090 23.830 21.540 ;
        RECT 25.730 16.500 26.030 29.090 ;
        RECT 26.370 24.460 26.540 29.330 ;
        RECT 26.880 24.040 27.170 29.330 ;
        RECT 28.090 22.950 28.470 23.000 ;
        RECT 27.140 22.590 28.470 22.950 ;
        RECT 28.090 22.540 28.470 22.590 ;
        RECT 26.880 16.090 27.170 21.540 ;
        RECT 29.065 16.500 29.365 29.090 ;
        RECT 31.260 24.040 31.550 29.330 ;
        RECT 31.890 24.460 32.060 29.330 ;
        RECT 32.400 24.040 32.690 29.330 ;
        RECT 29.960 22.950 30.340 23.000 ;
        RECT 33.610 22.950 33.990 23.000 ;
        RECT 29.960 22.590 31.290 22.950 ;
        RECT 32.660 22.590 33.990 22.950 ;
        RECT 29.960 22.540 30.340 22.590 ;
        RECT 33.610 22.540 33.990 22.590 ;
        RECT 31.260 16.090 31.550 21.540 ;
        RECT 32.400 16.090 32.690 21.540 ;
        RECT 34.585 16.500 34.885 29.090 ;
        RECT 36.780 24.040 37.070 29.330 ;
        RECT 37.410 24.460 37.580 29.330 ;
        RECT 37.920 24.030 38.210 29.330 ;
        RECT 35.480 22.950 35.860 23.000 ;
        RECT 39.130 22.950 39.510 23.000 ;
        RECT 35.480 22.590 36.810 22.950 ;
        RECT 38.180 22.590 39.510 22.950 ;
        RECT 35.480 22.540 35.860 22.590 ;
        RECT 39.130 22.540 39.510 22.590 ;
        RECT 36.780 16.090 37.070 21.540 ;
        RECT 37.920 16.090 38.210 21.540 ;
        RECT 40.110 16.500 40.410 29.090 ;
        RECT 41.250 24.030 41.540 29.330 ;
        RECT 42.460 22.950 42.840 23.000 ;
        RECT 41.510 22.590 42.840 22.950 ;
        RECT 42.460 22.540 42.840 22.590 ;
        RECT 41.250 16.090 41.540 21.540 ;
        RECT 43.440 16.500 43.740 29.090 ;
        RECT 44.080 24.460 44.250 29.330 ;
        RECT 44.590 24.040 44.880 29.330 ;
        RECT 45.800 22.950 46.180 23.000 ;
        RECT 44.850 22.590 46.180 22.950 ;
        RECT 45.800 22.540 46.180 22.590 ;
        RECT 44.590 16.090 44.880 21.540 ;
        RECT 46.775 16.500 47.075 29.090 ;
        RECT 48.970 24.040 49.260 29.330 ;
        RECT 49.600 24.460 49.770 29.330 ;
        RECT 50.110 24.040 50.400 29.330 ;
        RECT 47.670 22.950 48.050 23.000 ;
        RECT 51.320 22.950 51.700 23.000 ;
        RECT 47.670 22.590 49.000 22.950 ;
        RECT 50.370 22.590 51.700 22.950 ;
        RECT 47.670 22.540 48.050 22.590 ;
        RECT 51.320 22.540 51.700 22.590 ;
        RECT 48.970 16.090 49.260 21.540 ;
        RECT 50.110 16.090 50.400 21.540 ;
        RECT 52.295 16.500 52.595 29.090 ;
        RECT 54.490 24.040 54.780 29.330 ;
        RECT 55.120 24.460 55.290 29.330 ;
        RECT 55.630 24.030 55.920 29.330 ;
        RECT 53.190 22.950 53.570 23.000 ;
        RECT 56.840 22.950 57.220 23.000 ;
        RECT 53.190 22.590 54.520 22.950 ;
        RECT 55.890 22.590 57.220 22.950 ;
        RECT 53.190 22.540 53.570 22.590 ;
        RECT 56.840 22.540 57.220 22.590 ;
        RECT 54.490 16.090 54.780 21.540 ;
        RECT 55.630 16.090 55.920 21.540 ;
        RECT 57.820 16.500 58.120 29.090 ;
        RECT 58.960 24.030 59.250 29.330 ;
        RECT 60.170 22.950 60.550 23.000 ;
        RECT 59.220 22.590 60.550 22.950 ;
        RECT 60.170 22.540 60.550 22.590 ;
        RECT 58.960 16.090 59.250 21.540 ;
        RECT 61.150 16.500 61.450 29.090 ;
        RECT 61.790 24.460 61.960 29.330 ;
        RECT 62.300 24.040 62.590 29.330 ;
        RECT 63.510 22.950 63.890 23.000 ;
        RECT 62.560 22.590 63.890 22.950 ;
        RECT 63.510 22.540 63.890 22.590 ;
        RECT 62.300 16.090 62.590 21.540 ;
        RECT 64.485 16.500 64.785 29.090 ;
        RECT 66.680 24.040 66.970 29.330 ;
        RECT 67.310 24.460 67.480 29.330 ;
        RECT 67.820 24.040 68.110 29.330 ;
        RECT 65.380 22.950 65.760 23.000 ;
        RECT 69.030 22.950 69.410 23.000 ;
        RECT 65.380 22.590 66.710 22.950 ;
        RECT 68.080 22.590 69.410 22.950 ;
        RECT 65.380 22.540 65.760 22.590 ;
        RECT 69.030 22.540 69.410 22.590 ;
        RECT 66.680 16.090 66.970 21.540 ;
        RECT 67.820 16.090 68.110 21.540 ;
        RECT 70.005 16.500 70.305 29.090 ;
        RECT 72.200 24.040 72.490 29.330 ;
        RECT 72.830 24.460 73.000 29.330 ;
        RECT 73.340 24.030 73.630 29.330 ;
        RECT 70.900 22.950 71.280 23.000 ;
        RECT 74.550 22.950 74.930 23.000 ;
        RECT 70.900 22.590 72.230 22.950 ;
        RECT 73.600 22.590 74.930 22.950 ;
        RECT 70.900 22.540 71.280 22.590 ;
        RECT 74.550 22.540 74.930 22.590 ;
        RECT 72.200 16.090 72.490 21.540 ;
        RECT 73.340 16.090 73.630 21.540 ;
        RECT 75.530 16.500 75.830 29.090 ;
        RECT 76.670 24.030 76.960 29.330 ;
        RECT 77.880 22.950 78.260 23.000 ;
        RECT 76.930 22.590 78.260 22.950 ;
        RECT 77.880 22.540 78.260 22.590 ;
        RECT 76.670 16.090 76.960 21.540 ;
        RECT 78.860 16.500 79.160 29.090 ;
        RECT 79.500 24.460 79.670 29.330 ;
        RECT 80.010 24.040 80.300 29.330 ;
        RECT 81.220 22.950 81.600 23.000 ;
        RECT 80.270 22.590 81.600 22.950 ;
        RECT 81.220 22.540 81.600 22.590 ;
        RECT 80.010 16.090 80.300 21.540 ;
        RECT 82.195 16.500 82.495 29.090 ;
        RECT 84.390 24.040 84.680 29.330 ;
        RECT 85.020 24.460 85.190 29.330 ;
        RECT 85.530 24.040 85.820 29.330 ;
        RECT 83.090 22.950 83.470 23.000 ;
        RECT 86.740 22.950 87.120 23.000 ;
        RECT 83.090 22.590 84.420 22.950 ;
        RECT 85.790 22.590 87.120 22.950 ;
        RECT 83.090 22.540 83.470 22.590 ;
        RECT 86.740 22.540 87.120 22.590 ;
        RECT 84.390 16.090 84.680 21.540 ;
        RECT 85.530 16.090 85.820 21.540 ;
        RECT 87.715 16.500 88.015 29.090 ;
        RECT 89.910 24.040 90.200 29.330 ;
        RECT 90.540 24.460 90.710 29.330 ;
        RECT 91.050 24.030 91.340 29.330 ;
        RECT 88.610 22.950 88.990 23.000 ;
        RECT 92.260 22.950 92.640 23.000 ;
        RECT 88.610 22.590 89.940 22.950 ;
        RECT 91.310 22.590 92.640 22.950 ;
        RECT 88.610 22.540 88.990 22.590 ;
        RECT 92.260 22.540 92.640 22.590 ;
        RECT 89.910 16.090 90.200 21.540 ;
        RECT 91.050 16.090 91.340 21.540 ;
        RECT 93.240 16.500 93.540 29.090 ;
        RECT 94.380 24.030 94.670 29.330 ;
        RECT 95.590 22.950 95.970 23.000 ;
        RECT 94.640 22.590 95.970 22.950 ;
        RECT 95.590 22.540 95.970 22.590 ;
        RECT 94.380 16.090 94.670 21.540 ;
        RECT 96.570 16.500 96.870 29.090 ;
        RECT 101.000 24.015 103.000 24.380 ;
        RECT 101.000 19.500 103.000 19.865 ;
        RECT 102.000 18.500 103.365 19.500 ;
        RECT 103.000 17.500 103.365 18.500 ;
        RECT 107.515 18.500 108.500 19.500 ;
        RECT 107.515 17.500 107.880 18.500 ;
        RECT 8.660 15.730 10.550 16.090 ;
        RECT 12.340 15.730 16.190 16.090 ;
        RECT 17.850 15.730 21.700 16.090 ;
        RECT 23.540 15.730 24.940 16.090 ;
        RECT 26.370 15.730 28.260 16.090 ;
        RECT 30.050 15.730 33.900 16.090 ;
        RECT 35.560 15.730 39.410 16.090 ;
        RECT 41.250 15.730 42.650 16.090 ;
        RECT 44.080 15.730 45.970 16.090 ;
        RECT 47.760 15.730 51.610 16.090 ;
        RECT 53.270 15.730 57.120 16.090 ;
        RECT 58.960 15.730 60.360 16.090 ;
        RECT 61.790 15.730 63.680 16.090 ;
        RECT 65.470 15.730 69.320 16.090 ;
        RECT 70.980 15.730 74.830 16.090 ;
        RECT 76.670 15.730 78.070 16.090 ;
        RECT 79.500 15.730 81.390 16.090 ;
        RECT 83.180 15.730 87.030 16.090 ;
        RECT 88.690 15.730 92.540 16.090 ;
        RECT 94.380 15.730 95.780 16.090 ;
        RECT 1.770 13.750 3.170 14.110 ;
        RECT 5.010 13.750 8.860 14.110 ;
        RECT 10.520 13.750 14.370 14.110 ;
        RECT 16.160 13.750 18.050 14.110 ;
        RECT 19.480 13.750 20.880 14.110 ;
        RECT 22.720 13.750 26.570 14.110 ;
        RECT 28.230 13.750 32.080 14.110 ;
        RECT 33.870 13.750 35.760 14.110 ;
        RECT 37.190 13.750 38.590 14.110 ;
        RECT 40.430 13.750 44.280 14.110 ;
        RECT 45.940 13.750 49.790 14.110 ;
        RECT 51.580 13.750 53.470 14.110 ;
        RECT 54.900 13.750 56.300 14.110 ;
        RECT 58.140 13.750 61.990 14.110 ;
        RECT 63.650 13.750 67.500 14.110 ;
        RECT 69.290 13.750 71.180 14.110 ;
        RECT 72.610 13.750 74.010 14.110 ;
        RECT 75.850 13.750 79.700 14.110 ;
        RECT 81.360 13.750 85.210 14.110 ;
        RECT 87.000 13.750 88.890 14.110 ;
        RECT 90.320 13.750 91.720 14.110 ;
        RECT 93.560 13.750 97.410 14.110 ;
        RECT 99.070 13.750 102.920 14.110 ;
        RECT 104.710 13.750 106.600 14.110 ;
        RECT 0.680 0.750 0.980 13.340 ;
        RECT 2.880 8.300 3.170 13.750 ;
        RECT 1.580 7.250 1.960 7.300 ;
        RECT 1.580 6.890 2.910 7.250 ;
        RECT 1.580 6.840 1.960 6.890 ;
        RECT 2.880 0.510 3.170 5.810 ;
        RECT 4.010 0.750 4.310 13.340 ;
        RECT 6.210 8.300 6.500 13.750 ;
        RECT 7.350 8.300 7.640 13.750 ;
        RECT 4.910 7.250 5.290 7.300 ;
        RECT 8.560 7.250 8.940 7.300 ;
        RECT 4.910 6.890 6.240 7.250 ;
        RECT 7.610 6.890 8.940 7.250 ;
        RECT 4.910 6.840 5.290 6.890 ;
        RECT 8.560 6.840 8.940 6.890 ;
        RECT 6.210 0.510 6.500 5.810 ;
        RECT 6.840 0.510 7.010 5.380 ;
        RECT 7.350 0.510 7.640 5.800 ;
        RECT 9.535 0.750 9.835 13.340 ;
        RECT 11.730 8.300 12.020 13.750 ;
        RECT 12.870 8.300 13.160 13.750 ;
        RECT 10.430 7.250 10.810 7.300 ;
        RECT 14.080 7.250 14.460 7.300 ;
        RECT 10.430 6.890 11.760 7.250 ;
        RECT 13.130 6.890 14.460 7.250 ;
        RECT 10.430 6.840 10.810 6.890 ;
        RECT 14.080 6.840 14.460 6.890 ;
        RECT 11.730 0.510 12.020 5.800 ;
        RECT 12.360 0.510 12.530 5.380 ;
        RECT 12.870 0.510 13.160 5.800 ;
        RECT 15.055 0.750 15.355 13.340 ;
        RECT 17.250 8.300 17.540 13.750 ;
        RECT 15.950 7.250 16.330 7.300 ;
        RECT 15.950 6.890 17.280 7.250 ;
        RECT 15.950 6.840 16.330 6.890 ;
        RECT 17.250 0.510 17.540 5.800 ;
        RECT 17.880 0.510 18.050 5.380 ;
        RECT 18.390 0.750 18.690 13.340 ;
        RECT 20.590 8.300 20.880 13.750 ;
        RECT 19.290 7.250 19.670 7.300 ;
        RECT 19.290 6.890 20.620 7.250 ;
        RECT 19.290 6.840 19.670 6.890 ;
        RECT 20.590 0.510 20.880 5.810 ;
        RECT 21.720 0.750 22.020 13.340 ;
        RECT 23.920 8.300 24.210 13.750 ;
        RECT 25.060 8.300 25.350 13.750 ;
        RECT 22.620 7.250 23.000 7.300 ;
        RECT 26.270 7.250 26.650 7.300 ;
        RECT 22.620 6.890 23.950 7.250 ;
        RECT 25.320 6.890 26.650 7.250 ;
        RECT 22.620 6.840 23.000 6.890 ;
        RECT 26.270 6.840 26.650 6.890 ;
        RECT 23.920 0.510 24.210 5.810 ;
        RECT 24.550 0.510 24.720 5.380 ;
        RECT 25.060 0.510 25.350 5.800 ;
        RECT 27.245 0.750 27.545 13.340 ;
        RECT 29.440 8.300 29.730 13.750 ;
        RECT 30.580 8.300 30.870 13.750 ;
        RECT 28.140 7.250 28.520 7.300 ;
        RECT 31.790 7.250 32.170 7.300 ;
        RECT 28.140 6.890 29.470 7.250 ;
        RECT 30.840 6.890 32.170 7.250 ;
        RECT 28.140 6.840 28.520 6.890 ;
        RECT 31.790 6.840 32.170 6.890 ;
        RECT 29.440 0.510 29.730 5.800 ;
        RECT 30.070 0.510 30.240 5.380 ;
        RECT 30.580 0.510 30.870 5.800 ;
        RECT 32.765 0.750 33.065 13.340 ;
        RECT 34.960 8.300 35.250 13.750 ;
        RECT 33.660 7.250 34.040 7.300 ;
        RECT 33.660 6.890 34.990 7.250 ;
        RECT 33.660 6.840 34.040 6.890 ;
        RECT 34.960 0.510 35.250 5.800 ;
        RECT 35.590 0.510 35.760 5.380 ;
        RECT 36.100 0.750 36.400 13.340 ;
        RECT 38.300 8.300 38.590 13.750 ;
        RECT 37.000 7.250 37.380 7.300 ;
        RECT 37.000 6.890 38.330 7.250 ;
        RECT 37.000 6.840 37.380 6.890 ;
        RECT 38.300 0.510 38.590 5.810 ;
        RECT 39.430 0.750 39.730 13.340 ;
        RECT 41.630 8.300 41.920 13.750 ;
        RECT 42.770 8.300 43.060 13.750 ;
        RECT 40.330 7.250 40.710 7.300 ;
        RECT 43.980 7.250 44.360 7.300 ;
        RECT 40.330 6.890 41.660 7.250 ;
        RECT 43.030 6.890 44.360 7.250 ;
        RECT 40.330 6.840 40.710 6.890 ;
        RECT 43.980 6.840 44.360 6.890 ;
        RECT 41.630 0.510 41.920 5.810 ;
        RECT 42.260 0.510 42.430 5.380 ;
        RECT 42.770 0.510 43.060 5.800 ;
        RECT 44.955 0.750 45.255 13.340 ;
        RECT 47.150 8.300 47.440 13.750 ;
        RECT 48.290 8.300 48.580 13.750 ;
        RECT 45.850 7.250 46.230 7.300 ;
        RECT 49.500 7.250 49.880 7.300 ;
        RECT 45.850 6.890 47.180 7.250 ;
        RECT 48.550 6.890 49.880 7.250 ;
        RECT 45.850 6.840 46.230 6.890 ;
        RECT 49.500 6.840 49.880 6.890 ;
        RECT 47.150 0.510 47.440 5.800 ;
        RECT 47.780 0.510 47.950 5.380 ;
        RECT 48.290 0.510 48.580 5.800 ;
        RECT 50.475 0.750 50.775 13.340 ;
        RECT 52.670 8.300 52.960 13.750 ;
        RECT 51.370 7.250 51.750 7.300 ;
        RECT 51.370 6.890 52.700 7.250 ;
        RECT 51.370 6.840 51.750 6.890 ;
        RECT 52.670 0.510 52.960 5.800 ;
        RECT 53.300 0.510 53.470 5.380 ;
        RECT 53.810 0.750 54.110 13.340 ;
        RECT 56.010 8.300 56.300 13.750 ;
        RECT 54.710 7.250 55.090 7.300 ;
        RECT 54.710 6.890 56.040 7.250 ;
        RECT 54.710 6.840 55.090 6.890 ;
        RECT 56.010 0.510 56.300 5.810 ;
        RECT 57.140 0.750 57.440 13.340 ;
        RECT 59.340 8.300 59.630 13.750 ;
        RECT 60.480 8.300 60.770 13.750 ;
        RECT 58.040 7.250 58.420 7.300 ;
        RECT 61.690 7.250 62.070 7.300 ;
        RECT 58.040 6.890 59.370 7.250 ;
        RECT 60.740 6.890 62.070 7.250 ;
        RECT 58.040 6.840 58.420 6.890 ;
        RECT 61.690 6.840 62.070 6.890 ;
        RECT 59.340 0.510 59.630 5.810 ;
        RECT 59.970 0.510 60.140 5.380 ;
        RECT 60.480 0.510 60.770 5.800 ;
        RECT 62.665 0.750 62.965 13.340 ;
        RECT 64.860 8.300 65.150 13.750 ;
        RECT 66.000 8.300 66.290 13.750 ;
        RECT 63.560 7.250 63.940 7.300 ;
        RECT 67.210 7.250 67.590 7.300 ;
        RECT 63.560 6.890 64.890 7.250 ;
        RECT 66.260 6.890 67.590 7.250 ;
        RECT 63.560 6.840 63.940 6.890 ;
        RECT 67.210 6.840 67.590 6.890 ;
        RECT 64.860 0.510 65.150 5.800 ;
        RECT 65.490 0.510 65.660 5.380 ;
        RECT 66.000 0.510 66.290 5.800 ;
        RECT 68.185 0.750 68.485 13.340 ;
        RECT 70.380 8.300 70.670 13.750 ;
        RECT 69.080 7.250 69.460 7.300 ;
        RECT 69.080 6.890 70.410 7.250 ;
        RECT 69.080 6.840 69.460 6.890 ;
        RECT 70.380 0.510 70.670 5.800 ;
        RECT 71.010 0.510 71.180 5.380 ;
        RECT 71.520 0.750 71.820 13.340 ;
        RECT 73.720 8.300 74.010 13.750 ;
        RECT 72.420 7.250 72.800 7.300 ;
        RECT 72.420 6.890 73.750 7.250 ;
        RECT 72.420 6.840 72.800 6.890 ;
        RECT 73.720 0.510 74.010 5.810 ;
        RECT 74.850 0.750 75.150 13.340 ;
        RECT 77.050 8.300 77.340 13.750 ;
        RECT 78.190 8.300 78.480 13.750 ;
        RECT 75.750 7.250 76.130 7.300 ;
        RECT 79.400 7.250 79.780 7.300 ;
        RECT 75.750 6.890 77.080 7.250 ;
        RECT 78.450 6.890 79.780 7.250 ;
        RECT 75.750 6.840 76.130 6.890 ;
        RECT 79.400 6.840 79.780 6.890 ;
        RECT 77.050 0.510 77.340 5.810 ;
        RECT 77.680 0.510 77.850 5.380 ;
        RECT 78.190 0.510 78.480 5.800 ;
        RECT 80.375 0.750 80.675 13.340 ;
        RECT 82.570 8.300 82.860 13.750 ;
        RECT 83.710 8.300 84.000 13.750 ;
        RECT 81.270 7.250 81.650 7.300 ;
        RECT 84.920 7.250 85.300 7.300 ;
        RECT 81.270 6.890 82.600 7.250 ;
        RECT 83.970 6.890 85.300 7.250 ;
        RECT 81.270 6.840 81.650 6.890 ;
        RECT 84.920 6.840 85.300 6.890 ;
        RECT 82.570 0.510 82.860 5.800 ;
        RECT 83.200 0.510 83.370 5.380 ;
        RECT 83.710 0.510 84.000 5.800 ;
        RECT 85.895 0.750 86.195 13.340 ;
        RECT 88.090 8.300 88.380 13.750 ;
        RECT 86.790 7.250 87.170 7.300 ;
        RECT 86.790 6.890 88.120 7.250 ;
        RECT 86.790 6.840 87.170 6.890 ;
        RECT 88.090 0.510 88.380 5.800 ;
        RECT 88.720 0.510 88.890 5.380 ;
        RECT 89.230 0.750 89.530 13.340 ;
        RECT 91.430 8.300 91.720 13.750 ;
        RECT 90.130 7.250 90.510 7.300 ;
        RECT 90.130 6.890 91.460 7.250 ;
        RECT 90.130 6.840 90.510 6.890 ;
        RECT 91.430 0.510 91.720 5.810 ;
        RECT 92.560 0.750 92.860 13.340 ;
        RECT 94.760 8.300 95.050 13.750 ;
        RECT 95.900 8.300 96.190 13.750 ;
        RECT 93.460 7.250 93.840 7.300 ;
        RECT 97.110 7.250 97.490 7.300 ;
        RECT 93.460 6.890 94.790 7.250 ;
        RECT 96.160 6.890 97.490 7.250 ;
        RECT 93.460 6.840 93.840 6.890 ;
        RECT 97.110 6.840 97.490 6.890 ;
        RECT 94.760 0.510 95.050 5.810 ;
        RECT 95.390 0.510 95.560 5.380 ;
        RECT 95.900 0.510 96.190 5.800 ;
        RECT 98.085 0.750 98.385 13.340 ;
        RECT 100.280 8.300 100.570 13.750 ;
        RECT 101.420 8.300 101.710 13.750 ;
        RECT 98.980 7.250 99.360 7.300 ;
        RECT 102.630 7.250 103.010 7.300 ;
        RECT 98.980 6.890 100.310 7.250 ;
        RECT 101.680 6.890 103.010 7.250 ;
        RECT 98.980 6.840 99.360 6.890 ;
        RECT 102.630 6.840 103.010 6.890 ;
        RECT 100.280 0.510 100.570 5.800 ;
        RECT 100.910 0.510 101.080 5.380 ;
        RECT 101.420 0.510 101.710 5.800 ;
        RECT 103.605 0.750 103.905 13.340 ;
        RECT 105.800 8.300 106.090 13.750 ;
        RECT 104.500 7.250 104.880 7.300 ;
        RECT 104.500 6.890 105.830 7.250 ;
        RECT 104.500 6.840 104.880 6.890 ;
        RECT 105.800 0.510 106.090 5.800 ;
        RECT 106.430 0.510 106.600 5.380 ;
        RECT 1.770 0.350 3.170 0.510 ;
        RECT 5.010 0.350 8.860 0.510 ;
        RECT 10.520 0.350 14.370 0.510 ;
        RECT 16.160 0.350 18.050 0.510 ;
        RECT 19.480 0.350 20.880 0.510 ;
        RECT 22.720 0.350 26.570 0.510 ;
        RECT 28.230 0.350 32.080 0.510 ;
        RECT 33.870 0.350 35.760 0.510 ;
        RECT 37.190 0.350 38.590 0.510 ;
        RECT 40.430 0.350 44.280 0.510 ;
        RECT 45.940 0.350 49.790 0.510 ;
        RECT 51.580 0.350 53.470 0.510 ;
        RECT 54.900 0.350 56.300 0.510 ;
        RECT 58.140 0.350 61.990 0.510 ;
        RECT 63.650 0.350 67.500 0.510 ;
        RECT 69.290 0.350 71.180 0.510 ;
        RECT 72.610 0.350 74.010 0.510 ;
        RECT 75.850 0.350 79.700 0.510 ;
        RECT 81.360 0.350 85.210 0.510 ;
        RECT 87.000 0.350 88.890 0.510 ;
        RECT 90.320 0.350 91.720 0.510 ;
        RECT 93.560 0.350 97.410 0.510 ;
        RECT 99.070 0.350 102.920 0.510 ;
        RECT 104.710 0.350 106.600 0.510 ;
        RECT 0.180 0.180 106.600 0.350 ;
        RECT 1.770 0.150 3.170 0.180 ;
        RECT 5.010 0.150 8.860 0.180 ;
        RECT 10.520 0.150 14.370 0.180 ;
        RECT 16.160 0.150 18.050 0.180 ;
        RECT 19.480 0.150 20.880 0.180 ;
        RECT 22.720 0.150 26.570 0.180 ;
        RECT 28.230 0.150 32.080 0.180 ;
        RECT 33.870 0.150 35.760 0.180 ;
        RECT 37.190 0.150 38.590 0.180 ;
        RECT 40.430 0.150 44.280 0.180 ;
        RECT 45.940 0.150 49.790 0.180 ;
        RECT 51.580 0.150 53.470 0.180 ;
        RECT 54.900 0.150 56.300 0.180 ;
        RECT 58.140 0.150 61.990 0.180 ;
        RECT 63.650 0.150 67.500 0.180 ;
        RECT 69.290 0.150 71.180 0.180 ;
        RECT 72.610 0.150 74.010 0.180 ;
        RECT 75.850 0.150 79.700 0.180 ;
        RECT 81.360 0.150 85.210 0.180 ;
        RECT 87.000 0.150 88.890 0.180 ;
        RECT 90.320 0.150 91.720 0.180 ;
        RECT 93.560 0.150 97.410 0.180 ;
        RECT 99.070 0.150 102.920 0.180 ;
        RECT 104.710 0.150 106.600 0.180 ;
      LAYER mcon ;
        RECT 8.720 29.360 9.020 29.660 ;
        RECT 9.210 29.360 9.510 29.660 ;
        RECT 9.700 29.360 10.000 29.660 ;
        RECT 10.190 29.360 10.490 29.660 ;
        RECT 12.400 29.360 12.700 29.660 ;
        RECT 12.890 29.360 13.190 29.660 ;
        RECT 13.380 29.360 13.680 29.660 ;
        RECT 13.870 29.360 14.170 29.660 ;
        RECT 14.360 29.360 14.660 29.660 ;
        RECT 14.850 29.360 15.150 29.660 ;
        RECT 15.340 29.360 15.640 29.660 ;
        RECT 15.830 29.360 16.130 29.660 ;
        RECT 17.910 29.360 18.210 29.660 ;
        RECT 18.400 29.360 18.700 29.660 ;
        RECT 18.890 29.360 19.190 29.660 ;
        RECT 19.380 29.360 19.680 29.660 ;
        RECT 19.870 29.360 20.170 29.660 ;
        RECT 20.360 29.360 20.660 29.660 ;
        RECT 20.850 29.360 21.150 29.660 ;
        RECT 21.340 29.360 21.640 29.660 ;
        RECT 23.600 29.360 23.900 29.660 ;
        RECT 24.090 29.360 24.390 29.660 ;
        RECT 24.580 29.360 24.880 29.660 ;
        RECT 26.430 29.360 26.730 29.660 ;
        RECT 26.920 29.360 27.220 29.660 ;
        RECT 27.410 29.360 27.710 29.660 ;
        RECT 27.900 29.360 28.200 29.660 ;
        RECT 30.110 29.360 30.410 29.660 ;
        RECT 30.600 29.360 30.900 29.660 ;
        RECT 31.090 29.360 31.390 29.660 ;
        RECT 31.580 29.360 31.880 29.660 ;
        RECT 32.070 29.360 32.370 29.660 ;
        RECT 32.560 29.360 32.860 29.660 ;
        RECT 33.050 29.360 33.350 29.660 ;
        RECT 33.540 29.360 33.840 29.660 ;
        RECT 35.620 29.360 35.920 29.660 ;
        RECT 36.110 29.360 36.410 29.660 ;
        RECT 36.600 29.360 36.900 29.660 ;
        RECT 37.090 29.360 37.390 29.660 ;
        RECT 37.580 29.360 37.880 29.660 ;
        RECT 38.070 29.360 38.370 29.660 ;
        RECT 38.560 29.360 38.860 29.660 ;
        RECT 39.050 29.360 39.350 29.660 ;
        RECT 41.310 29.360 41.610 29.660 ;
        RECT 41.800 29.360 42.100 29.660 ;
        RECT 42.290 29.360 42.590 29.660 ;
        RECT 44.140 29.360 44.440 29.660 ;
        RECT 44.630 29.360 44.930 29.660 ;
        RECT 45.120 29.360 45.420 29.660 ;
        RECT 45.610 29.360 45.910 29.660 ;
        RECT 47.820 29.360 48.120 29.660 ;
        RECT 48.310 29.360 48.610 29.660 ;
        RECT 48.800 29.360 49.100 29.660 ;
        RECT 49.290 29.360 49.590 29.660 ;
        RECT 49.780 29.360 50.080 29.660 ;
        RECT 50.270 29.360 50.570 29.660 ;
        RECT 50.760 29.360 51.060 29.660 ;
        RECT 51.250 29.360 51.550 29.660 ;
        RECT 53.330 29.360 53.630 29.660 ;
        RECT 53.820 29.360 54.120 29.660 ;
        RECT 54.310 29.360 54.610 29.660 ;
        RECT 54.800 29.360 55.100 29.660 ;
        RECT 55.290 29.360 55.590 29.660 ;
        RECT 55.780 29.360 56.080 29.660 ;
        RECT 56.270 29.360 56.570 29.660 ;
        RECT 56.760 29.360 57.060 29.660 ;
        RECT 59.020 29.360 59.320 29.660 ;
        RECT 59.510 29.360 59.810 29.660 ;
        RECT 60.000 29.360 60.300 29.660 ;
        RECT 61.850 29.360 62.150 29.660 ;
        RECT 62.340 29.360 62.640 29.660 ;
        RECT 62.830 29.360 63.130 29.660 ;
        RECT 63.320 29.360 63.620 29.660 ;
        RECT 65.530 29.360 65.830 29.660 ;
        RECT 66.020 29.360 66.320 29.660 ;
        RECT 66.510 29.360 66.810 29.660 ;
        RECT 67.000 29.360 67.300 29.660 ;
        RECT 67.490 29.360 67.790 29.660 ;
        RECT 67.980 29.360 68.280 29.660 ;
        RECT 68.470 29.360 68.770 29.660 ;
        RECT 68.960 29.360 69.260 29.660 ;
        RECT 71.040 29.360 71.340 29.660 ;
        RECT 71.530 29.360 71.830 29.660 ;
        RECT 72.020 29.360 72.320 29.660 ;
        RECT 72.510 29.360 72.810 29.660 ;
        RECT 73.000 29.360 73.300 29.660 ;
        RECT 73.490 29.360 73.790 29.660 ;
        RECT 73.980 29.360 74.280 29.660 ;
        RECT 74.470 29.360 74.770 29.660 ;
        RECT 76.730 29.360 77.030 29.660 ;
        RECT 77.220 29.360 77.520 29.660 ;
        RECT 77.710 29.360 78.010 29.660 ;
        RECT 79.560 29.360 79.860 29.660 ;
        RECT 80.050 29.360 80.350 29.660 ;
        RECT 80.540 29.360 80.840 29.660 ;
        RECT 81.030 29.360 81.330 29.660 ;
        RECT 83.240 29.360 83.540 29.660 ;
        RECT 83.730 29.360 84.030 29.660 ;
        RECT 84.220 29.360 84.520 29.660 ;
        RECT 84.710 29.360 85.010 29.660 ;
        RECT 85.200 29.360 85.500 29.660 ;
        RECT 85.690 29.360 85.990 29.660 ;
        RECT 86.180 29.360 86.480 29.660 ;
        RECT 86.670 29.360 86.970 29.660 ;
        RECT 88.750 29.360 89.050 29.660 ;
        RECT 89.240 29.360 89.540 29.660 ;
        RECT 89.730 29.360 90.030 29.660 ;
        RECT 90.220 29.360 90.520 29.660 ;
        RECT 90.710 29.360 91.010 29.660 ;
        RECT 91.200 29.360 91.500 29.660 ;
        RECT 91.690 29.360 91.990 29.660 ;
        RECT 92.180 29.360 92.480 29.660 ;
        RECT 94.440 29.360 94.740 29.660 ;
        RECT 94.930 29.360 95.230 29.660 ;
        RECT 95.420 29.360 95.720 29.660 ;
        RECT -0.665 25.435 -0.495 25.605 ;
        RECT -0.205 25.435 -0.035 25.605 ;
        RECT 0.255 25.435 0.425 25.605 ;
        RECT 0.715 25.435 0.885 25.605 ;
        RECT 1.175 25.435 1.345 25.605 ;
        RECT 3.330 25.435 3.500 25.605 ;
        RECT 3.790 25.435 3.960 25.605 ;
        RECT 4.250 25.435 4.420 25.605 ;
        RECT -7.880 24.020 -7.620 24.280 ;
        RECT 2.240 24.040 2.480 24.280 ;
        RECT 11.355 23.980 11.655 24.280 ;
        RECT -0.665 22.715 -0.495 22.885 ;
        RECT -0.205 22.715 -0.035 22.885 ;
        RECT 0.255 22.715 0.425 22.885 ;
        RECT 0.715 22.715 0.885 22.885 ;
        RECT 1.175 22.715 1.345 22.885 ;
        RECT 3.330 22.715 3.500 22.885 ;
        RECT 3.790 22.715 3.960 22.885 ;
        RECT 4.250 22.715 4.420 22.885 ;
        RECT 9.430 22.620 9.730 22.920 ;
        RECT 9.920 22.620 10.220 22.920 ;
        RECT 10.410 22.620 10.710 22.920 ;
        RECT 12.300 22.620 12.600 22.920 ;
        RECT 12.790 22.620 13.090 22.920 ;
        RECT 13.280 22.620 13.580 22.920 ;
        RECT 14.950 22.620 15.250 22.920 ;
        RECT 15.440 22.620 15.740 22.920 ;
        RECT 15.930 22.620 16.230 22.920 ;
        RECT 17.820 22.620 18.120 22.920 ;
        RECT 18.310 22.620 18.610 22.920 ;
        RECT 18.800 22.620 19.100 22.920 ;
        RECT 20.470 22.620 20.770 22.920 ;
        RECT 20.960 22.620 21.260 22.920 ;
        RECT 21.450 22.620 21.750 22.920 ;
        RECT 16.875 21.260 17.175 21.560 ;
        RECT 25.730 23.980 26.030 24.280 ;
        RECT 23.800 22.620 24.100 22.920 ;
        RECT 24.290 22.620 24.590 22.920 ;
        RECT 24.780 22.620 25.080 22.920 ;
        RECT 22.400 21.260 22.700 21.560 ;
        RECT 29.065 23.980 29.365 24.280 ;
        RECT 27.140 22.620 27.440 22.920 ;
        RECT 27.630 22.620 27.930 22.920 ;
        RECT 28.120 22.620 28.420 22.920 ;
        RECT 30.010 22.620 30.310 22.920 ;
        RECT 30.500 22.620 30.800 22.920 ;
        RECT 30.990 22.620 31.290 22.920 ;
        RECT 32.660 22.620 32.960 22.920 ;
        RECT 33.150 22.620 33.450 22.920 ;
        RECT 33.640 22.620 33.940 22.920 ;
        RECT 35.530 22.620 35.830 22.920 ;
        RECT 36.020 22.620 36.320 22.920 ;
        RECT 36.510 22.620 36.810 22.920 ;
        RECT 38.180 22.620 38.480 22.920 ;
        RECT 38.670 22.620 38.970 22.920 ;
        RECT 39.160 22.620 39.460 22.920 ;
        RECT 34.585 21.260 34.885 21.560 ;
        RECT 43.440 23.980 43.740 24.280 ;
        RECT 41.510 22.620 41.810 22.920 ;
        RECT 42.000 22.620 42.300 22.920 ;
        RECT 42.490 22.620 42.790 22.920 ;
        RECT 40.110 21.260 40.410 21.560 ;
        RECT 46.775 23.980 47.075 24.280 ;
        RECT 44.850 22.620 45.150 22.920 ;
        RECT 45.340 22.620 45.640 22.920 ;
        RECT 45.830 22.620 46.130 22.920 ;
        RECT 47.720 22.620 48.020 22.920 ;
        RECT 48.210 22.620 48.510 22.920 ;
        RECT 48.700 22.620 49.000 22.920 ;
        RECT 50.370 22.620 50.670 22.920 ;
        RECT 50.860 22.620 51.160 22.920 ;
        RECT 51.350 22.620 51.650 22.920 ;
        RECT 53.240 22.620 53.540 22.920 ;
        RECT 53.730 22.620 54.030 22.920 ;
        RECT 54.220 22.620 54.520 22.920 ;
        RECT 55.890 22.620 56.190 22.920 ;
        RECT 56.380 22.620 56.680 22.920 ;
        RECT 56.870 22.620 57.170 22.920 ;
        RECT 52.295 21.260 52.595 21.560 ;
        RECT 61.150 23.980 61.450 24.280 ;
        RECT 59.220 22.620 59.520 22.920 ;
        RECT 59.710 22.620 60.010 22.920 ;
        RECT 60.200 22.620 60.500 22.920 ;
        RECT 57.820 21.260 58.120 21.560 ;
        RECT 64.485 23.980 64.785 24.280 ;
        RECT 62.560 22.620 62.860 22.920 ;
        RECT 63.050 22.620 63.350 22.920 ;
        RECT 63.540 22.620 63.840 22.920 ;
        RECT 65.430 22.620 65.730 22.920 ;
        RECT 65.920 22.620 66.220 22.920 ;
        RECT 66.410 22.620 66.710 22.920 ;
        RECT 68.080 22.620 68.380 22.920 ;
        RECT 68.570 22.620 68.870 22.920 ;
        RECT 69.060 22.620 69.360 22.920 ;
        RECT 70.950 22.620 71.250 22.920 ;
        RECT 71.440 22.620 71.740 22.920 ;
        RECT 71.930 22.620 72.230 22.920 ;
        RECT 73.600 22.620 73.900 22.920 ;
        RECT 74.090 22.620 74.390 22.920 ;
        RECT 74.580 22.620 74.880 22.920 ;
        RECT 70.005 21.260 70.305 21.560 ;
        RECT 78.860 23.980 79.160 24.280 ;
        RECT 76.930 22.620 77.230 22.920 ;
        RECT 77.420 22.620 77.720 22.920 ;
        RECT 77.910 22.620 78.210 22.920 ;
        RECT 75.530 21.260 75.830 21.560 ;
        RECT 82.195 23.980 82.495 24.280 ;
        RECT 80.270 22.620 80.570 22.920 ;
        RECT 80.760 22.620 81.060 22.920 ;
        RECT 81.250 22.620 81.550 22.920 ;
        RECT 83.140 22.620 83.440 22.920 ;
        RECT 83.630 22.620 83.930 22.920 ;
        RECT 84.120 22.620 84.420 22.920 ;
        RECT 85.790 22.620 86.090 22.920 ;
        RECT 86.280 22.620 86.580 22.920 ;
        RECT 86.770 22.620 87.070 22.920 ;
        RECT 88.660 22.620 88.960 22.920 ;
        RECT 89.150 22.620 89.450 22.920 ;
        RECT 89.640 22.620 89.940 22.920 ;
        RECT 91.310 22.620 91.610 22.920 ;
        RECT 91.800 22.620 92.100 22.920 ;
        RECT 92.290 22.620 92.590 22.920 ;
        RECT 87.715 21.260 88.015 21.560 ;
        RECT 96.570 23.980 96.870 24.280 ;
        RECT 101.100 24.050 101.400 24.350 ;
        RECT 101.600 24.050 101.900 24.350 ;
        RECT 102.100 24.050 102.400 24.350 ;
        RECT 102.600 24.050 102.900 24.350 ;
        RECT 94.640 22.620 94.940 22.920 ;
        RECT 95.130 22.620 95.430 22.920 ;
        RECT 95.620 22.620 95.920 22.920 ;
        RECT 93.240 21.260 93.540 21.560 ;
        RECT 102.090 19.120 102.390 19.420 ;
        RECT 102.610 19.120 102.910 19.420 ;
        RECT 102.090 18.600 102.390 18.900 ;
        RECT 102.610 18.600 102.910 18.900 ;
        RECT 107.605 19.100 107.905 19.400 ;
        RECT 108.095 19.100 108.395 19.400 ;
        RECT 107.605 18.600 107.905 18.900 ;
        RECT 108.095 18.600 108.395 18.900 ;
        RECT 8.720 15.760 9.020 16.060 ;
        RECT 9.210 15.760 9.510 16.060 ;
        RECT 9.700 15.760 10.000 16.060 ;
        RECT 10.190 15.760 10.490 16.060 ;
        RECT 12.400 15.760 12.700 16.060 ;
        RECT 12.890 15.760 13.190 16.060 ;
        RECT 13.380 15.760 13.680 16.060 ;
        RECT 13.870 15.760 14.170 16.060 ;
        RECT 14.360 15.760 14.660 16.060 ;
        RECT 14.850 15.760 15.150 16.060 ;
        RECT 15.340 15.760 15.640 16.060 ;
        RECT 15.830 15.760 16.130 16.060 ;
        RECT 17.910 15.760 18.210 16.060 ;
        RECT 18.400 15.760 18.700 16.060 ;
        RECT 18.890 15.760 19.190 16.060 ;
        RECT 19.380 15.760 19.680 16.060 ;
        RECT 19.870 15.760 20.170 16.060 ;
        RECT 20.360 15.760 20.660 16.060 ;
        RECT 20.850 15.760 21.150 16.060 ;
        RECT 21.340 15.760 21.640 16.060 ;
        RECT 23.600 15.760 23.900 16.060 ;
        RECT 24.090 15.760 24.390 16.060 ;
        RECT 24.580 15.760 24.880 16.060 ;
        RECT 26.430 15.760 26.730 16.060 ;
        RECT 26.920 15.760 27.220 16.060 ;
        RECT 27.410 15.760 27.710 16.060 ;
        RECT 27.900 15.760 28.200 16.060 ;
        RECT 30.110 15.760 30.410 16.060 ;
        RECT 30.600 15.760 30.900 16.060 ;
        RECT 31.090 15.760 31.390 16.060 ;
        RECT 31.580 15.760 31.880 16.060 ;
        RECT 32.070 15.760 32.370 16.060 ;
        RECT 32.560 15.760 32.860 16.060 ;
        RECT 33.050 15.760 33.350 16.060 ;
        RECT 33.540 15.760 33.840 16.060 ;
        RECT 35.620 15.760 35.920 16.060 ;
        RECT 36.110 15.760 36.410 16.060 ;
        RECT 36.600 15.760 36.900 16.060 ;
        RECT 37.090 15.760 37.390 16.060 ;
        RECT 37.580 15.760 37.880 16.060 ;
        RECT 38.070 15.760 38.370 16.060 ;
        RECT 38.560 15.760 38.860 16.060 ;
        RECT 39.050 15.760 39.350 16.060 ;
        RECT 41.310 15.760 41.610 16.060 ;
        RECT 41.800 15.760 42.100 16.060 ;
        RECT 42.290 15.760 42.590 16.060 ;
        RECT 44.140 15.760 44.440 16.060 ;
        RECT 44.630 15.760 44.930 16.060 ;
        RECT 45.120 15.760 45.420 16.060 ;
        RECT 45.610 15.760 45.910 16.060 ;
        RECT 47.820 15.760 48.120 16.060 ;
        RECT 48.310 15.760 48.610 16.060 ;
        RECT 48.800 15.760 49.100 16.060 ;
        RECT 49.290 15.760 49.590 16.060 ;
        RECT 49.780 15.760 50.080 16.060 ;
        RECT 50.270 15.760 50.570 16.060 ;
        RECT 50.760 15.760 51.060 16.060 ;
        RECT 51.250 15.760 51.550 16.060 ;
        RECT 53.330 15.760 53.630 16.060 ;
        RECT 53.820 15.760 54.120 16.060 ;
        RECT 54.310 15.760 54.610 16.060 ;
        RECT 54.800 15.760 55.100 16.060 ;
        RECT 55.290 15.760 55.590 16.060 ;
        RECT 55.780 15.760 56.080 16.060 ;
        RECT 56.270 15.760 56.570 16.060 ;
        RECT 56.760 15.760 57.060 16.060 ;
        RECT 59.020 15.760 59.320 16.060 ;
        RECT 59.510 15.760 59.810 16.060 ;
        RECT 60.000 15.760 60.300 16.060 ;
        RECT 61.850 15.760 62.150 16.060 ;
        RECT 62.340 15.760 62.640 16.060 ;
        RECT 62.830 15.760 63.130 16.060 ;
        RECT 63.320 15.760 63.620 16.060 ;
        RECT 65.530 15.760 65.830 16.060 ;
        RECT 66.020 15.760 66.320 16.060 ;
        RECT 66.510 15.760 66.810 16.060 ;
        RECT 67.000 15.760 67.300 16.060 ;
        RECT 67.490 15.760 67.790 16.060 ;
        RECT 67.980 15.760 68.280 16.060 ;
        RECT 68.470 15.760 68.770 16.060 ;
        RECT 68.960 15.760 69.260 16.060 ;
        RECT 71.040 15.760 71.340 16.060 ;
        RECT 71.530 15.760 71.830 16.060 ;
        RECT 72.020 15.760 72.320 16.060 ;
        RECT 72.510 15.760 72.810 16.060 ;
        RECT 73.000 15.760 73.300 16.060 ;
        RECT 73.490 15.760 73.790 16.060 ;
        RECT 73.980 15.760 74.280 16.060 ;
        RECT 74.470 15.760 74.770 16.060 ;
        RECT 76.730 15.760 77.030 16.060 ;
        RECT 77.220 15.760 77.520 16.060 ;
        RECT 77.710 15.760 78.010 16.060 ;
        RECT 79.560 15.760 79.860 16.060 ;
        RECT 80.050 15.760 80.350 16.060 ;
        RECT 80.540 15.760 80.840 16.060 ;
        RECT 81.030 15.760 81.330 16.060 ;
        RECT 83.240 15.760 83.540 16.060 ;
        RECT 83.730 15.760 84.030 16.060 ;
        RECT 84.220 15.760 84.520 16.060 ;
        RECT 84.710 15.760 85.010 16.060 ;
        RECT 85.200 15.760 85.500 16.060 ;
        RECT 85.690 15.760 85.990 16.060 ;
        RECT 86.180 15.760 86.480 16.060 ;
        RECT 86.670 15.760 86.970 16.060 ;
        RECT 88.750 15.760 89.050 16.060 ;
        RECT 89.240 15.760 89.540 16.060 ;
        RECT 89.730 15.760 90.030 16.060 ;
        RECT 90.220 15.760 90.520 16.060 ;
        RECT 90.710 15.760 91.010 16.060 ;
        RECT 91.200 15.760 91.500 16.060 ;
        RECT 91.690 15.760 91.990 16.060 ;
        RECT 92.180 15.760 92.480 16.060 ;
        RECT 94.440 15.760 94.740 16.060 ;
        RECT 94.930 15.760 95.230 16.060 ;
        RECT 95.420 15.760 95.720 16.060 ;
        RECT 1.830 13.780 2.130 14.080 ;
        RECT 2.320 13.780 2.620 14.080 ;
        RECT 2.810 13.780 3.110 14.080 ;
        RECT 5.070 13.780 5.370 14.080 ;
        RECT 5.560 13.780 5.860 14.080 ;
        RECT 6.050 13.780 6.350 14.080 ;
        RECT 6.540 13.780 6.840 14.080 ;
        RECT 7.030 13.780 7.330 14.080 ;
        RECT 7.520 13.780 7.820 14.080 ;
        RECT 8.010 13.780 8.310 14.080 ;
        RECT 8.500 13.780 8.800 14.080 ;
        RECT 10.580 13.780 10.880 14.080 ;
        RECT 11.070 13.780 11.370 14.080 ;
        RECT 11.560 13.780 11.860 14.080 ;
        RECT 12.050 13.780 12.350 14.080 ;
        RECT 12.540 13.780 12.840 14.080 ;
        RECT 13.030 13.780 13.330 14.080 ;
        RECT 13.520 13.780 13.820 14.080 ;
        RECT 14.010 13.780 14.310 14.080 ;
        RECT 16.220 13.780 16.520 14.080 ;
        RECT 16.710 13.780 17.010 14.080 ;
        RECT 17.200 13.780 17.500 14.080 ;
        RECT 17.690 13.780 17.990 14.080 ;
        RECT 19.540 13.780 19.840 14.080 ;
        RECT 20.030 13.780 20.330 14.080 ;
        RECT 20.520 13.780 20.820 14.080 ;
        RECT 22.780 13.780 23.080 14.080 ;
        RECT 23.270 13.780 23.570 14.080 ;
        RECT 23.760 13.780 24.060 14.080 ;
        RECT 24.250 13.780 24.550 14.080 ;
        RECT 24.740 13.780 25.040 14.080 ;
        RECT 25.230 13.780 25.530 14.080 ;
        RECT 25.720 13.780 26.020 14.080 ;
        RECT 26.210 13.780 26.510 14.080 ;
        RECT 28.290 13.780 28.590 14.080 ;
        RECT 28.780 13.780 29.080 14.080 ;
        RECT 29.270 13.780 29.570 14.080 ;
        RECT 29.760 13.780 30.060 14.080 ;
        RECT 30.250 13.780 30.550 14.080 ;
        RECT 30.740 13.780 31.040 14.080 ;
        RECT 31.230 13.780 31.530 14.080 ;
        RECT 31.720 13.780 32.020 14.080 ;
        RECT 33.930 13.780 34.230 14.080 ;
        RECT 34.420 13.780 34.720 14.080 ;
        RECT 34.910 13.780 35.210 14.080 ;
        RECT 35.400 13.780 35.700 14.080 ;
        RECT 37.250 13.780 37.550 14.080 ;
        RECT 37.740 13.780 38.040 14.080 ;
        RECT 38.230 13.780 38.530 14.080 ;
        RECT 40.490 13.780 40.790 14.080 ;
        RECT 40.980 13.780 41.280 14.080 ;
        RECT 41.470 13.780 41.770 14.080 ;
        RECT 41.960 13.780 42.260 14.080 ;
        RECT 42.450 13.780 42.750 14.080 ;
        RECT 42.940 13.780 43.240 14.080 ;
        RECT 43.430 13.780 43.730 14.080 ;
        RECT 43.920 13.780 44.220 14.080 ;
        RECT 46.000 13.780 46.300 14.080 ;
        RECT 46.490 13.780 46.790 14.080 ;
        RECT 46.980 13.780 47.280 14.080 ;
        RECT 47.470 13.780 47.770 14.080 ;
        RECT 47.960 13.780 48.260 14.080 ;
        RECT 48.450 13.780 48.750 14.080 ;
        RECT 48.940 13.780 49.240 14.080 ;
        RECT 49.430 13.780 49.730 14.080 ;
        RECT 51.640 13.780 51.940 14.080 ;
        RECT 52.130 13.780 52.430 14.080 ;
        RECT 52.620 13.780 52.920 14.080 ;
        RECT 53.110 13.780 53.410 14.080 ;
        RECT 54.960 13.780 55.260 14.080 ;
        RECT 55.450 13.780 55.750 14.080 ;
        RECT 55.940 13.780 56.240 14.080 ;
        RECT 58.200 13.780 58.500 14.080 ;
        RECT 58.690 13.780 58.990 14.080 ;
        RECT 59.180 13.780 59.480 14.080 ;
        RECT 59.670 13.780 59.970 14.080 ;
        RECT 60.160 13.780 60.460 14.080 ;
        RECT 60.650 13.780 60.950 14.080 ;
        RECT 61.140 13.780 61.440 14.080 ;
        RECT 61.630 13.780 61.930 14.080 ;
        RECT 63.710 13.780 64.010 14.080 ;
        RECT 64.200 13.780 64.500 14.080 ;
        RECT 64.690 13.780 64.990 14.080 ;
        RECT 65.180 13.780 65.480 14.080 ;
        RECT 65.670 13.780 65.970 14.080 ;
        RECT 66.160 13.780 66.460 14.080 ;
        RECT 66.650 13.780 66.950 14.080 ;
        RECT 67.140 13.780 67.440 14.080 ;
        RECT 69.350 13.780 69.650 14.080 ;
        RECT 69.840 13.780 70.140 14.080 ;
        RECT 70.330 13.780 70.630 14.080 ;
        RECT 70.820 13.780 71.120 14.080 ;
        RECT 72.670 13.780 72.970 14.080 ;
        RECT 73.160 13.780 73.460 14.080 ;
        RECT 73.650 13.780 73.950 14.080 ;
        RECT 75.910 13.780 76.210 14.080 ;
        RECT 76.400 13.780 76.700 14.080 ;
        RECT 76.890 13.780 77.190 14.080 ;
        RECT 77.380 13.780 77.680 14.080 ;
        RECT 77.870 13.780 78.170 14.080 ;
        RECT 78.360 13.780 78.660 14.080 ;
        RECT 78.850 13.780 79.150 14.080 ;
        RECT 79.340 13.780 79.640 14.080 ;
        RECT 81.420 13.780 81.720 14.080 ;
        RECT 81.910 13.780 82.210 14.080 ;
        RECT 82.400 13.780 82.700 14.080 ;
        RECT 82.890 13.780 83.190 14.080 ;
        RECT 83.380 13.780 83.680 14.080 ;
        RECT 83.870 13.780 84.170 14.080 ;
        RECT 84.360 13.780 84.660 14.080 ;
        RECT 84.850 13.780 85.150 14.080 ;
        RECT 87.060 13.780 87.360 14.080 ;
        RECT 87.550 13.780 87.850 14.080 ;
        RECT 88.040 13.780 88.340 14.080 ;
        RECT 88.530 13.780 88.830 14.080 ;
        RECT 90.380 13.780 90.680 14.080 ;
        RECT 90.870 13.780 91.170 14.080 ;
        RECT 91.360 13.780 91.660 14.080 ;
        RECT 93.620 13.780 93.920 14.080 ;
        RECT 94.110 13.780 94.410 14.080 ;
        RECT 94.600 13.780 94.900 14.080 ;
        RECT 95.090 13.780 95.390 14.080 ;
        RECT 95.580 13.780 95.880 14.080 ;
        RECT 96.070 13.780 96.370 14.080 ;
        RECT 96.560 13.780 96.860 14.080 ;
        RECT 97.050 13.780 97.350 14.080 ;
        RECT 99.130 13.780 99.430 14.080 ;
        RECT 99.620 13.780 99.920 14.080 ;
        RECT 100.110 13.780 100.410 14.080 ;
        RECT 100.600 13.780 100.900 14.080 ;
        RECT 101.090 13.780 101.390 14.080 ;
        RECT 101.580 13.780 101.880 14.080 ;
        RECT 102.070 13.780 102.370 14.080 ;
        RECT 102.560 13.780 102.860 14.080 ;
        RECT 104.770 13.780 105.070 14.080 ;
        RECT 105.260 13.780 105.560 14.080 ;
        RECT 105.750 13.780 106.050 14.080 ;
        RECT 106.240 13.780 106.540 14.080 ;
        RECT 4.010 8.280 4.310 8.580 ;
        RECT 1.630 6.920 1.930 7.220 ;
        RECT 2.120 6.920 2.420 7.220 ;
        RECT 2.610 6.920 2.910 7.220 ;
        RECT 0.680 5.560 0.980 5.860 ;
        RECT 9.535 8.280 9.835 8.580 ;
        RECT 4.960 6.920 5.260 7.220 ;
        RECT 5.450 6.920 5.750 7.220 ;
        RECT 5.940 6.920 6.240 7.220 ;
        RECT 7.610 6.920 7.910 7.220 ;
        RECT 8.100 6.920 8.400 7.220 ;
        RECT 8.590 6.920 8.890 7.220 ;
        RECT 10.480 6.920 10.780 7.220 ;
        RECT 10.970 6.920 11.270 7.220 ;
        RECT 11.460 6.920 11.760 7.220 ;
        RECT 13.130 6.920 13.430 7.220 ;
        RECT 13.620 6.920 13.920 7.220 ;
        RECT 14.110 6.920 14.410 7.220 ;
        RECT 16.000 6.920 16.300 7.220 ;
        RECT 16.490 6.920 16.790 7.220 ;
        RECT 16.980 6.920 17.280 7.220 ;
        RECT 15.055 5.560 15.355 5.860 ;
        RECT 21.720 8.280 22.020 8.580 ;
        RECT 19.340 6.920 19.640 7.220 ;
        RECT 19.830 6.920 20.130 7.220 ;
        RECT 20.320 6.920 20.620 7.220 ;
        RECT 18.390 5.560 18.690 5.860 ;
        RECT 27.245 8.280 27.545 8.580 ;
        RECT 22.670 6.920 22.970 7.220 ;
        RECT 23.160 6.920 23.460 7.220 ;
        RECT 23.650 6.920 23.950 7.220 ;
        RECT 25.320 6.920 25.620 7.220 ;
        RECT 25.810 6.920 26.110 7.220 ;
        RECT 26.300 6.920 26.600 7.220 ;
        RECT 28.190 6.920 28.490 7.220 ;
        RECT 28.680 6.920 28.980 7.220 ;
        RECT 29.170 6.920 29.470 7.220 ;
        RECT 30.840 6.920 31.140 7.220 ;
        RECT 31.330 6.920 31.630 7.220 ;
        RECT 31.820 6.920 32.120 7.220 ;
        RECT 33.710 6.920 34.010 7.220 ;
        RECT 34.200 6.920 34.500 7.220 ;
        RECT 34.690 6.920 34.990 7.220 ;
        RECT 32.765 5.560 33.065 5.860 ;
        RECT 39.430 8.280 39.730 8.580 ;
        RECT 37.050 6.920 37.350 7.220 ;
        RECT 37.540 6.920 37.840 7.220 ;
        RECT 38.030 6.920 38.330 7.220 ;
        RECT 36.100 5.560 36.400 5.860 ;
        RECT 44.955 8.280 45.255 8.580 ;
        RECT 40.380 6.920 40.680 7.220 ;
        RECT 40.870 6.920 41.170 7.220 ;
        RECT 41.360 6.920 41.660 7.220 ;
        RECT 43.030 6.920 43.330 7.220 ;
        RECT 43.520 6.920 43.820 7.220 ;
        RECT 44.010 6.920 44.310 7.220 ;
        RECT 45.900 6.920 46.200 7.220 ;
        RECT 46.390 6.920 46.690 7.220 ;
        RECT 46.880 6.920 47.180 7.220 ;
        RECT 48.550 6.920 48.850 7.220 ;
        RECT 49.040 6.920 49.340 7.220 ;
        RECT 49.530 6.920 49.830 7.220 ;
        RECT 51.420 6.920 51.720 7.220 ;
        RECT 51.910 6.920 52.210 7.220 ;
        RECT 52.400 6.920 52.700 7.220 ;
        RECT 50.475 5.560 50.775 5.860 ;
        RECT 57.140 8.280 57.440 8.580 ;
        RECT 54.760 6.920 55.060 7.220 ;
        RECT 55.250 6.920 55.550 7.220 ;
        RECT 55.740 6.920 56.040 7.220 ;
        RECT 53.810 5.560 54.110 5.860 ;
        RECT 62.665 8.280 62.965 8.580 ;
        RECT 58.090 6.920 58.390 7.220 ;
        RECT 58.580 6.920 58.880 7.220 ;
        RECT 59.070 6.920 59.370 7.220 ;
        RECT 60.740 6.920 61.040 7.220 ;
        RECT 61.230 6.920 61.530 7.220 ;
        RECT 61.720 6.920 62.020 7.220 ;
        RECT 63.610 6.920 63.910 7.220 ;
        RECT 64.100 6.920 64.400 7.220 ;
        RECT 64.590 6.920 64.890 7.220 ;
        RECT 66.260 6.920 66.560 7.220 ;
        RECT 66.750 6.920 67.050 7.220 ;
        RECT 67.240 6.920 67.540 7.220 ;
        RECT 69.130 6.920 69.430 7.220 ;
        RECT 69.620 6.920 69.920 7.220 ;
        RECT 70.110 6.920 70.410 7.220 ;
        RECT 68.185 5.560 68.485 5.860 ;
        RECT 74.850 8.280 75.150 8.580 ;
        RECT 72.470 6.920 72.770 7.220 ;
        RECT 72.960 6.920 73.260 7.220 ;
        RECT 73.450 6.920 73.750 7.220 ;
        RECT 71.520 5.560 71.820 5.860 ;
        RECT 80.375 8.280 80.675 8.580 ;
        RECT 75.800 6.920 76.100 7.220 ;
        RECT 76.290 6.920 76.590 7.220 ;
        RECT 76.780 6.920 77.080 7.220 ;
        RECT 78.450 6.920 78.750 7.220 ;
        RECT 78.940 6.920 79.240 7.220 ;
        RECT 79.430 6.920 79.730 7.220 ;
        RECT 81.320 6.920 81.620 7.220 ;
        RECT 81.810 6.920 82.110 7.220 ;
        RECT 82.300 6.920 82.600 7.220 ;
        RECT 83.970 6.920 84.270 7.220 ;
        RECT 84.460 6.920 84.760 7.220 ;
        RECT 84.950 6.920 85.250 7.220 ;
        RECT 86.840 6.920 87.140 7.220 ;
        RECT 87.330 6.920 87.630 7.220 ;
        RECT 87.820 6.920 88.120 7.220 ;
        RECT 85.895 5.560 86.195 5.860 ;
        RECT 92.560 8.280 92.860 8.580 ;
        RECT 90.180 6.920 90.480 7.220 ;
        RECT 90.670 6.920 90.970 7.220 ;
        RECT 91.160 6.920 91.460 7.220 ;
        RECT 89.230 5.560 89.530 5.860 ;
        RECT 98.085 8.280 98.385 8.580 ;
        RECT 93.510 6.920 93.810 7.220 ;
        RECT 94.000 6.920 94.300 7.220 ;
        RECT 94.490 6.920 94.790 7.220 ;
        RECT 96.160 6.920 96.460 7.220 ;
        RECT 96.650 6.920 96.950 7.220 ;
        RECT 97.140 6.920 97.440 7.220 ;
        RECT 99.030 6.920 99.330 7.220 ;
        RECT 99.520 6.920 99.820 7.220 ;
        RECT 100.010 6.920 100.310 7.220 ;
        RECT 101.680 6.920 101.980 7.220 ;
        RECT 102.170 6.920 102.470 7.220 ;
        RECT 102.660 6.920 102.960 7.220 ;
        RECT 104.550 6.920 104.850 7.220 ;
        RECT 105.040 6.920 105.340 7.220 ;
        RECT 105.530 6.920 105.830 7.220 ;
        RECT 103.605 5.560 103.905 5.860 ;
        RECT 1.830 0.180 2.130 0.480 ;
        RECT 2.320 0.180 2.620 0.480 ;
        RECT 2.810 0.180 3.110 0.480 ;
        RECT 5.070 0.180 5.370 0.480 ;
        RECT 5.560 0.180 5.860 0.480 ;
        RECT 6.050 0.180 6.350 0.480 ;
        RECT 6.540 0.180 6.840 0.480 ;
        RECT 7.030 0.180 7.330 0.480 ;
        RECT 7.520 0.180 7.820 0.480 ;
        RECT 8.010 0.180 8.310 0.480 ;
        RECT 8.500 0.180 8.800 0.480 ;
        RECT 10.580 0.180 10.880 0.480 ;
        RECT 11.070 0.180 11.370 0.480 ;
        RECT 11.560 0.180 11.860 0.480 ;
        RECT 12.050 0.180 12.350 0.480 ;
        RECT 12.540 0.180 12.840 0.480 ;
        RECT 13.030 0.180 13.330 0.480 ;
        RECT 13.520 0.180 13.820 0.480 ;
        RECT 14.010 0.180 14.310 0.480 ;
        RECT 16.220 0.180 16.520 0.480 ;
        RECT 16.710 0.180 17.010 0.480 ;
        RECT 17.200 0.180 17.500 0.480 ;
        RECT 17.690 0.180 17.990 0.480 ;
        RECT 19.540 0.180 19.840 0.480 ;
        RECT 20.030 0.180 20.330 0.480 ;
        RECT 20.520 0.180 20.820 0.480 ;
        RECT 22.780 0.180 23.080 0.480 ;
        RECT 23.270 0.180 23.570 0.480 ;
        RECT 23.760 0.180 24.060 0.480 ;
        RECT 24.250 0.180 24.550 0.480 ;
        RECT 24.740 0.180 25.040 0.480 ;
        RECT 25.230 0.180 25.530 0.480 ;
        RECT 25.720 0.180 26.020 0.480 ;
        RECT 26.210 0.180 26.510 0.480 ;
        RECT 28.290 0.180 28.590 0.480 ;
        RECT 28.780 0.180 29.080 0.480 ;
        RECT 29.270 0.180 29.570 0.480 ;
        RECT 29.760 0.180 30.060 0.480 ;
        RECT 30.250 0.180 30.550 0.480 ;
        RECT 30.740 0.180 31.040 0.480 ;
        RECT 31.230 0.180 31.530 0.480 ;
        RECT 31.720 0.180 32.020 0.480 ;
        RECT 33.930 0.180 34.230 0.480 ;
        RECT 34.420 0.180 34.720 0.480 ;
        RECT 34.910 0.180 35.210 0.480 ;
        RECT 35.400 0.180 35.700 0.480 ;
        RECT 37.250 0.180 37.550 0.480 ;
        RECT 37.740 0.180 38.040 0.480 ;
        RECT 38.230 0.180 38.530 0.480 ;
        RECT 40.490 0.180 40.790 0.480 ;
        RECT 40.980 0.180 41.280 0.480 ;
        RECT 41.470 0.180 41.770 0.480 ;
        RECT 41.960 0.180 42.260 0.480 ;
        RECT 42.450 0.180 42.750 0.480 ;
        RECT 42.940 0.180 43.240 0.480 ;
        RECT 43.430 0.180 43.730 0.480 ;
        RECT 43.920 0.180 44.220 0.480 ;
        RECT 46.000 0.180 46.300 0.480 ;
        RECT 46.490 0.180 46.790 0.480 ;
        RECT 46.980 0.180 47.280 0.480 ;
        RECT 47.470 0.180 47.770 0.480 ;
        RECT 47.960 0.180 48.260 0.480 ;
        RECT 48.450 0.180 48.750 0.480 ;
        RECT 48.940 0.180 49.240 0.480 ;
        RECT 49.430 0.180 49.730 0.480 ;
        RECT 51.640 0.180 51.940 0.480 ;
        RECT 52.130 0.180 52.430 0.480 ;
        RECT 52.620 0.180 52.920 0.480 ;
        RECT 53.110 0.180 53.410 0.480 ;
        RECT 54.960 0.180 55.260 0.480 ;
        RECT 55.450 0.180 55.750 0.480 ;
        RECT 55.940 0.180 56.240 0.480 ;
        RECT 58.200 0.180 58.500 0.480 ;
        RECT 58.690 0.180 58.990 0.480 ;
        RECT 59.180 0.180 59.480 0.480 ;
        RECT 59.670 0.180 59.970 0.480 ;
        RECT 60.160 0.180 60.460 0.480 ;
        RECT 60.650 0.180 60.950 0.480 ;
        RECT 61.140 0.180 61.440 0.480 ;
        RECT 61.630 0.180 61.930 0.480 ;
        RECT 63.710 0.180 64.010 0.480 ;
        RECT 64.200 0.180 64.500 0.480 ;
        RECT 64.690 0.180 64.990 0.480 ;
        RECT 65.180 0.180 65.480 0.480 ;
        RECT 65.670 0.180 65.970 0.480 ;
        RECT 66.160 0.180 66.460 0.480 ;
        RECT 66.650 0.180 66.950 0.480 ;
        RECT 67.140 0.180 67.440 0.480 ;
        RECT 69.350 0.180 69.650 0.480 ;
        RECT 69.840 0.180 70.140 0.480 ;
        RECT 70.330 0.180 70.630 0.480 ;
        RECT 70.820 0.180 71.120 0.480 ;
        RECT 72.670 0.180 72.970 0.480 ;
        RECT 73.160 0.180 73.460 0.480 ;
        RECT 73.650 0.180 73.950 0.480 ;
        RECT 75.910 0.180 76.210 0.480 ;
        RECT 76.400 0.180 76.700 0.480 ;
        RECT 76.890 0.180 77.190 0.480 ;
        RECT 77.380 0.180 77.680 0.480 ;
        RECT 77.870 0.180 78.170 0.480 ;
        RECT 78.360 0.180 78.660 0.480 ;
        RECT 78.850 0.180 79.150 0.480 ;
        RECT 79.340 0.180 79.640 0.480 ;
        RECT 81.420 0.180 81.720 0.480 ;
        RECT 81.910 0.180 82.210 0.480 ;
        RECT 82.400 0.180 82.700 0.480 ;
        RECT 82.890 0.180 83.190 0.480 ;
        RECT 83.380 0.180 83.680 0.480 ;
        RECT 83.870 0.180 84.170 0.480 ;
        RECT 84.360 0.180 84.660 0.480 ;
        RECT 84.850 0.180 85.150 0.480 ;
        RECT 87.060 0.180 87.360 0.480 ;
        RECT 87.550 0.180 87.850 0.480 ;
        RECT 88.040 0.180 88.340 0.480 ;
        RECT 88.530 0.180 88.830 0.480 ;
        RECT 90.380 0.180 90.680 0.480 ;
        RECT 90.870 0.180 91.170 0.480 ;
        RECT 91.360 0.180 91.660 0.480 ;
        RECT 93.620 0.180 93.920 0.480 ;
        RECT 94.110 0.180 94.410 0.480 ;
        RECT 94.600 0.180 94.900 0.480 ;
        RECT 95.090 0.180 95.390 0.480 ;
        RECT 95.580 0.180 95.880 0.480 ;
        RECT 96.070 0.180 96.370 0.480 ;
        RECT 96.560 0.180 96.860 0.480 ;
        RECT 97.050 0.180 97.350 0.480 ;
        RECT 99.130 0.180 99.430 0.480 ;
        RECT 99.620 0.180 99.920 0.480 ;
        RECT 100.110 0.180 100.410 0.480 ;
        RECT 100.600 0.180 100.900 0.480 ;
        RECT 101.090 0.180 101.390 0.480 ;
        RECT 101.580 0.180 101.880 0.480 ;
        RECT 102.070 0.180 102.370 0.480 ;
        RECT 102.560 0.180 102.860 0.480 ;
        RECT 104.770 0.180 105.070 0.480 ;
        RECT 105.260 0.180 105.560 0.480 ;
        RECT 105.750 0.180 106.050 0.480 ;
        RECT 106.240 0.180 106.540 0.480 ;
      LAYER met1 ;
        RECT 8.400 29.270 97.550 29.750 ;
        RECT -1.000 25.280 4.565 25.760 ;
        RECT -7.950 23.950 -7.550 24.350 ;
        RECT 2.180 24.010 10.340 24.310 ;
        RECT 5.760 23.950 10.340 24.010 ;
        RECT 11.295 23.950 28.050 24.310 ;
        RECT 29.005 23.950 45.760 24.310 ;
        RECT 46.715 23.950 63.470 24.310 ;
        RECT 64.425 23.950 81.180 24.310 ;
        RECT 82.135 23.950 100.220 24.310 ;
        RECT 101.000 24.015 103.005 24.380 ;
        RECT -1.000 22.560 4.565 23.040 ;
        RECT 5.760 17.360 6.120 23.950 ;
        RECT 9.980 22.950 10.340 23.950 ;
        RECT 20.960 22.950 21.320 23.950 ;
        RECT 27.690 22.950 28.050 23.950 ;
        RECT 38.670 22.950 39.030 23.950 ;
        RECT 45.400 22.950 45.760 23.950 ;
        RECT 56.380 22.950 56.740 23.950 ;
        RECT 63.110 22.950 63.470 23.950 ;
        RECT 74.090 22.950 74.450 23.950 ;
        RECT 80.820 22.950 81.180 23.950 ;
        RECT 91.800 22.950 92.160 23.950 ;
        RECT 9.370 22.590 13.640 22.950 ;
        RECT 14.890 22.590 19.160 22.950 ;
        RECT 20.410 22.590 21.910 22.950 ;
        RECT 23.740 22.590 25.240 22.950 ;
        RECT 27.080 22.590 31.350 22.950 ;
        RECT 32.600 22.590 36.870 22.950 ;
        RECT 38.120 22.590 39.620 22.950 ;
        RECT 41.450 22.590 42.950 22.950 ;
        RECT 44.790 22.590 49.060 22.950 ;
        RECT 50.310 22.590 54.580 22.950 ;
        RECT 55.830 22.590 57.330 22.950 ;
        RECT 59.160 22.590 60.660 22.950 ;
        RECT 62.500 22.590 66.770 22.950 ;
        RECT 68.020 22.590 72.290 22.950 ;
        RECT 73.540 22.590 75.040 22.950 ;
        RECT 76.870 22.590 78.370 22.950 ;
        RECT 80.210 22.590 84.480 22.950 ;
        RECT 85.730 22.590 90.000 22.950 ;
        RECT 91.250 22.590 92.750 22.950 ;
        RECT 94.580 22.590 96.080 22.950 ;
        RECT 15.505 21.590 15.865 22.590 ;
        RECT 24.290 21.590 24.650 22.590 ;
        RECT 33.215 21.590 33.575 22.590 ;
        RECT 42.000 21.590 42.360 22.590 ;
        RECT 50.925 21.590 51.285 22.590 ;
        RECT 59.710 21.590 60.070 22.590 ;
        RECT 68.635 21.590 68.995 22.590 ;
        RECT 77.420 21.590 77.780 22.590 ;
        RECT 86.345 21.590 86.705 22.590 ;
        RECT 95.130 21.590 95.490 22.590 ;
        RECT -2.510 17.000 6.120 17.360 ;
        RECT 7.120 21.230 15.865 21.590 ;
        RECT 16.815 21.230 33.575 21.590 ;
        RECT 34.525 21.230 51.285 21.590 ;
        RECT 52.235 21.230 68.995 21.590 ;
        RECT 69.945 21.230 86.705 21.590 ;
        RECT 87.655 21.230 98.860 21.590 ;
        RECT -2.510 5.890 -2.150 17.000 ;
        RECT 7.120 16.000 7.480 21.230 ;
        RECT -1.150 15.640 7.480 16.000 ;
        RECT 8.480 15.670 97.550 16.150 ;
        RECT 98.500 16.000 98.860 21.230 ;
        RECT 99.860 17.360 100.220 23.950 ;
        RECT 102.000 18.500 103.000 19.515 ;
        RECT 107.515 18.500 108.500 19.500 ;
        RECT 99.860 17.000 109.360 17.360 ;
        RECT 98.500 15.640 108.000 16.000 ;
        RECT -1.150 8.610 -0.790 15.640 ;
        RECT 0.000 13.690 106.780 14.170 ;
        RECT 107.640 8.610 108.000 15.640 ;
        RECT -1.150 8.250 9.895 8.610 ;
        RECT 10.845 8.250 27.605 8.610 ;
        RECT 28.555 8.250 45.315 8.610 ;
        RECT 46.265 8.250 63.025 8.610 ;
        RECT 63.975 8.250 80.735 8.610 ;
        RECT 81.685 8.250 98.445 8.610 ;
        RECT 99.395 8.250 108.000 8.610 ;
        RECT 2.060 7.250 2.420 8.250 ;
        RECT 10.845 7.250 11.205 8.250 ;
        RECT 19.770 7.250 20.130 8.250 ;
        RECT 28.555 7.250 28.915 8.250 ;
        RECT 37.480 7.250 37.840 8.250 ;
        RECT 46.265 7.250 46.625 8.250 ;
        RECT 55.190 7.250 55.550 8.250 ;
        RECT 63.975 7.250 64.335 8.250 ;
        RECT 72.900 7.250 73.260 8.250 ;
        RECT 81.685 7.250 82.045 8.250 ;
        RECT 90.610 7.250 90.970 8.250 ;
        RECT 99.395 7.250 99.755 8.250 ;
        RECT 1.470 6.890 2.970 7.250 ;
        RECT 4.800 6.890 6.300 7.250 ;
        RECT 7.550 6.890 11.820 7.250 ;
        RECT 13.070 6.890 17.340 7.250 ;
        RECT 19.180 6.890 20.680 7.250 ;
        RECT 22.510 6.890 24.010 7.250 ;
        RECT 25.260 6.890 29.530 7.250 ;
        RECT 30.780 6.890 35.050 7.250 ;
        RECT 36.890 6.890 38.390 7.250 ;
        RECT 40.220 6.890 41.720 7.250 ;
        RECT 42.970 6.890 47.240 7.250 ;
        RECT 48.490 6.890 52.760 7.250 ;
        RECT 54.600 6.890 56.100 7.250 ;
        RECT 57.930 6.890 59.430 7.250 ;
        RECT 60.680 6.890 64.950 7.250 ;
        RECT 66.200 6.890 70.470 7.250 ;
        RECT 72.310 6.890 73.810 7.250 ;
        RECT 75.640 6.890 77.140 7.250 ;
        RECT 78.390 6.890 82.660 7.250 ;
        RECT 83.910 6.890 88.180 7.250 ;
        RECT 90.020 6.890 91.520 7.250 ;
        RECT 93.350 6.890 94.850 7.250 ;
        RECT 96.100 6.890 100.370 7.250 ;
        RECT 101.620 6.890 105.890 7.250 ;
        RECT 5.390 5.890 5.750 6.890 ;
        RECT 16.370 5.890 16.730 6.890 ;
        RECT 23.100 5.890 23.460 6.890 ;
        RECT 34.080 5.890 34.440 6.890 ;
        RECT 40.810 5.890 41.170 6.890 ;
        RECT 51.790 5.890 52.150 6.890 ;
        RECT 58.520 5.890 58.880 6.890 ;
        RECT 69.500 5.890 69.860 6.890 ;
        RECT 76.230 5.890 76.590 6.890 ;
        RECT 87.210 5.890 87.570 6.890 ;
        RECT 93.940 5.890 94.300 6.890 ;
        RECT 104.920 5.890 105.280 6.890 ;
        RECT 109.000 5.890 109.360 17.000 ;
        RECT -2.510 5.530 15.415 5.890 ;
        RECT 16.370 5.530 33.125 5.890 ;
        RECT 34.080 5.530 50.835 5.890 ;
        RECT 51.790 5.530 68.545 5.890 ;
        RECT 69.500 5.530 86.255 5.890 ;
        RECT 87.210 5.530 103.965 5.890 ;
        RECT 104.920 5.530 109.360 5.890 ;
        RECT 0.000 0.090 106.780 0.570 ;
      LAYER via ;
        RECT 19.610 23.950 19.970 24.310 ;
        RECT 43.980 23.950 44.340 24.310 ;
        RECT 60.770 23.950 61.130 24.310 ;
        RECT 76.070 23.950 76.430 24.310 ;
        RECT 98.500 23.950 98.860 24.310 ;
        RECT 12.000 15.770 12.260 16.030 ;
        RECT 12.370 15.770 12.630 16.030 ;
        RECT 12.740 15.770 13.000 16.030 ;
        RECT 18.000 15.770 18.260 16.030 ;
        RECT 18.370 15.770 18.630 16.030 ;
        RECT 18.740 15.770 19.000 16.030 ;
        RECT 24.000 15.770 24.260 16.030 ;
        RECT 24.370 15.770 24.630 16.030 ;
        RECT 24.740 15.770 25.000 16.030 ;
        RECT 30.000 15.770 30.260 16.030 ;
        RECT 30.370 15.770 30.630 16.030 ;
        RECT 30.740 15.770 31.000 16.030 ;
        RECT 36.000 15.770 36.260 16.030 ;
        RECT 36.370 15.770 36.630 16.030 ;
        RECT 36.740 15.770 37.000 16.030 ;
        RECT 42.000 15.770 42.260 16.030 ;
        RECT 42.370 15.770 42.630 16.030 ;
        RECT 42.740 15.770 43.000 16.030 ;
        RECT 48.000 15.770 48.260 16.030 ;
        RECT 48.370 15.770 48.630 16.030 ;
        RECT 48.740 15.770 49.000 16.030 ;
        RECT 54.000 15.770 54.260 16.030 ;
        RECT 54.370 15.770 54.630 16.030 ;
        RECT 54.740 15.770 55.000 16.030 ;
        RECT 60.000 15.770 60.260 16.030 ;
        RECT 60.370 15.770 60.630 16.030 ;
        RECT 60.740 15.770 61.000 16.030 ;
        RECT 66.000 15.770 66.260 16.030 ;
        RECT 66.370 15.770 66.630 16.030 ;
        RECT 66.740 15.770 67.000 16.030 ;
        RECT 72.000 15.770 72.260 16.030 ;
        RECT 72.370 15.770 72.630 16.030 ;
        RECT 72.740 15.770 73.000 16.030 ;
        RECT 78.000 15.770 78.260 16.030 ;
        RECT 78.370 15.770 78.630 16.030 ;
        RECT 78.740 15.770 79.000 16.030 ;
        RECT 84.000 15.770 84.260 16.030 ;
        RECT 84.370 15.770 84.630 16.030 ;
        RECT 84.740 15.770 85.000 16.030 ;
        RECT 90.000 15.770 90.260 16.030 ;
        RECT 90.370 15.770 90.630 16.030 ;
        RECT 90.740 15.770 91.000 16.030 ;
        RECT 96.000 15.770 96.260 16.030 ;
        RECT 96.370 15.770 96.630 16.030 ;
        RECT 96.740 15.770 97.000 16.030 ;
        RECT 102.070 19.100 102.410 19.440 ;
        RECT 102.590 19.100 102.930 19.440 ;
        RECT 102.070 18.580 102.410 18.920 ;
        RECT 102.590 18.580 102.930 18.920 ;
        RECT 107.585 19.080 107.925 19.420 ;
        RECT 108.075 19.080 108.415 19.420 ;
        RECT 107.585 18.580 107.925 18.920 ;
        RECT 108.075 18.580 108.415 18.920 ;
        RECT 0.000 13.790 0.260 14.050 ;
        RECT 0.370 13.790 0.630 14.050 ;
        RECT 0.740 13.790 1.000 14.050 ;
        RECT 6.000 13.790 6.260 14.050 ;
        RECT 6.370 13.790 6.630 14.050 ;
        RECT 6.740 13.790 7.000 14.050 ;
        RECT 12.000 13.790 12.260 14.050 ;
        RECT 12.370 13.790 12.630 14.050 ;
        RECT 12.740 13.790 13.000 14.050 ;
        RECT 18.000 13.790 18.260 14.050 ;
        RECT 18.370 13.790 18.630 14.050 ;
        RECT 18.740 13.790 19.000 14.050 ;
        RECT 24.000 13.790 24.260 14.050 ;
        RECT 24.370 13.790 24.630 14.050 ;
        RECT 24.740 13.790 25.000 14.050 ;
        RECT 30.000 13.790 30.260 14.050 ;
        RECT 30.370 13.790 30.630 14.050 ;
        RECT 30.740 13.790 31.000 14.050 ;
        RECT 36.000 13.790 36.260 14.050 ;
        RECT 36.370 13.790 36.630 14.050 ;
        RECT 36.740 13.790 37.000 14.050 ;
        RECT 42.000 13.790 42.260 14.050 ;
        RECT 42.370 13.790 42.630 14.050 ;
        RECT 42.740 13.790 43.000 14.050 ;
        RECT 48.000 13.790 48.260 14.050 ;
        RECT 48.370 13.790 48.630 14.050 ;
        RECT 48.740 13.790 49.000 14.050 ;
        RECT 54.000 13.790 54.260 14.050 ;
        RECT 54.370 13.790 54.630 14.050 ;
        RECT 54.740 13.790 55.000 14.050 ;
        RECT 60.000 13.790 60.260 14.050 ;
        RECT 60.370 13.790 60.630 14.050 ;
        RECT 60.740 13.790 61.000 14.050 ;
        RECT 66.000 13.790 66.260 14.050 ;
        RECT 66.370 13.790 66.630 14.050 ;
        RECT 66.740 13.790 67.000 14.050 ;
        RECT 72.000 13.790 72.260 14.050 ;
        RECT 72.370 13.790 72.630 14.050 ;
        RECT 72.740 13.790 73.000 14.050 ;
        RECT 78.000 13.790 78.260 14.050 ;
        RECT 78.370 13.790 78.630 14.050 ;
        RECT 78.740 13.790 79.000 14.050 ;
        RECT 84.000 13.790 84.260 14.050 ;
        RECT 84.370 13.790 84.630 14.050 ;
        RECT 84.740 13.790 85.000 14.050 ;
        RECT 90.000 13.790 90.260 14.050 ;
        RECT 90.370 13.790 90.630 14.050 ;
        RECT 90.740 13.790 91.000 14.050 ;
        RECT 96.000 13.790 96.260 14.050 ;
        RECT 96.370 13.790 96.630 14.050 ;
        RECT 96.740 13.790 97.000 14.050 ;
        RECT 102.000 13.790 102.260 14.050 ;
        RECT 102.370 13.790 102.630 14.050 ;
        RECT 102.740 13.790 103.000 14.050 ;
        RECT 105.780 13.790 106.040 14.050 ;
        RECT 106.150 13.790 106.410 14.050 ;
        RECT 106.520 13.790 106.780 14.050 ;
        RECT -0.360 5.530 0.000 5.890 ;
        RECT 17.780 5.530 18.140 5.890 ;
        RECT 35.530 5.530 35.890 5.890 ;
        RECT 58.520 5.530 58.880 5.890 ;
        RECT 71.840 5.530 72.200 5.890 ;
        RECT 88.640 5.530 89.000 5.890 ;
      LAYER met2 ;
        RECT 19.580 23.950 20.000 31.500 ;
        RECT 43.950 23.950 44.370 31.500 ;
        RECT 60.740 23.950 61.160 31.500 ;
        RECT 76.040 23.950 76.460 31.500 ;
        RECT 98.470 23.950 98.890 31.500 ;
        RECT 102.000 18.500 103.000 19.515 ;
        RECT 107.515 19.000 115.600 19.500 ;
        RECT 107.515 18.500 108.500 19.000 ;
        RECT 12.000 15.700 13.000 16.100 ;
        RECT 18.000 15.700 19.000 16.100 ;
        RECT 24.000 15.700 25.000 16.100 ;
        RECT 30.000 15.700 31.000 16.100 ;
        RECT 36.000 15.700 37.000 16.100 ;
        RECT 42.000 15.700 43.000 16.100 ;
        RECT 48.000 15.700 49.000 16.100 ;
        RECT 54.000 15.700 55.000 16.100 ;
        RECT 60.000 15.700 61.000 16.100 ;
        RECT 66.000 15.700 67.000 16.100 ;
        RECT 72.000 15.700 73.000 16.100 ;
        RECT 78.000 15.700 79.000 16.100 ;
        RECT 84.000 15.700 85.000 16.100 ;
        RECT 90.000 15.700 91.000 16.100 ;
        RECT 96.000 15.700 97.000 16.100 ;
        RECT 0.000 13.720 1.000 14.120 ;
        RECT 6.000 13.720 7.000 14.120 ;
        RECT 12.000 13.720 13.000 14.120 ;
        RECT 18.000 13.720 19.000 14.120 ;
        RECT 24.000 13.720 25.000 14.120 ;
        RECT 30.000 13.720 31.000 14.120 ;
        RECT 36.000 13.720 37.000 14.120 ;
        RECT 42.000 13.720 43.000 14.120 ;
        RECT 48.000 13.720 49.000 14.120 ;
        RECT 54.000 13.720 55.000 14.120 ;
        RECT 60.000 13.720 61.000 14.120 ;
        RECT 66.000 13.720 67.000 14.120 ;
        RECT 72.000 13.720 73.000 14.120 ;
        RECT 78.000 13.720 79.000 14.120 ;
        RECT 84.000 13.720 85.000 14.120 ;
        RECT 90.000 13.720 91.000 14.120 ;
        RECT 96.000 13.720 97.000 14.120 ;
        RECT 102.000 13.720 103.000 14.120 ;
        RECT 105.780 13.720 106.780 14.120 ;
        RECT -0.390 -1.720 0.030 5.890 ;
        RECT 17.750 -1.720 18.170 5.890 ;
        RECT 35.500 -1.720 35.920 5.890 ;
        RECT 58.490 -1.720 58.910 5.890 ;
        RECT 71.810 -1.720 72.230 5.890 ;
        RECT 88.610 -1.720 89.030 5.890 ;
      LAYER via2 ;
        RECT 102.040 19.070 102.440 19.470 ;
        RECT 102.560 19.070 102.960 19.470 ;
        RECT 102.040 18.550 102.440 18.950 ;
        RECT 102.560 18.550 102.960 18.950 ;
        RECT 12.100 15.750 12.400 16.050 ;
        RECT 12.600 15.750 12.900 16.050 ;
        RECT 18.100 15.750 18.400 16.050 ;
        RECT 18.600 15.750 18.900 16.050 ;
        RECT 24.100 15.750 24.400 16.050 ;
        RECT 24.600 15.750 24.900 16.050 ;
        RECT 30.100 15.750 30.400 16.050 ;
        RECT 30.600 15.750 30.900 16.050 ;
        RECT 36.100 15.750 36.400 16.050 ;
        RECT 36.600 15.750 36.900 16.050 ;
        RECT 42.100 15.750 42.400 16.050 ;
        RECT 42.600 15.750 42.900 16.050 ;
        RECT 48.100 15.750 48.400 16.050 ;
        RECT 48.600 15.750 48.900 16.050 ;
        RECT 54.100 15.750 54.400 16.050 ;
        RECT 54.600 15.750 54.900 16.050 ;
        RECT 60.100 15.750 60.400 16.050 ;
        RECT 60.600 15.750 60.900 16.050 ;
        RECT 66.100 15.750 66.400 16.050 ;
        RECT 66.600 15.750 66.900 16.050 ;
        RECT 72.100 15.750 72.400 16.050 ;
        RECT 72.600 15.750 72.900 16.050 ;
        RECT 78.100 15.750 78.400 16.050 ;
        RECT 78.600 15.750 78.900 16.050 ;
        RECT 84.100 15.750 84.400 16.050 ;
        RECT 84.600 15.750 84.900 16.050 ;
        RECT 90.100 15.750 90.400 16.050 ;
        RECT 90.600 15.750 90.900 16.050 ;
        RECT 96.100 15.750 96.400 16.050 ;
        RECT 96.600 15.750 96.900 16.050 ;
        RECT 0.100 13.770 0.400 14.070 ;
        RECT 0.600 13.770 0.900 14.070 ;
        RECT 6.100 13.770 6.400 14.070 ;
        RECT 6.600 13.770 6.900 14.070 ;
        RECT 12.100 13.770 12.400 14.070 ;
        RECT 12.600 13.770 12.900 14.070 ;
        RECT 18.100 13.770 18.400 14.070 ;
        RECT 18.600 13.770 18.900 14.070 ;
        RECT 24.100 13.770 24.400 14.070 ;
        RECT 24.600 13.770 24.900 14.070 ;
        RECT 30.100 13.770 30.400 14.070 ;
        RECT 30.600 13.770 30.900 14.070 ;
        RECT 36.100 13.770 36.400 14.070 ;
        RECT 36.600 13.770 36.900 14.070 ;
        RECT 42.100 13.770 42.400 14.070 ;
        RECT 42.600 13.770 42.900 14.070 ;
        RECT 48.100 13.770 48.400 14.070 ;
        RECT 48.600 13.770 48.900 14.070 ;
        RECT 54.100 13.770 54.400 14.070 ;
        RECT 54.600 13.770 54.900 14.070 ;
        RECT 60.100 13.770 60.400 14.070 ;
        RECT 60.600 13.770 60.900 14.070 ;
        RECT 66.100 13.770 66.400 14.070 ;
        RECT 66.600 13.770 66.900 14.070 ;
        RECT 72.100 13.770 72.400 14.070 ;
        RECT 72.600 13.770 72.900 14.070 ;
        RECT 78.100 13.770 78.400 14.070 ;
        RECT 78.600 13.770 78.900 14.070 ;
        RECT 84.100 13.770 84.400 14.070 ;
        RECT 84.600 13.770 84.900 14.070 ;
        RECT 90.100 13.770 90.400 14.070 ;
        RECT 90.600 13.770 90.900 14.070 ;
        RECT 96.100 13.770 96.400 14.070 ;
        RECT 96.600 13.770 96.900 14.070 ;
        RECT 102.100 13.770 102.400 14.070 ;
        RECT 102.600 13.770 102.900 14.070 ;
        RECT 105.880 13.770 106.180 14.070 ;
        RECT 106.380 13.770 106.680 14.070 ;
      LAYER met3 ;
        RECT 12.000 15.670 13.000 16.150 ;
        RECT 18.000 15.670 19.000 16.150 ;
        RECT 24.000 15.670 25.000 16.150 ;
        RECT 30.000 15.670 31.000 16.150 ;
        RECT 36.000 15.670 37.000 16.150 ;
        RECT 42.000 15.670 43.000 16.150 ;
        RECT 48.000 15.670 49.000 16.150 ;
        RECT 54.000 15.670 55.000 16.150 ;
        RECT 60.000 15.670 61.000 16.150 ;
        RECT 66.000 15.670 67.000 16.150 ;
        RECT 72.000 15.670 73.000 16.150 ;
        RECT 78.000 15.670 79.000 16.150 ;
        RECT 84.000 15.670 85.000 16.150 ;
        RECT 90.000 15.670 91.000 16.150 ;
        RECT 96.000 15.670 97.000 16.150 ;
        RECT 102.000 15.670 103.000 19.515 ;
        RECT 0.000 14.170 106.780 15.670 ;
        RECT 0.000 13.690 1.000 14.170 ;
        RECT 6.000 13.690 7.000 14.170 ;
        RECT 12.000 13.690 13.000 14.170 ;
        RECT 18.000 13.690 19.000 14.170 ;
        RECT 24.000 13.690 25.000 14.170 ;
        RECT 30.000 13.690 31.000 14.170 ;
        RECT 36.000 13.690 37.000 14.170 ;
        RECT 42.000 13.690 43.000 14.170 ;
        RECT 48.000 13.690 49.000 14.170 ;
        RECT 54.000 13.690 55.000 14.170 ;
        RECT 60.000 13.690 61.000 14.170 ;
        RECT 66.000 13.690 67.000 14.170 ;
        RECT 72.000 13.690 73.000 14.170 ;
        RECT 78.000 13.690 79.000 14.170 ;
        RECT 84.000 13.690 85.000 14.170 ;
        RECT 90.000 13.690 91.000 14.170 ;
        RECT 96.000 13.690 97.000 14.170 ;
        RECT 102.000 13.690 103.000 14.170 ;
        RECT 105.780 13.690 106.780 14.170 ;
  END
END ring_osc
MACRO pwell_co_ring
  CLASS BLOCK ;
  FOREIGN pwell_co_ring ;
  ORIGIN 8.400 31.800 ;
  SIZE 109.125 BY 32.100 ;
  OBS
      LAYER li1 ;
        RECT -0.100 0.000 90.900 0.300 ;
        RECT -0.100 -15.630 0.200 0.000 ;
        RECT 90.600 -15.630 90.900 0.000 ;
        RECT -8.400 -15.930 100.725 -15.630 ;
        RECT -8.400 -31.500 -8.100 -15.930 ;
        RECT 100.400 -16.000 100.725 -15.930 ;
        RECT 100.400 -31.500 100.700 -16.000 ;
        RECT -8.400 -31.800 100.700 -31.500 ;
  END
END pwell_co_ring
MACRO via_m4_li
  CLASS BLOCK ;
  FOREIGN via_m4_li ;
  ORIGIN 0.000 -0.010 ;
  SIZE 2.000 BY 0.480 ;
  OBS
      LAYER li1 ;
        RECT 0.000 0.100 2.000 0.400 ;
      LAYER mcon ;
        RECT 0.110 0.100 0.410 0.400 ;
        RECT 0.600 0.100 0.900 0.400 ;
        RECT 1.100 0.100 1.400 0.400 ;
        RECT 1.590 0.100 1.890 0.400 ;
      LAYER met1 ;
        RECT 0.080 0.010 1.920 0.490 ;
      LAYER via ;
        RECT 0.130 0.100 0.430 0.400 ;
        RECT 0.490 0.100 0.790 0.400 ;
        RECT 0.850 0.100 1.150 0.400 ;
        RECT 1.210 0.100 1.510 0.400 ;
        RECT 1.570 0.100 1.870 0.400 ;
      LAYER met2 ;
        RECT 0.000 0.010 2.000 0.490 ;
      LAYER via2 ;
        RECT 0.180 0.090 0.500 0.410 ;
        RECT 0.620 0.090 0.940 0.410 ;
        RECT 1.060 0.090 1.380 0.410 ;
        RECT 1.500 0.090 1.820 0.410 ;
      LAYER met3 ;
        RECT 0.000 0.010 2.000 0.490 ;
      LAYER via3 ;
        RECT 0.160 0.070 0.520 0.435 ;
        RECT 0.600 0.070 0.960 0.435 ;
        RECT 1.040 0.070 1.400 0.435 ;
        RECT 1.480 0.070 1.840 0.435 ;
      LAYER met4 ;
        RECT 0.000 0.010 2.000 0.490 ;
  END
END via_m4_li
MACRO via_m1
  CLASS BLOCK ;
  FOREIGN via_m1 ;
  ORIGIN -54.490 -34.780 ;
  SIZE 2.000 BY 0.480 ;
  OBS
      LAYER met1 ;
        RECT 54.620 34.780 56.360 35.260 ;
      LAYER via ;
        RECT 54.620 34.870 54.920 35.170 ;
        RECT 54.980 34.870 55.280 35.170 ;
        RECT 55.340 34.870 55.640 35.170 ;
        RECT 55.700 34.870 56.000 35.170 ;
        RECT 56.060 34.870 56.360 35.170 ;
      LAYER met2 ;
        RECT 54.490 34.780 56.490 35.260 ;
      LAYER via2 ;
        RECT 54.670 34.860 54.990 35.180 ;
        RECT 55.110 34.860 55.430 35.180 ;
        RECT 55.550 34.860 55.870 35.180 ;
        RECT 55.990 34.860 56.310 35.180 ;
      LAYER met3 ;
        RECT 54.490 34.780 56.490 35.260 ;
      LAYER via3 ;
        RECT 54.650 34.840 55.010 35.205 ;
        RECT 55.090 34.840 55.450 35.205 ;
        RECT 55.530 34.840 55.890 35.205 ;
        RECT 55.970 34.840 56.330 35.205 ;
      LAYER met4 ;
        RECT 54.490 34.780 56.490 35.260 ;
  END
END via_m1
MACRO vco_w6_r100
  CLASS BLOCK ;
  FOREIGN vco_w6_r100 ;
  ORIGIN 0.450 12.000 ;
  SIZE 123.550 BY 105.000 ;
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 92.420 33.250 92.800 33.300 ;
        RECT 91.470 32.890 92.800 33.250 ;
        RECT 92.420 32.840 92.800 32.890 ;
        RECT 94.290 33.250 94.670 33.300 ;
        RECT 94.290 32.890 95.620 33.250 ;
        RECT 94.290 32.840 94.670 32.890 ;
        RECT 96.730 26.750 97.030 39.340 ;
        RECT 100.960 33.250 101.340 33.300 ;
        RECT 100.960 32.890 102.290 33.250 ;
        RECT 100.960 32.840 101.340 32.890 ;
        RECT 111.105 26.750 111.405 39.340 ;
      LAYER mcon ;
        RECT 91.470 32.920 91.770 33.220 ;
        RECT 91.960 32.920 92.260 33.220 ;
        RECT 92.450 32.920 92.750 33.220 ;
        RECT 94.340 32.920 94.640 33.220 ;
        RECT 94.830 32.920 95.130 33.220 ;
        RECT 95.320 32.920 95.620 33.220 ;
        RECT 101.010 32.920 101.310 33.220 ;
        RECT 101.500 32.920 101.800 33.220 ;
        RECT 101.990 32.920 102.290 33.220 ;
        RECT 96.730 31.560 97.030 31.860 ;
        RECT 111.105 31.560 111.405 31.860 ;
      LAYER met1 ;
        RECT 91.410 32.890 95.680 33.250 ;
        RECT 100.850 32.890 102.350 33.250 ;
        RECT 94.710 31.890 95.070 32.890 ;
        RECT 101.440 31.890 101.800 32.890 ;
        RECT 94.710 31.530 111.465 31.890 ;
      LAYER via ;
        RECT 96.140 31.530 96.500 31.890 ;
      LAYER met2 ;
        RECT 96.110 24.280 96.530 31.890 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 74.710 33.250 75.090 33.300 ;
        RECT 73.760 32.890 75.090 33.250 ;
        RECT 74.710 32.840 75.090 32.890 ;
        RECT 76.580 33.250 76.960 33.300 ;
        RECT 76.580 32.890 77.910 33.250 ;
        RECT 76.580 32.840 76.960 32.890 ;
        RECT 79.020 26.750 79.320 39.340 ;
        RECT 83.250 33.250 83.630 33.300 ;
        RECT 83.250 32.890 84.580 33.250 ;
        RECT 83.250 32.840 83.630 32.890 ;
        RECT 93.395 26.750 93.695 39.340 ;
      LAYER mcon ;
        RECT 73.760 32.920 74.060 33.220 ;
        RECT 74.250 32.920 74.550 33.220 ;
        RECT 74.740 32.920 75.040 33.220 ;
        RECT 76.630 32.920 76.930 33.220 ;
        RECT 77.120 32.920 77.420 33.220 ;
        RECT 77.610 32.920 77.910 33.220 ;
        RECT 83.300 32.920 83.600 33.220 ;
        RECT 83.790 32.920 84.090 33.220 ;
        RECT 84.280 32.920 84.580 33.220 ;
        RECT 79.020 31.560 79.320 31.860 ;
        RECT 93.395 31.560 93.695 31.860 ;
      LAYER met1 ;
        RECT 73.700 32.890 77.970 33.250 ;
        RECT 83.140 32.890 84.640 33.250 ;
        RECT 77.000 31.890 77.360 32.890 ;
        RECT 83.730 31.890 84.090 32.890 ;
        RECT 77.000 31.530 93.755 31.890 ;
      LAYER via ;
        RECT 79.340 31.530 79.700 31.890 ;
      LAYER met2 ;
        RECT 79.310 24.280 79.730 31.890 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 57.000 33.250 57.380 33.300 ;
        RECT 56.050 32.890 57.380 33.250 ;
        RECT 57.000 32.840 57.380 32.890 ;
        RECT 58.870 33.250 59.250 33.300 ;
        RECT 58.870 32.890 60.200 33.250 ;
        RECT 58.870 32.840 59.250 32.890 ;
        RECT 61.310 26.750 61.610 39.340 ;
        RECT 65.540 33.250 65.920 33.300 ;
        RECT 65.540 32.890 66.870 33.250 ;
        RECT 65.540 32.840 65.920 32.890 ;
        RECT 75.685 26.750 75.985 39.340 ;
      LAYER mcon ;
        RECT 56.050 32.920 56.350 33.220 ;
        RECT 56.540 32.920 56.840 33.220 ;
        RECT 57.030 32.920 57.330 33.220 ;
        RECT 58.920 32.920 59.220 33.220 ;
        RECT 59.410 32.920 59.710 33.220 ;
        RECT 59.900 32.920 60.200 33.220 ;
        RECT 65.590 32.920 65.890 33.220 ;
        RECT 66.080 32.920 66.380 33.220 ;
        RECT 66.570 32.920 66.870 33.220 ;
        RECT 61.310 31.560 61.610 31.860 ;
        RECT 75.685 31.560 75.985 31.860 ;
      LAYER met1 ;
        RECT 55.990 32.890 60.260 33.250 ;
        RECT 65.430 32.890 66.930 33.250 ;
        RECT 59.290 31.890 59.650 32.890 ;
        RECT 66.020 31.890 66.380 32.890 ;
        RECT 59.290 31.530 76.045 31.890 ;
      LAYER via ;
        RECT 66.020 31.530 66.380 31.890 ;
      LAYER met2 ;
        RECT 65.990 24.280 66.410 31.890 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 39.290 33.250 39.670 33.300 ;
        RECT 38.340 32.890 39.670 33.250 ;
        RECT 39.290 32.840 39.670 32.890 ;
        RECT 41.160 33.250 41.540 33.300 ;
        RECT 41.160 32.890 42.490 33.250 ;
        RECT 41.160 32.840 41.540 32.890 ;
        RECT 43.600 26.750 43.900 39.340 ;
        RECT 47.830 33.250 48.210 33.300 ;
        RECT 47.830 32.890 49.160 33.250 ;
        RECT 47.830 32.840 48.210 32.890 ;
        RECT 57.975 26.750 58.275 39.340 ;
      LAYER mcon ;
        RECT 38.340 32.920 38.640 33.220 ;
        RECT 38.830 32.920 39.130 33.220 ;
        RECT 39.320 32.920 39.620 33.220 ;
        RECT 41.210 32.920 41.510 33.220 ;
        RECT 41.700 32.920 42.000 33.220 ;
        RECT 42.190 32.920 42.490 33.220 ;
        RECT 47.880 32.920 48.180 33.220 ;
        RECT 48.370 32.920 48.670 33.220 ;
        RECT 48.860 32.920 49.160 33.220 ;
        RECT 43.600 31.560 43.900 31.860 ;
        RECT 57.975 31.560 58.275 31.860 ;
      LAYER met1 ;
        RECT 38.280 32.890 42.550 33.250 ;
        RECT 47.720 32.890 49.220 33.250 ;
        RECT 41.580 31.890 41.940 32.890 ;
        RECT 48.310 31.890 48.670 32.890 ;
        RECT 41.580 31.530 58.335 31.890 ;
      LAYER via ;
        RECT 43.030 31.530 43.390 31.890 ;
      LAYER met2 ;
        RECT 43.000 24.280 43.420 31.890 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 21.580 33.250 21.960 33.300 ;
        RECT 20.630 32.890 21.960 33.250 ;
        RECT 21.580 32.840 21.960 32.890 ;
        RECT 23.450 33.250 23.830 33.300 ;
        RECT 23.450 32.890 24.780 33.250 ;
        RECT 23.450 32.840 23.830 32.890 ;
        RECT 25.890 26.750 26.190 39.340 ;
        RECT 30.120 33.250 30.500 33.300 ;
        RECT 30.120 32.890 31.450 33.250 ;
        RECT 30.120 32.840 30.500 32.890 ;
        RECT 40.265 26.750 40.565 39.340 ;
      LAYER mcon ;
        RECT 20.630 32.920 20.930 33.220 ;
        RECT 21.120 32.920 21.420 33.220 ;
        RECT 21.610 32.920 21.910 33.220 ;
        RECT 23.500 32.920 23.800 33.220 ;
        RECT 23.990 32.920 24.290 33.220 ;
        RECT 24.480 32.920 24.780 33.220 ;
        RECT 30.170 32.920 30.470 33.220 ;
        RECT 30.660 32.920 30.960 33.220 ;
        RECT 31.150 32.920 31.450 33.220 ;
        RECT 25.890 31.560 26.190 31.860 ;
        RECT 40.265 31.560 40.565 31.860 ;
      LAYER met1 ;
        RECT 20.570 32.890 24.840 33.250 ;
        RECT 30.010 32.890 31.510 33.250 ;
        RECT 23.870 31.890 24.230 32.890 ;
        RECT 30.600 31.890 30.960 32.890 ;
        RECT 23.870 31.530 40.625 31.890 ;
      LAYER via ;
        RECT 25.280 31.530 25.640 31.890 ;
      LAYER met2 ;
        RECT 25.250 24.280 25.670 31.890 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 6.245500 ;
    PORT
      LAYER li1 ;
        RECT 8.310 50.925 8.905 51.265 ;
        RECT 8.310 49.605 8.485 50.925 ;
        RECT 8.310 49.480 8.905 49.605 ;
        RECT 9.710 49.480 10.010 50.310 ;
        RECT 8.310 49.180 10.010 49.480 ;
        RECT 8.310 49.055 8.905 49.180 ;
        RECT 17.880 48.950 18.260 49.000 ;
        RECT 16.930 48.590 18.260 48.950 ;
        RECT 17.880 48.540 18.260 48.590 ;
        RECT 19.750 48.950 20.130 49.000 ;
        RECT 19.750 48.590 21.080 48.950 ;
        RECT 19.750 48.540 20.130 48.590 ;
        RECT 8.180 26.750 8.480 39.340 ;
        RECT 12.410 33.250 12.790 33.300 ;
        RECT 12.410 32.890 13.740 33.250 ;
        RECT 12.410 32.840 12.790 32.890 ;
        RECT 22.555 26.750 22.855 39.340 ;
      LAYER mcon ;
        RECT 9.740 50.040 9.980 50.280 ;
        RECT 16.930 48.620 17.230 48.920 ;
        RECT 17.420 48.620 17.720 48.920 ;
        RECT 17.910 48.620 18.210 48.920 ;
        RECT 19.800 48.620 20.100 48.920 ;
        RECT 20.290 48.620 20.590 48.920 ;
        RECT 20.780 48.620 21.080 48.920 ;
        RECT 12.460 32.920 12.760 33.220 ;
        RECT 12.950 32.920 13.250 33.220 ;
        RECT 13.440 32.920 13.740 33.220 ;
        RECT 8.180 31.560 8.480 31.860 ;
        RECT 22.555 31.560 22.855 31.860 ;
      LAYER met1 ;
        RECT 9.680 50.010 17.840 50.310 ;
        RECT 13.260 49.950 17.840 50.010 ;
        RECT 13.260 43.360 13.620 49.950 ;
        RECT 17.480 48.950 17.840 49.950 ;
        RECT 16.870 48.590 21.140 48.950 ;
        RECT 4.990 43.000 13.620 43.360 ;
        RECT 4.990 31.890 5.350 43.000 ;
        RECT 12.300 32.890 13.800 33.250 ;
        RECT 12.890 31.890 13.250 32.890 ;
        RECT 4.990 31.530 22.915 31.890 ;
      LAYER via ;
        RECT 7.140 31.530 7.500 31.890 ;
      LAYER met2 ;
        RECT 7.110 24.280 7.530 31.890 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 18.855 42.500 19.155 55.090 ;
        RECT 28.920 48.950 29.300 49.000 ;
        RECT 27.970 48.590 29.300 48.950 ;
        RECT 28.920 48.540 29.300 48.590 ;
        RECT 33.230 42.500 33.530 55.090 ;
        RECT 35.590 48.950 35.970 49.000 ;
        RECT 34.640 48.590 35.970 48.950 ;
        RECT 35.590 48.540 35.970 48.590 ;
        RECT 37.460 48.950 37.840 49.000 ;
        RECT 37.460 48.590 38.790 48.950 ;
        RECT 37.460 48.540 37.840 48.590 ;
      LAYER mcon ;
        RECT 18.855 49.980 19.155 50.280 ;
        RECT 33.230 49.980 33.530 50.280 ;
        RECT 27.970 48.620 28.270 48.920 ;
        RECT 28.460 48.620 28.760 48.920 ;
        RECT 28.950 48.620 29.250 48.920 ;
        RECT 34.640 48.620 34.940 48.920 ;
        RECT 35.130 48.620 35.430 48.920 ;
        RECT 35.620 48.620 35.920 48.920 ;
        RECT 37.510 48.620 37.810 48.920 ;
        RECT 38.000 48.620 38.300 48.920 ;
        RECT 38.490 48.620 38.790 48.920 ;
      LAYER met1 ;
        RECT 18.795 49.950 35.550 50.310 ;
        RECT 28.460 48.950 28.820 49.950 ;
        RECT 35.190 48.950 35.550 49.950 ;
        RECT 27.910 48.590 29.410 48.950 ;
        RECT 34.580 48.590 38.850 48.950 ;
      LAYER via ;
        RECT 27.110 49.950 27.470 50.310 ;
      LAYER met2 ;
        RECT 27.080 49.950 27.500 57.500 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 36.565 42.500 36.865 55.090 ;
        RECT 46.630 48.950 47.010 49.000 ;
        RECT 45.680 48.590 47.010 48.950 ;
        RECT 46.630 48.540 47.010 48.590 ;
        RECT 50.940 42.500 51.240 55.090 ;
        RECT 53.300 48.950 53.680 49.000 ;
        RECT 52.350 48.590 53.680 48.950 ;
        RECT 53.300 48.540 53.680 48.590 ;
        RECT 55.170 48.950 55.550 49.000 ;
        RECT 55.170 48.590 56.500 48.950 ;
        RECT 55.170 48.540 55.550 48.590 ;
      LAYER mcon ;
        RECT 36.565 49.980 36.865 50.280 ;
        RECT 50.940 49.980 51.240 50.280 ;
        RECT 45.680 48.620 45.980 48.920 ;
        RECT 46.170 48.620 46.470 48.920 ;
        RECT 46.660 48.620 46.960 48.920 ;
        RECT 52.350 48.620 52.650 48.920 ;
        RECT 52.840 48.620 53.140 48.920 ;
        RECT 53.330 48.620 53.630 48.920 ;
        RECT 55.220 48.620 55.520 48.920 ;
        RECT 55.710 48.620 56.010 48.920 ;
        RECT 56.200 48.620 56.500 48.920 ;
      LAYER met1 ;
        RECT 36.505 49.950 53.260 50.310 ;
        RECT 46.170 48.950 46.530 49.950 ;
        RECT 52.900 48.950 53.260 49.950 ;
        RECT 45.620 48.590 47.120 48.950 ;
        RECT 52.290 48.590 56.560 48.950 ;
      LAYER via ;
        RECT 51.480 49.950 51.840 50.310 ;
      LAYER met2 ;
        RECT 51.450 49.950 51.870 57.500 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 54.275 42.500 54.575 55.090 ;
        RECT 64.340 48.950 64.720 49.000 ;
        RECT 63.390 48.590 64.720 48.950 ;
        RECT 64.340 48.540 64.720 48.590 ;
        RECT 68.650 42.500 68.950 55.090 ;
        RECT 71.010 48.950 71.390 49.000 ;
        RECT 70.060 48.590 71.390 48.950 ;
        RECT 71.010 48.540 71.390 48.590 ;
        RECT 72.880 48.950 73.260 49.000 ;
        RECT 72.880 48.590 74.210 48.950 ;
        RECT 72.880 48.540 73.260 48.590 ;
      LAYER mcon ;
        RECT 54.275 49.980 54.575 50.280 ;
        RECT 68.650 49.980 68.950 50.280 ;
        RECT 63.390 48.620 63.690 48.920 ;
        RECT 63.880 48.620 64.180 48.920 ;
        RECT 64.370 48.620 64.670 48.920 ;
        RECT 70.060 48.620 70.360 48.920 ;
        RECT 70.550 48.620 70.850 48.920 ;
        RECT 71.040 48.620 71.340 48.920 ;
        RECT 72.930 48.620 73.230 48.920 ;
        RECT 73.420 48.620 73.720 48.920 ;
        RECT 73.910 48.620 74.210 48.920 ;
      LAYER met1 ;
        RECT 54.215 49.950 70.970 50.310 ;
        RECT 63.880 48.950 64.240 49.950 ;
        RECT 70.610 48.950 70.970 49.950 ;
        RECT 63.330 48.590 64.830 48.950 ;
        RECT 70.000 48.590 74.270 48.950 ;
      LAYER via ;
        RECT 68.270 49.950 68.630 50.310 ;
      LAYER met2 ;
        RECT 68.240 49.950 68.660 57.500 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 71.985 42.500 72.285 55.090 ;
        RECT 82.050 48.950 82.430 49.000 ;
        RECT 81.100 48.590 82.430 48.950 ;
        RECT 82.050 48.540 82.430 48.590 ;
        RECT 86.360 42.500 86.660 55.090 ;
        RECT 88.720 48.950 89.100 49.000 ;
        RECT 87.770 48.590 89.100 48.950 ;
        RECT 88.720 48.540 89.100 48.590 ;
        RECT 90.590 48.950 90.970 49.000 ;
        RECT 90.590 48.590 91.920 48.950 ;
        RECT 90.590 48.540 90.970 48.590 ;
      LAYER mcon ;
        RECT 71.985 49.980 72.285 50.280 ;
        RECT 86.360 49.980 86.660 50.280 ;
        RECT 81.100 48.620 81.400 48.920 ;
        RECT 81.590 48.620 81.890 48.920 ;
        RECT 82.080 48.620 82.380 48.920 ;
        RECT 87.770 48.620 88.070 48.920 ;
        RECT 88.260 48.620 88.560 48.920 ;
        RECT 88.750 48.620 89.050 48.920 ;
        RECT 90.640 48.620 90.940 48.920 ;
        RECT 91.130 48.620 91.430 48.920 ;
        RECT 91.620 48.620 91.920 48.920 ;
      LAYER met1 ;
        RECT 71.925 49.950 88.680 50.310 ;
        RECT 81.590 48.950 81.950 49.950 ;
        RECT 88.320 48.950 88.680 49.950 ;
        RECT 81.040 48.590 82.540 48.950 ;
        RECT 87.710 48.590 91.980 48.950 ;
      LAYER via ;
        RECT 83.570 49.950 83.930 50.310 ;
      LAYER met2 ;
        RECT 83.540 49.950 83.960 57.500 ;
    END
  END p[9]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 57.000000 ;
    ANTENNADIFFAREA 5.800000 ;
    PORT
      LAYER li1 ;
        RECT 89.695 42.500 89.995 55.090 ;
        RECT 99.760 48.950 100.140 49.000 ;
        RECT 98.810 48.590 100.140 48.950 ;
        RECT 99.760 48.540 100.140 48.590 ;
        RECT 104.070 42.500 104.370 55.090 ;
        RECT 110.130 33.250 110.510 33.300 ;
        RECT 109.180 32.890 110.510 33.250 ;
        RECT 110.130 32.840 110.510 32.890 ;
        RECT 112.000 33.250 112.380 33.300 ;
        RECT 112.000 32.890 113.330 33.250 ;
        RECT 112.000 32.840 112.380 32.890 ;
      LAYER mcon ;
        RECT 89.695 49.980 89.995 50.280 ;
        RECT 104.070 49.980 104.370 50.280 ;
        RECT 98.810 48.620 99.110 48.920 ;
        RECT 99.300 48.620 99.600 48.920 ;
        RECT 99.790 48.620 100.090 48.920 ;
        RECT 109.180 32.920 109.480 33.220 ;
        RECT 109.670 32.920 109.970 33.220 ;
        RECT 110.160 32.920 110.460 33.220 ;
        RECT 112.050 32.920 112.350 33.220 ;
        RECT 112.540 32.920 112.840 33.220 ;
        RECT 113.030 32.920 113.330 33.220 ;
      LAYER met1 ;
        RECT 89.635 49.950 107.720 50.310 ;
        RECT 99.300 48.950 99.660 49.950 ;
        RECT 98.750 48.590 100.250 48.950 ;
        RECT 107.360 43.360 107.720 49.950 ;
        RECT 107.360 43.000 116.860 43.360 ;
        RECT 109.120 32.890 113.390 33.250 ;
        RECT 112.420 31.890 112.780 32.890 ;
        RECT 116.500 31.890 116.860 43.000 ;
        RECT 112.420 31.530 116.860 31.890 ;
      LAYER via ;
        RECT 106.000 49.950 106.360 50.310 ;
      LAYER met2 ;
        RECT 105.970 49.950 106.390 57.500 ;
    END
  END p[10]
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER li1 ;
        RECT 6.775 50.300 7.235 50.525 ;
        RECT -0.400 50.000 7.235 50.300 ;
        RECT 6.775 49.795 7.235 50.000 ;
      LAYER mcon ;
        RECT -0.380 50.020 -0.120 50.280 ;
      LAYER met1 ;
        RECT -0.450 49.950 -0.050 50.350 ;
    END
  END enb
  PIN input_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 115.015 44.500 116.000 45.500 ;
        RECT 115.015 43.500 115.380 44.500 ;
      LAYER mcon ;
        RECT 115.105 45.100 115.405 45.400 ;
        RECT 115.595 45.100 115.895 45.400 ;
        RECT 115.105 44.600 115.405 44.900 ;
        RECT 115.595 44.600 115.895 44.900 ;
      LAYER met1 ;
        RECT 115.015 44.500 116.000 45.500 ;
      LAYER via ;
        RECT 115.085 45.080 115.425 45.420 ;
        RECT 115.575 45.080 115.915 45.420 ;
        RECT 115.085 44.580 115.425 44.920 ;
        RECT 115.575 44.580 115.915 44.920 ;
      LAYER met2 ;
        RECT 115.015 45.000 123.100 45.500 ;
        RECT 115.015 44.500 116.000 45.000 ;
    END
  END input_analog
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 6.500 50.105 9.180 51.950 ;
        RECT 10.495 50.105 12.255 51.950 ;
        RECT 15.980 48.965 105.050 55.840 ;
        RECT 27.020 48.960 34.210 48.965 ;
        RECT 44.730 48.960 51.920 48.965 ;
        RECT 62.440 48.960 69.630 48.965 ;
        RECT 80.150 48.960 87.340 48.965 ;
        RECT 97.860 48.960 105.050 48.965 ;
        RECT 7.500 32.875 14.690 32.880 ;
        RECT 25.210 32.875 32.400 32.880 ;
        RECT 42.920 32.875 50.110 32.880 ;
        RECT 60.630 32.875 67.820 32.880 ;
        RECT 78.340 32.875 85.530 32.880 ;
        RECT 96.050 32.875 103.240 32.880 ;
        RECT 7.500 26.000 114.280 32.875 ;
      LAYER li1 ;
        RECT 16.160 55.660 18.050 55.690 ;
        RECT 19.840 55.660 23.690 55.690 ;
        RECT 25.350 55.660 29.200 55.690 ;
        RECT 31.040 55.660 32.440 55.690 ;
        RECT 33.870 55.660 35.760 55.690 ;
        RECT 37.550 55.660 41.400 55.690 ;
        RECT 43.060 55.660 46.910 55.690 ;
        RECT 48.750 55.660 50.150 55.690 ;
        RECT 51.580 55.660 53.470 55.690 ;
        RECT 55.260 55.660 59.110 55.690 ;
        RECT 60.770 55.660 64.620 55.690 ;
        RECT 66.460 55.660 67.860 55.690 ;
        RECT 69.290 55.660 71.180 55.690 ;
        RECT 72.970 55.660 76.820 55.690 ;
        RECT 78.480 55.660 82.330 55.690 ;
        RECT 84.170 55.660 85.570 55.690 ;
        RECT 87.000 55.660 88.890 55.690 ;
        RECT 90.680 55.660 94.530 55.690 ;
        RECT 96.190 55.660 100.040 55.690 ;
        RECT 101.880 55.660 103.280 55.690 ;
        RECT 16.160 55.490 104.870 55.660 ;
        RECT 16.160 55.330 18.050 55.490 ;
        RECT 19.840 55.330 23.690 55.490 ;
        RECT 25.350 55.330 29.200 55.490 ;
        RECT 31.040 55.330 32.440 55.490 ;
        RECT 33.870 55.330 35.760 55.490 ;
        RECT 37.550 55.330 41.400 55.490 ;
        RECT 43.060 55.330 46.910 55.490 ;
        RECT 48.750 55.330 50.150 55.490 ;
        RECT 51.580 55.330 53.470 55.490 ;
        RECT 55.260 55.330 59.110 55.490 ;
        RECT 60.770 55.330 64.620 55.490 ;
        RECT 66.460 55.330 67.860 55.490 ;
        RECT 69.290 55.330 71.180 55.490 ;
        RECT 72.970 55.330 76.820 55.490 ;
        RECT 78.480 55.330 82.330 55.490 ;
        RECT 84.170 55.330 85.570 55.490 ;
        RECT 87.000 55.330 88.890 55.490 ;
        RECT 90.680 55.330 94.530 55.490 ;
        RECT 96.190 55.330 100.040 55.490 ;
        RECT 101.880 55.330 103.280 55.490 ;
        RECT 6.690 51.605 7.690 51.770 ;
        RECT 10.685 51.605 11.685 51.770 ;
        RECT 6.690 51.435 8.990 51.605 ;
        RECT 10.685 51.435 12.065 51.605 ;
        RECT 7.205 51.035 8.140 51.435 ;
        RECT 10.960 50.710 11.290 51.435 ;
        RECT 16.160 50.460 16.330 55.330 ;
        RECT 16.670 50.040 16.960 55.330 ;
        RECT 21.050 50.040 21.340 55.330 ;
        RECT 21.680 50.460 21.850 55.330 ;
        RECT 22.190 50.040 22.480 55.330 ;
        RECT 26.570 50.040 26.860 55.330 ;
        RECT 27.200 50.460 27.370 55.330 ;
        RECT 27.710 50.030 28.000 55.330 ;
        RECT 31.040 50.030 31.330 55.330 ;
        RECT 33.870 50.460 34.040 55.330 ;
        RECT 34.380 50.040 34.670 55.330 ;
        RECT 38.760 50.040 39.050 55.330 ;
        RECT 39.390 50.460 39.560 55.330 ;
        RECT 39.900 50.040 40.190 55.330 ;
        RECT 44.280 50.040 44.570 55.330 ;
        RECT 44.910 50.460 45.080 55.330 ;
        RECT 45.420 50.030 45.710 55.330 ;
        RECT 48.750 50.030 49.040 55.330 ;
        RECT 51.580 50.460 51.750 55.330 ;
        RECT 52.090 50.040 52.380 55.330 ;
        RECT 56.470 50.040 56.760 55.330 ;
        RECT 57.100 50.460 57.270 55.330 ;
        RECT 57.610 50.040 57.900 55.330 ;
        RECT 61.990 50.040 62.280 55.330 ;
        RECT 62.620 50.460 62.790 55.330 ;
        RECT 63.130 50.030 63.420 55.330 ;
        RECT 66.460 50.030 66.750 55.330 ;
        RECT 69.290 50.460 69.460 55.330 ;
        RECT 69.800 50.040 70.090 55.330 ;
        RECT 74.180 50.040 74.470 55.330 ;
        RECT 74.810 50.460 74.980 55.330 ;
        RECT 75.320 50.040 75.610 55.330 ;
        RECT 79.700 50.040 79.990 55.330 ;
        RECT 80.330 50.460 80.500 55.330 ;
        RECT 80.840 50.030 81.130 55.330 ;
        RECT 84.170 50.030 84.460 55.330 ;
        RECT 87.000 50.460 87.170 55.330 ;
        RECT 87.510 50.040 87.800 55.330 ;
        RECT 91.890 50.040 92.180 55.330 ;
        RECT 92.520 50.460 92.690 55.330 ;
        RECT 93.030 50.040 93.320 55.330 ;
        RECT 97.410 50.040 97.700 55.330 ;
        RECT 98.040 50.460 98.210 55.330 ;
        RECT 98.550 50.030 98.840 55.330 ;
        RECT 101.880 50.030 102.170 55.330 ;
        RECT 10.380 26.510 10.670 31.810 ;
        RECT 13.710 26.510 14.000 31.810 ;
        RECT 14.340 26.510 14.510 31.380 ;
        RECT 14.850 26.510 15.140 31.800 ;
        RECT 19.230 26.510 19.520 31.800 ;
        RECT 19.860 26.510 20.030 31.380 ;
        RECT 20.370 26.510 20.660 31.800 ;
        RECT 24.750 26.510 25.040 31.800 ;
        RECT 25.380 26.510 25.550 31.380 ;
        RECT 28.090 26.510 28.380 31.810 ;
        RECT 31.420 26.510 31.710 31.810 ;
        RECT 32.050 26.510 32.220 31.380 ;
        RECT 32.560 26.510 32.850 31.800 ;
        RECT 36.940 26.510 37.230 31.800 ;
        RECT 37.570 26.510 37.740 31.380 ;
        RECT 38.080 26.510 38.370 31.800 ;
        RECT 42.460 26.510 42.750 31.800 ;
        RECT 43.090 26.510 43.260 31.380 ;
        RECT 45.800 26.510 46.090 31.810 ;
        RECT 49.130 26.510 49.420 31.810 ;
        RECT 49.760 26.510 49.930 31.380 ;
        RECT 50.270 26.510 50.560 31.800 ;
        RECT 54.650 26.510 54.940 31.800 ;
        RECT 55.280 26.510 55.450 31.380 ;
        RECT 55.790 26.510 56.080 31.800 ;
        RECT 60.170 26.510 60.460 31.800 ;
        RECT 60.800 26.510 60.970 31.380 ;
        RECT 63.510 26.510 63.800 31.810 ;
        RECT 66.840 26.510 67.130 31.810 ;
        RECT 67.470 26.510 67.640 31.380 ;
        RECT 67.980 26.510 68.270 31.800 ;
        RECT 72.360 26.510 72.650 31.800 ;
        RECT 72.990 26.510 73.160 31.380 ;
        RECT 73.500 26.510 73.790 31.800 ;
        RECT 77.880 26.510 78.170 31.800 ;
        RECT 78.510 26.510 78.680 31.380 ;
        RECT 81.220 26.510 81.510 31.810 ;
        RECT 84.550 26.510 84.840 31.810 ;
        RECT 85.180 26.510 85.350 31.380 ;
        RECT 85.690 26.510 85.980 31.800 ;
        RECT 90.070 26.510 90.360 31.800 ;
        RECT 90.700 26.510 90.870 31.380 ;
        RECT 91.210 26.510 91.500 31.800 ;
        RECT 95.590 26.510 95.880 31.800 ;
        RECT 96.220 26.510 96.390 31.380 ;
        RECT 98.930 26.510 99.220 31.810 ;
        RECT 102.260 26.510 102.550 31.810 ;
        RECT 102.890 26.510 103.060 31.380 ;
        RECT 103.400 26.510 103.690 31.800 ;
        RECT 107.780 26.510 108.070 31.800 ;
        RECT 108.410 26.510 108.580 31.380 ;
        RECT 108.920 26.510 109.210 31.800 ;
        RECT 113.300 26.510 113.590 31.800 ;
        RECT 113.930 26.510 114.100 31.380 ;
        RECT 9.270 26.350 10.670 26.510 ;
        RECT 12.510 26.350 16.360 26.510 ;
        RECT 18.020 26.350 21.870 26.510 ;
        RECT 23.660 26.350 25.550 26.510 ;
        RECT 26.980 26.350 28.380 26.510 ;
        RECT 30.220 26.350 34.070 26.510 ;
        RECT 35.730 26.350 39.580 26.510 ;
        RECT 41.370 26.350 43.260 26.510 ;
        RECT 44.690 26.350 46.090 26.510 ;
        RECT 47.930 26.350 51.780 26.510 ;
        RECT 53.440 26.350 57.290 26.510 ;
        RECT 59.080 26.350 60.970 26.510 ;
        RECT 62.400 26.350 63.800 26.510 ;
        RECT 65.640 26.350 69.490 26.510 ;
        RECT 71.150 26.350 75.000 26.510 ;
        RECT 76.790 26.350 78.680 26.510 ;
        RECT 80.110 26.350 81.510 26.510 ;
        RECT 83.350 26.350 87.200 26.510 ;
        RECT 88.860 26.350 92.710 26.510 ;
        RECT 94.500 26.350 96.390 26.510 ;
        RECT 97.820 26.350 99.220 26.510 ;
        RECT 101.060 26.350 104.910 26.510 ;
        RECT 106.570 26.350 110.420 26.510 ;
        RECT 112.210 26.350 114.100 26.510 ;
        RECT 7.680 26.180 114.100 26.350 ;
        RECT 9.270 26.150 10.670 26.180 ;
        RECT 12.510 26.150 16.360 26.180 ;
        RECT 18.020 26.150 21.870 26.180 ;
        RECT 23.660 26.150 25.550 26.180 ;
        RECT 26.980 26.150 28.380 26.180 ;
        RECT 30.220 26.150 34.070 26.180 ;
        RECT 35.730 26.150 39.580 26.180 ;
        RECT 41.370 26.150 43.260 26.180 ;
        RECT 44.690 26.150 46.090 26.180 ;
        RECT 47.930 26.150 51.780 26.180 ;
        RECT 53.440 26.150 57.290 26.180 ;
        RECT 59.080 26.150 60.970 26.180 ;
        RECT 62.400 26.150 63.800 26.180 ;
        RECT 65.640 26.150 69.490 26.180 ;
        RECT 71.150 26.150 75.000 26.180 ;
        RECT 76.790 26.150 78.680 26.180 ;
        RECT 80.110 26.150 81.510 26.180 ;
        RECT 83.350 26.150 87.200 26.180 ;
        RECT 88.860 26.150 92.710 26.180 ;
        RECT 94.500 26.150 96.390 26.180 ;
        RECT 97.820 26.150 99.220 26.180 ;
        RECT 101.060 26.150 104.910 26.180 ;
        RECT 106.570 26.150 110.420 26.180 ;
        RECT 112.210 26.150 114.100 26.180 ;
      LAYER mcon ;
        RECT 16.220 55.360 16.520 55.660 ;
        RECT 16.710 55.360 17.010 55.660 ;
        RECT 17.200 55.360 17.500 55.660 ;
        RECT 17.690 55.360 17.990 55.660 ;
        RECT 19.900 55.360 20.200 55.660 ;
        RECT 20.390 55.360 20.690 55.660 ;
        RECT 20.880 55.360 21.180 55.660 ;
        RECT 21.370 55.360 21.670 55.660 ;
        RECT 21.860 55.360 22.160 55.660 ;
        RECT 22.350 55.360 22.650 55.660 ;
        RECT 22.840 55.360 23.140 55.660 ;
        RECT 23.330 55.360 23.630 55.660 ;
        RECT 25.410 55.360 25.710 55.660 ;
        RECT 25.900 55.360 26.200 55.660 ;
        RECT 26.390 55.360 26.690 55.660 ;
        RECT 26.880 55.360 27.180 55.660 ;
        RECT 27.370 55.360 27.670 55.660 ;
        RECT 27.860 55.360 28.160 55.660 ;
        RECT 28.350 55.360 28.650 55.660 ;
        RECT 28.840 55.360 29.140 55.660 ;
        RECT 31.100 55.360 31.400 55.660 ;
        RECT 31.590 55.360 31.890 55.660 ;
        RECT 32.080 55.360 32.380 55.660 ;
        RECT 33.930 55.360 34.230 55.660 ;
        RECT 34.420 55.360 34.720 55.660 ;
        RECT 34.910 55.360 35.210 55.660 ;
        RECT 35.400 55.360 35.700 55.660 ;
        RECT 37.610 55.360 37.910 55.660 ;
        RECT 38.100 55.360 38.400 55.660 ;
        RECT 38.590 55.360 38.890 55.660 ;
        RECT 39.080 55.360 39.380 55.660 ;
        RECT 39.570 55.360 39.870 55.660 ;
        RECT 40.060 55.360 40.360 55.660 ;
        RECT 40.550 55.360 40.850 55.660 ;
        RECT 41.040 55.360 41.340 55.660 ;
        RECT 43.120 55.360 43.420 55.660 ;
        RECT 43.610 55.360 43.910 55.660 ;
        RECT 44.100 55.360 44.400 55.660 ;
        RECT 44.590 55.360 44.890 55.660 ;
        RECT 45.080 55.360 45.380 55.660 ;
        RECT 45.570 55.360 45.870 55.660 ;
        RECT 46.060 55.360 46.360 55.660 ;
        RECT 46.550 55.360 46.850 55.660 ;
        RECT 48.810 55.360 49.110 55.660 ;
        RECT 49.300 55.360 49.600 55.660 ;
        RECT 49.790 55.360 50.090 55.660 ;
        RECT 51.640 55.360 51.940 55.660 ;
        RECT 52.130 55.360 52.430 55.660 ;
        RECT 52.620 55.360 52.920 55.660 ;
        RECT 53.110 55.360 53.410 55.660 ;
        RECT 55.320 55.360 55.620 55.660 ;
        RECT 55.810 55.360 56.110 55.660 ;
        RECT 56.300 55.360 56.600 55.660 ;
        RECT 56.790 55.360 57.090 55.660 ;
        RECT 57.280 55.360 57.580 55.660 ;
        RECT 57.770 55.360 58.070 55.660 ;
        RECT 58.260 55.360 58.560 55.660 ;
        RECT 58.750 55.360 59.050 55.660 ;
        RECT 60.830 55.360 61.130 55.660 ;
        RECT 61.320 55.360 61.620 55.660 ;
        RECT 61.810 55.360 62.110 55.660 ;
        RECT 62.300 55.360 62.600 55.660 ;
        RECT 62.790 55.360 63.090 55.660 ;
        RECT 63.280 55.360 63.580 55.660 ;
        RECT 63.770 55.360 64.070 55.660 ;
        RECT 64.260 55.360 64.560 55.660 ;
        RECT 66.520 55.360 66.820 55.660 ;
        RECT 67.010 55.360 67.310 55.660 ;
        RECT 67.500 55.360 67.800 55.660 ;
        RECT 69.350 55.360 69.650 55.660 ;
        RECT 69.840 55.360 70.140 55.660 ;
        RECT 70.330 55.360 70.630 55.660 ;
        RECT 70.820 55.360 71.120 55.660 ;
        RECT 73.030 55.360 73.330 55.660 ;
        RECT 73.520 55.360 73.820 55.660 ;
        RECT 74.010 55.360 74.310 55.660 ;
        RECT 74.500 55.360 74.800 55.660 ;
        RECT 74.990 55.360 75.290 55.660 ;
        RECT 75.480 55.360 75.780 55.660 ;
        RECT 75.970 55.360 76.270 55.660 ;
        RECT 76.460 55.360 76.760 55.660 ;
        RECT 78.540 55.360 78.840 55.660 ;
        RECT 79.030 55.360 79.330 55.660 ;
        RECT 79.520 55.360 79.820 55.660 ;
        RECT 80.010 55.360 80.310 55.660 ;
        RECT 80.500 55.360 80.800 55.660 ;
        RECT 80.990 55.360 81.290 55.660 ;
        RECT 81.480 55.360 81.780 55.660 ;
        RECT 81.970 55.360 82.270 55.660 ;
        RECT 84.230 55.360 84.530 55.660 ;
        RECT 84.720 55.360 85.020 55.660 ;
        RECT 85.210 55.360 85.510 55.660 ;
        RECT 87.060 55.360 87.360 55.660 ;
        RECT 87.550 55.360 87.850 55.660 ;
        RECT 88.040 55.360 88.340 55.660 ;
        RECT 88.530 55.360 88.830 55.660 ;
        RECT 90.740 55.360 91.040 55.660 ;
        RECT 91.230 55.360 91.530 55.660 ;
        RECT 91.720 55.360 92.020 55.660 ;
        RECT 92.210 55.360 92.510 55.660 ;
        RECT 92.700 55.360 93.000 55.660 ;
        RECT 93.190 55.360 93.490 55.660 ;
        RECT 93.680 55.360 93.980 55.660 ;
        RECT 94.170 55.360 94.470 55.660 ;
        RECT 96.250 55.360 96.550 55.660 ;
        RECT 96.740 55.360 97.040 55.660 ;
        RECT 97.230 55.360 97.530 55.660 ;
        RECT 97.720 55.360 98.020 55.660 ;
        RECT 98.210 55.360 98.510 55.660 ;
        RECT 98.700 55.360 99.000 55.660 ;
        RECT 99.190 55.360 99.490 55.660 ;
        RECT 99.680 55.360 99.980 55.660 ;
        RECT 101.940 55.360 102.240 55.660 ;
        RECT 102.430 55.360 102.730 55.660 ;
        RECT 102.920 55.360 103.220 55.660 ;
        RECT 6.835 51.435 7.005 51.605 ;
        RECT 7.295 51.435 7.465 51.605 ;
        RECT 7.755 51.435 7.925 51.605 ;
        RECT 8.215 51.435 8.385 51.605 ;
        RECT 8.675 51.435 8.845 51.605 ;
        RECT 10.830 51.435 11.000 51.605 ;
        RECT 11.290 51.435 11.460 51.605 ;
        RECT 11.750 51.435 11.920 51.605 ;
        RECT 9.330 26.180 9.630 26.480 ;
        RECT 9.820 26.180 10.120 26.480 ;
        RECT 10.310 26.180 10.610 26.480 ;
        RECT 12.570 26.180 12.870 26.480 ;
        RECT 13.060 26.180 13.360 26.480 ;
        RECT 13.550 26.180 13.850 26.480 ;
        RECT 14.040 26.180 14.340 26.480 ;
        RECT 14.530 26.180 14.830 26.480 ;
        RECT 15.020 26.180 15.320 26.480 ;
        RECT 15.510 26.180 15.810 26.480 ;
        RECT 16.000 26.180 16.300 26.480 ;
        RECT 18.080 26.180 18.380 26.480 ;
        RECT 18.570 26.180 18.870 26.480 ;
        RECT 19.060 26.180 19.360 26.480 ;
        RECT 19.550 26.180 19.850 26.480 ;
        RECT 20.040 26.180 20.340 26.480 ;
        RECT 20.530 26.180 20.830 26.480 ;
        RECT 21.020 26.180 21.320 26.480 ;
        RECT 21.510 26.180 21.810 26.480 ;
        RECT 23.720 26.180 24.020 26.480 ;
        RECT 24.210 26.180 24.510 26.480 ;
        RECT 24.700 26.180 25.000 26.480 ;
        RECT 25.190 26.180 25.490 26.480 ;
        RECT 27.040 26.180 27.340 26.480 ;
        RECT 27.530 26.180 27.830 26.480 ;
        RECT 28.020 26.180 28.320 26.480 ;
        RECT 30.280 26.180 30.580 26.480 ;
        RECT 30.770 26.180 31.070 26.480 ;
        RECT 31.260 26.180 31.560 26.480 ;
        RECT 31.750 26.180 32.050 26.480 ;
        RECT 32.240 26.180 32.540 26.480 ;
        RECT 32.730 26.180 33.030 26.480 ;
        RECT 33.220 26.180 33.520 26.480 ;
        RECT 33.710 26.180 34.010 26.480 ;
        RECT 35.790 26.180 36.090 26.480 ;
        RECT 36.280 26.180 36.580 26.480 ;
        RECT 36.770 26.180 37.070 26.480 ;
        RECT 37.260 26.180 37.560 26.480 ;
        RECT 37.750 26.180 38.050 26.480 ;
        RECT 38.240 26.180 38.540 26.480 ;
        RECT 38.730 26.180 39.030 26.480 ;
        RECT 39.220 26.180 39.520 26.480 ;
        RECT 41.430 26.180 41.730 26.480 ;
        RECT 41.920 26.180 42.220 26.480 ;
        RECT 42.410 26.180 42.710 26.480 ;
        RECT 42.900 26.180 43.200 26.480 ;
        RECT 44.750 26.180 45.050 26.480 ;
        RECT 45.240 26.180 45.540 26.480 ;
        RECT 45.730 26.180 46.030 26.480 ;
        RECT 47.990 26.180 48.290 26.480 ;
        RECT 48.480 26.180 48.780 26.480 ;
        RECT 48.970 26.180 49.270 26.480 ;
        RECT 49.460 26.180 49.760 26.480 ;
        RECT 49.950 26.180 50.250 26.480 ;
        RECT 50.440 26.180 50.740 26.480 ;
        RECT 50.930 26.180 51.230 26.480 ;
        RECT 51.420 26.180 51.720 26.480 ;
        RECT 53.500 26.180 53.800 26.480 ;
        RECT 53.990 26.180 54.290 26.480 ;
        RECT 54.480 26.180 54.780 26.480 ;
        RECT 54.970 26.180 55.270 26.480 ;
        RECT 55.460 26.180 55.760 26.480 ;
        RECT 55.950 26.180 56.250 26.480 ;
        RECT 56.440 26.180 56.740 26.480 ;
        RECT 56.930 26.180 57.230 26.480 ;
        RECT 59.140 26.180 59.440 26.480 ;
        RECT 59.630 26.180 59.930 26.480 ;
        RECT 60.120 26.180 60.420 26.480 ;
        RECT 60.610 26.180 60.910 26.480 ;
        RECT 62.460 26.180 62.760 26.480 ;
        RECT 62.950 26.180 63.250 26.480 ;
        RECT 63.440 26.180 63.740 26.480 ;
        RECT 65.700 26.180 66.000 26.480 ;
        RECT 66.190 26.180 66.490 26.480 ;
        RECT 66.680 26.180 66.980 26.480 ;
        RECT 67.170 26.180 67.470 26.480 ;
        RECT 67.660 26.180 67.960 26.480 ;
        RECT 68.150 26.180 68.450 26.480 ;
        RECT 68.640 26.180 68.940 26.480 ;
        RECT 69.130 26.180 69.430 26.480 ;
        RECT 71.210 26.180 71.510 26.480 ;
        RECT 71.700 26.180 72.000 26.480 ;
        RECT 72.190 26.180 72.490 26.480 ;
        RECT 72.680 26.180 72.980 26.480 ;
        RECT 73.170 26.180 73.470 26.480 ;
        RECT 73.660 26.180 73.960 26.480 ;
        RECT 74.150 26.180 74.450 26.480 ;
        RECT 74.640 26.180 74.940 26.480 ;
        RECT 76.850 26.180 77.150 26.480 ;
        RECT 77.340 26.180 77.640 26.480 ;
        RECT 77.830 26.180 78.130 26.480 ;
        RECT 78.320 26.180 78.620 26.480 ;
        RECT 80.170 26.180 80.470 26.480 ;
        RECT 80.660 26.180 80.960 26.480 ;
        RECT 81.150 26.180 81.450 26.480 ;
        RECT 83.410 26.180 83.710 26.480 ;
        RECT 83.900 26.180 84.200 26.480 ;
        RECT 84.390 26.180 84.690 26.480 ;
        RECT 84.880 26.180 85.180 26.480 ;
        RECT 85.370 26.180 85.670 26.480 ;
        RECT 85.860 26.180 86.160 26.480 ;
        RECT 86.350 26.180 86.650 26.480 ;
        RECT 86.840 26.180 87.140 26.480 ;
        RECT 88.920 26.180 89.220 26.480 ;
        RECT 89.410 26.180 89.710 26.480 ;
        RECT 89.900 26.180 90.200 26.480 ;
        RECT 90.390 26.180 90.690 26.480 ;
        RECT 90.880 26.180 91.180 26.480 ;
        RECT 91.370 26.180 91.670 26.480 ;
        RECT 91.860 26.180 92.160 26.480 ;
        RECT 92.350 26.180 92.650 26.480 ;
        RECT 94.560 26.180 94.860 26.480 ;
        RECT 95.050 26.180 95.350 26.480 ;
        RECT 95.540 26.180 95.840 26.480 ;
        RECT 96.030 26.180 96.330 26.480 ;
        RECT 97.880 26.180 98.180 26.480 ;
        RECT 98.370 26.180 98.670 26.480 ;
        RECT 98.860 26.180 99.160 26.480 ;
        RECT 101.120 26.180 101.420 26.480 ;
        RECT 101.610 26.180 101.910 26.480 ;
        RECT 102.100 26.180 102.400 26.480 ;
        RECT 102.590 26.180 102.890 26.480 ;
        RECT 103.080 26.180 103.380 26.480 ;
        RECT 103.570 26.180 103.870 26.480 ;
        RECT 104.060 26.180 104.360 26.480 ;
        RECT 104.550 26.180 104.850 26.480 ;
        RECT 106.630 26.180 106.930 26.480 ;
        RECT 107.120 26.180 107.420 26.480 ;
        RECT 107.610 26.180 107.910 26.480 ;
        RECT 108.100 26.180 108.400 26.480 ;
        RECT 108.590 26.180 108.890 26.480 ;
        RECT 109.080 26.180 109.380 26.480 ;
        RECT 109.570 26.180 109.870 26.480 ;
        RECT 110.060 26.180 110.360 26.480 ;
        RECT 112.270 26.180 112.570 26.480 ;
        RECT 112.760 26.180 113.060 26.480 ;
        RECT 113.250 26.180 113.550 26.480 ;
        RECT 113.740 26.180 114.040 26.480 ;
      LAYER met1 ;
        RECT 15.900 55.270 105.050 55.750 ;
        RECT 0.000 51.280 12.065 51.760 ;
        RECT 7.500 26.090 114.280 26.570 ;
      LAYER via ;
        RECT 18.130 55.360 18.430 55.660 ;
        RECT 18.490 55.360 18.790 55.660 ;
        RECT 18.850 55.360 19.150 55.660 ;
        RECT 19.210 55.360 19.510 55.660 ;
        RECT 19.570 55.360 19.870 55.660 ;
        RECT 46.130 55.360 46.430 55.660 ;
        RECT 46.490 55.360 46.790 55.660 ;
        RECT 46.850 55.360 47.150 55.660 ;
        RECT 47.210 55.360 47.510 55.660 ;
        RECT 47.570 55.360 47.870 55.660 ;
        RECT 74.130 55.360 74.430 55.660 ;
        RECT 74.490 55.360 74.790 55.660 ;
        RECT 74.850 55.360 75.150 55.660 ;
        RECT 75.210 55.360 75.510 55.660 ;
        RECT 75.570 55.360 75.870 55.660 ;
        RECT 102.130 55.360 102.430 55.660 ;
        RECT 102.490 55.360 102.790 55.660 ;
        RECT 102.850 55.360 103.150 55.660 ;
        RECT 103.210 55.360 103.510 55.660 ;
        RECT 103.570 55.360 103.870 55.660 ;
        RECT 0.130 51.370 0.430 51.670 ;
        RECT 0.490 51.370 0.790 51.670 ;
        RECT 0.850 51.370 1.150 51.670 ;
        RECT 1.210 51.370 1.510 51.670 ;
        RECT 1.570 51.370 1.870 51.670 ;
        RECT 18.130 26.180 18.430 26.480 ;
        RECT 18.490 26.180 18.790 26.480 ;
        RECT 18.850 26.180 19.150 26.480 ;
        RECT 19.210 26.180 19.510 26.480 ;
        RECT 19.570 26.180 19.870 26.480 ;
        RECT 46.130 26.180 46.430 26.480 ;
        RECT 46.490 26.180 46.790 26.480 ;
        RECT 46.850 26.180 47.150 26.480 ;
        RECT 47.210 26.180 47.510 26.480 ;
        RECT 47.570 26.180 47.870 26.480 ;
        RECT 74.130 26.180 74.430 26.480 ;
        RECT 74.490 26.180 74.790 26.480 ;
        RECT 74.850 26.180 75.150 26.480 ;
        RECT 75.210 26.180 75.510 26.480 ;
        RECT 75.570 26.180 75.870 26.480 ;
        RECT 102.130 26.180 102.430 26.480 ;
        RECT 102.490 26.180 102.790 26.480 ;
        RECT 102.850 26.180 103.150 26.480 ;
        RECT 103.210 26.180 103.510 26.480 ;
        RECT 103.570 26.180 103.870 26.480 ;
      LAYER met2 ;
        RECT 18.000 55.270 20.000 55.750 ;
        RECT 46.000 55.270 48.000 55.750 ;
        RECT 74.000 55.270 76.000 55.750 ;
        RECT 102.000 55.270 104.000 55.750 ;
        RECT 0.000 51.280 2.000 51.760 ;
        RECT 18.000 26.090 20.000 26.570 ;
        RECT 46.000 26.090 48.000 26.570 ;
        RECT 74.000 26.090 76.000 26.570 ;
        RECT 102.000 26.090 104.000 26.570 ;
      LAYER via2 ;
        RECT 18.180 55.350 18.500 55.670 ;
        RECT 18.620 55.350 18.940 55.670 ;
        RECT 19.060 55.350 19.380 55.670 ;
        RECT 19.500 55.350 19.820 55.670 ;
        RECT 46.180 55.350 46.500 55.670 ;
        RECT 46.620 55.350 46.940 55.670 ;
        RECT 47.060 55.350 47.380 55.670 ;
        RECT 47.500 55.350 47.820 55.670 ;
        RECT 74.180 55.350 74.500 55.670 ;
        RECT 74.620 55.350 74.940 55.670 ;
        RECT 75.060 55.350 75.380 55.670 ;
        RECT 75.500 55.350 75.820 55.670 ;
        RECT 102.180 55.350 102.500 55.670 ;
        RECT 102.620 55.350 102.940 55.670 ;
        RECT 103.060 55.350 103.380 55.670 ;
        RECT 103.500 55.350 103.820 55.670 ;
        RECT 0.180 51.360 0.500 51.680 ;
        RECT 0.620 51.360 0.940 51.680 ;
        RECT 1.060 51.360 1.380 51.680 ;
        RECT 1.500 51.360 1.820 51.680 ;
        RECT 18.180 26.170 18.500 26.490 ;
        RECT 18.620 26.170 18.940 26.490 ;
        RECT 19.060 26.170 19.380 26.490 ;
        RECT 19.500 26.170 19.820 26.490 ;
        RECT 46.180 26.170 46.500 26.490 ;
        RECT 46.620 26.170 46.940 26.490 ;
        RECT 47.060 26.170 47.380 26.490 ;
        RECT 47.500 26.170 47.820 26.490 ;
        RECT 74.180 26.170 74.500 26.490 ;
        RECT 74.620 26.170 74.940 26.490 ;
        RECT 75.060 26.170 75.380 26.490 ;
        RECT 75.500 26.170 75.820 26.490 ;
        RECT 102.180 26.170 102.500 26.490 ;
        RECT 102.620 26.170 102.940 26.490 ;
        RECT 103.060 26.170 103.380 26.490 ;
        RECT 103.500 26.170 103.820 26.490 ;
      LAYER met3 ;
        RECT 0.000 91.000 122.000 93.000 ;
        RECT 18.000 55.270 20.000 55.750 ;
        RECT 46.000 55.270 48.000 55.750 ;
        RECT 74.000 55.270 76.000 55.750 ;
        RECT 102.000 55.270 104.000 55.750 ;
        RECT 0.000 51.280 2.000 51.760 ;
        RECT 18.000 26.090 20.000 26.570 ;
        RECT 46.000 26.090 48.000 26.570 ;
        RECT 74.000 26.090 76.000 26.570 ;
        RECT 102.000 26.090 104.000 26.570 ;
        RECT 0.000 -12.000 122.000 -10.000 ;
      LAYER via3 ;
        RECT 0.200 92.400 0.600 92.800 ;
        RECT 0.800 92.400 1.200 92.800 ;
        RECT 1.400 92.400 1.800 92.800 ;
        RECT 18.200 92.400 18.600 92.800 ;
        RECT 18.800 92.400 19.200 92.800 ;
        RECT 19.400 92.400 19.800 92.800 ;
        RECT 46.200 92.400 46.600 92.800 ;
        RECT 46.800 92.400 47.200 92.800 ;
        RECT 47.400 92.400 47.800 92.800 ;
        RECT 74.200 92.400 74.600 92.800 ;
        RECT 74.800 92.400 75.200 92.800 ;
        RECT 75.400 92.400 75.800 92.800 ;
        RECT 102.200 92.400 102.600 92.800 ;
        RECT 102.800 92.400 103.200 92.800 ;
        RECT 103.400 92.400 103.800 92.800 ;
        RECT 120.200 92.400 120.600 92.800 ;
        RECT 120.800 92.400 121.200 92.800 ;
        RECT 121.400 92.400 121.800 92.800 ;
        RECT 0.200 91.800 0.600 92.200 ;
        RECT 0.800 91.800 1.200 92.200 ;
        RECT 1.400 91.800 1.800 92.200 ;
        RECT 18.200 91.800 18.600 92.200 ;
        RECT 18.800 91.800 19.200 92.200 ;
        RECT 19.400 91.800 19.800 92.200 ;
        RECT 46.200 91.800 46.600 92.200 ;
        RECT 46.800 91.800 47.200 92.200 ;
        RECT 47.400 91.800 47.800 92.200 ;
        RECT 74.200 91.800 74.600 92.200 ;
        RECT 74.800 91.800 75.200 92.200 ;
        RECT 75.400 91.800 75.800 92.200 ;
        RECT 102.200 91.800 102.600 92.200 ;
        RECT 102.800 91.800 103.200 92.200 ;
        RECT 103.400 91.800 103.800 92.200 ;
        RECT 120.200 91.800 120.600 92.200 ;
        RECT 120.800 91.800 121.200 92.200 ;
        RECT 121.400 91.800 121.800 92.200 ;
        RECT 0.200 91.200 0.600 91.600 ;
        RECT 0.800 91.200 1.200 91.600 ;
        RECT 1.400 91.200 1.800 91.600 ;
        RECT 18.200 91.200 18.600 91.600 ;
        RECT 18.800 91.200 19.200 91.600 ;
        RECT 19.400 91.200 19.800 91.600 ;
        RECT 46.200 91.200 46.600 91.600 ;
        RECT 46.800 91.200 47.200 91.600 ;
        RECT 47.400 91.200 47.800 91.600 ;
        RECT 74.200 91.200 74.600 91.600 ;
        RECT 74.800 91.200 75.200 91.600 ;
        RECT 75.400 91.200 75.800 91.600 ;
        RECT 102.200 91.200 102.600 91.600 ;
        RECT 102.800 91.200 103.200 91.600 ;
        RECT 103.400 91.200 103.800 91.600 ;
        RECT 120.200 91.200 120.600 91.600 ;
        RECT 120.800 91.200 121.200 91.600 ;
        RECT 121.400 91.200 121.800 91.600 ;
        RECT 18.160 55.330 18.520 55.695 ;
        RECT 18.600 55.330 18.960 55.695 ;
        RECT 19.040 55.330 19.400 55.695 ;
        RECT 19.480 55.330 19.840 55.695 ;
        RECT 46.160 55.330 46.520 55.695 ;
        RECT 46.600 55.330 46.960 55.695 ;
        RECT 47.040 55.330 47.400 55.695 ;
        RECT 47.480 55.330 47.840 55.695 ;
        RECT 74.160 55.330 74.520 55.695 ;
        RECT 74.600 55.330 74.960 55.695 ;
        RECT 75.040 55.330 75.400 55.695 ;
        RECT 75.480 55.330 75.840 55.695 ;
        RECT 102.160 55.330 102.520 55.695 ;
        RECT 102.600 55.330 102.960 55.695 ;
        RECT 103.040 55.330 103.400 55.695 ;
        RECT 103.480 55.330 103.840 55.695 ;
        RECT 0.160 51.340 0.520 51.705 ;
        RECT 0.600 51.340 0.960 51.705 ;
        RECT 1.040 51.340 1.400 51.705 ;
        RECT 1.480 51.340 1.840 51.705 ;
        RECT 18.160 26.150 18.520 26.515 ;
        RECT 18.600 26.150 18.960 26.515 ;
        RECT 19.040 26.150 19.400 26.515 ;
        RECT 19.480 26.150 19.840 26.515 ;
        RECT 46.160 26.150 46.520 26.515 ;
        RECT 46.600 26.150 46.960 26.515 ;
        RECT 47.040 26.150 47.400 26.515 ;
        RECT 47.480 26.150 47.840 26.515 ;
        RECT 74.160 26.150 74.520 26.515 ;
        RECT 74.600 26.150 74.960 26.515 ;
        RECT 75.040 26.150 75.400 26.515 ;
        RECT 75.480 26.150 75.840 26.515 ;
        RECT 102.160 26.150 102.520 26.515 ;
        RECT 102.600 26.150 102.960 26.515 ;
        RECT 103.040 26.150 103.400 26.515 ;
        RECT 103.480 26.150 103.840 26.515 ;
        RECT 0.200 -10.600 0.600 -10.200 ;
        RECT 0.800 -10.600 1.200 -10.200 ;
        RECT 1.400 -10.600 1.800 -10.200 ;
        RECT 18.200 -10.600 18.600 -10.200 ;
        RECT 18.800 -10.600 19.200 -10.200 ;
        RECT 19.400 -10.600 19.800 -10.200 ;
        RECT 46.200 -10.600 46.600 -10.200 ;
        RECT 46.800 -10.600 47.200 -10.200 ;
        RECT 47.400 -10.600 47.800 -10.200 ;
        RECT 74.200 -10.600 74.600 -10.200 ;
        RECT 74.800 -10.600 75.200 -10.200 ;
        RECT 75.400 -10.600 75.800 -10.200 ;
        RECT 102.200 -10.600 102.600 -10.200 ;
        RECT 102.800 -10.600 103.200 -10.200 ;
        RECT 103.400 -10.600 103.800 -10.200 ;
        RECT 120.200 -10.600 120.600 -10.200 ;
        RECT 120.800 -10.600 121.200 -10.200 ;
        RECT 121.400 -10.600 121.800 -10.200 ;
        RECT 0.200 -11.200 0.600 -10.800 ;
        RECT 0.800 -11.200 1.200 -10.800 ;
        RECT 1.400 -11.200 1.800 -10.800 ;
        RECT 18.200 -11.200 18.600 -10.800 ;
        RECT 18.800 -11.200 19.200 -10.800 ;
        RECT 19.400 -11.200 19.800 -10.800 ;
        RECT 46.200 -11.200 46.600 -10.800 ;
        RECT 46.800 -11.200 47.200 -10.800 ;
        RECT 47.400 -11.200 47.800 -10.800 ;
        RECT 74.200 -11.200 74.600 -10.800 ;
        RECT 74.800 -11.200 75.200 -10.800 ;
        RECT 75.400 -11.200 75.800 -10.800 ;
        RECT 102.200 -11.200 102.600 -10.800 ;
        RECT 102.800 -11.200 103.200 -10.800 ;
        RECT 103.400 -11.200 103.800 -10.800 ;
        RECT 120.200 -11.200 120.600 -10.800 ;
        RECT 120.800 -11.200 121.200 -10.800 ;
        RECT 121.400 -11.200 121.800 -10.800 ;
        RECT 0.200 -11.800 0.600 -11.400 ;
        RECT 0.800 -11.800 1.200 -11.400 ;
        RECT 1.400 -11.800 1.800 -11.400 ;
        RECT 18.200 -11.800 18.600 -11.400 ;
        RECT 18.800 -11.800 19.200 -11.400 ;
        RECT 19.400 -11.800 19.800 -11.400 ;
        RECT 46.200 -11.800 46.600 -11.400 ;
        RECT 46.800 -11.800 47.200 -11.400 ;
        RECT 47.400 -11.800 47.800 -11.400 ;
        RECT 74.200 -11.800 74.600 -11.400 ;
        RECT 74.800 -11.800 75.200 -11.400 ;
        RECT 75.400 -11.800 75.800 -11.400 ;
        RECT 102.200 -11.800 102.600 -11.400 ;
        RECT 102.800 -11.800 103.200 -11.400 ;
        RECT 103.400 -11.800 103.800 -11.400 ;
        RECT 120.200 -11.800 120.600 -11.400 ;
        RECT 120.800 -11.800 121.200 -11.400 ;
        RECT 121.400 -11.800 121.800 -11.400 ;
      LAYER met4 ;
        RECT 0.000 -12.000 2.000 93.000 ;
        RECT 18.000 -12.000 20.000 93.000 ;
        RECT 46.000 -12.000 48.000 93.000 ;
        RECT 74.000 -12.000 76.000 93.000 ;
        RECT 102.000 -12.000 104.000 93.000 ;
        RECT 120.000 -12.000 122.000 93.000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 15.000 56.700 106.000 57.000 ;
        RECT 7.205 48.885 8.140 49.285 ;
        RECT 11.460 48.885 11.800 49.545 ;
        RECT 6.690 48.715 8.990 48.885 ;
        RECT 10.685 48.715 12.065 48.885 ;
        RECT 15.000 41.070 15.300 56.700 ;
        RECT 105.700 41.070 106.000 56.700 ;
        RECT 108.500 50.015 110.500 50.380 ;
        RECT 6.700 40.770 115.825 41.070 ;
        RECT 6.700 25.200 7.000 40.770 ;
        RECT 115.500 40.700 115.825 40.770 ;
        RECT 115.500 25.200 115.800 40.700 ;
        RECT 6.700 24.900 115.800 25.200 ;
      LAYER mcon ;
        RECT 32.110 56.700 32.410 57.000 ;
        RECT 32.600 56.700 32.900 57.000 ;
        RECT 33.100 56.700 33.400 57.000 ;
        RECT 33.590 56.700 33.890 57.000 ;
        RECT 60.110 56.700 60.410 57.000 ;
        RECT 60.600 56.700 60.900 57.000 ;
        RECT 61.100 56.700 61.400 57.000 ;
        RECT 61.590 56.700 61.890 57.000 ;
        RECT 88.110 56.700 88.410 57.000 ;
        RECT 88.600 56.700 88.900 57.000 ;
        RECT 89.100 56.700 89.400 57.000 ;
        RECT 89.590 56.700 89.890 57.000 ;
        RECT 6.835 48.715 7.005 48.885 ;
        RECT 7.295 48.715 7.465 48.885 ;
        RECT 7.755 48.715 7.925 48.885 ;
        RECT 8.215 48.715 8.385 48.885 ;
        RECT 8.675 48.715 8.845 48.885 ;
        RECT 10.830 48.715 11.000 48.885 ;
        RECT 11.290 48.715 11.460 48.885 ;
        RECT 11.750 48.715 11.920 48.885 ;
        RECT 108.600 50.050 108.900 50.350 ;
        RECT 109.100 50.050 109.400 50.350 ;
        RECT 109.600 50.050 109.900 50.350 ;
        RECT 110.100 50.050 110.400 50.350 ;
        RECT 32.110 24.900 32.410 25.200 ;
        RECT 32.600 24.900 32.900 25.200 ;
        RECT 33.100 24.900 33.400 25.200 ;
        RECT 33.590 24.900 33.890 25.200 ;
        RECT 60.110 24.900 60.410 25.200 ;
        RECT 60.600 24.900 60.900 25.200 ;
        RECT 61.100 24.900 61.400 25.200 ;
        RECT 61.590 24.900 61.890 25.200 ;
      LAYER met1 ;
        RECT 32.080 56.610 33.920 57.090 ;
        RECT 60.080 56.610 61.920 57.090 ;
        RECT 88.080 56.610 89.920 57.090 ;
        RECT 116.130 50.380 117.870 50.440 ;
        RECT 108.500 50.020 118.000 50.380 ;
        RECT 108.500 50.015 110.505 50.020 ;
        RECT 116.130 49.960 117.870 50.020 ;
        RECT 4.000 48.560 12.065 49.040 ;
        RECT 32.080 24.810 33.920 25.290 ;
        RECT 60.080 24.810 61.920 25.290 ;
      LAYER via ;
        RECT 32.130 56.700 32.430 57.000 ;
        RECT 32.490 56.700 32.790 57.000 ;
        RECT 32.850 56.700 33.150 57.000 ;
        RECT 33.210 56.700 33.510 57.000 ;
        RECT 33.570 56.700 33.870 57.000 ;
        RECT 60.130 56.700 60.430 57.000 ;
        RECT 60.490 56.700 60.790 57.000 ;
        RECT 60.850 56.700 61.150 57.000 ;
        RECT 61.210 56.700 61.510 57.000 ;
        RECT 61.570 56.700 61.870 57.000 ;
        RECT 88.130 56.700 88.430 57.000 ;
        RECT 88.490 56.700 88.790 57.000 ;
        RECT 88.850 56.700 89.150 57.000 ;
        RECT 89.210 56.700 89.510 57.000 ;
        RECT 89.570 56.700 89.870 57.000 ;
        RECT 116.130 50.050 116.430 50.350 ;
        RECT 116.490 50.050 116.790 50.350 ;
        RECT 116.850 50.050 117.150 50.350 ;
        RECT 117.210 50.050 117.510 50.350 ;
        RECT 117.570 50.050 117.870 50.350 ;
        RECT 4.130 48.650 4.430 48.950 ;
        RECT 4.490 48.650 4.790 48.950 ;
        RECT 4.850 48.650 5.150 48.950 ;
        RECT 5.210 48.650 5.510 48.950 ;
        RECT 5.570 48.650 5.870 48.950 ;
        RECT 32.130 24.900 32.430 25.200 ;
        RECT 32.490 24.900 32.790 25.200 ;
        RECT 32.850 24.900 33.150 25.200 ;
        RECT 33.210 24.900 33.510 25.200 ;
        RECT 33.570 24.900 33.870 25.200 ;
        RECT 60.130 24.900 60.430 25.200 ;
        RECT 60.490 24.900 60.790 25.200 ;
        RECT 60.850 24.900 61.150 25.200 ;
        RECT 61.210 24.900 61.510 25.200 ;
        RECT 61.570 24.900 61.870 25.200 ;
      LAYER met2 ;
        RECT 32.000 56.610 34.000 57.090 ;
        RECT 60.000 56.610 62.000 57.090 ;
        RECT 88.000 56.610 90.000 57.090 ;
        RECT 116.000 49.960 118.000 50.440 ;
        RECT 4.000 48.560 6.000 49.040 ;
        RECT 32.000 24.810 34.000 25.290 ;
        RECT 60.000 24.810 62.000 25.290 ;
      LAYER via2 ;
        RECT 32.180 56.690 32.500 57.010 ;
        RECT 32.620 56.690 32.940 57.010 ;
        RECT 33.060 56.690 33.380 57.010 ;
        RECT 33.500 56.690 33.820 57.010 ;
        RECT 60.180 56.690 60.500 57.010 ;
        RECT 60.620 56.690 60.940 57.010 ;
        RECT 61.060 56.690 61.380 57.010 ;
        RECT 61.500 56.690 61.820 57.010 ;
        RECT 88.180 56.690 88.500 57.010 ;
        RECT 88.620 56.690 88.940 57.010 ;
        RECT 89.060 56.690 89.380 57.010 ;
        RECT 89.500 56.690 89.820 57.010 ;
        RECT 116.180 50.040 116.500 50.360 ;
        RECT 116.620 50.040 116.940 50.360 ;
        RECT 117.060 50.040 117.380 50.360 ;
        RECT 117.500 50.040 117.820 50.360 ;
        RECT 4.180 48.640 4.500 48.960 ;
        RECT 4.620 48.640 4.940 48.960 ;
        RECT 5.060 48.640 5.380 48.960 ;
        RECT 5.500 48.640 5.820 48.960 ;
        RECT 32.180 24.890 32.500 25.210 ;
        RECT 32.620 24.890 32.940 25.210 ;
        RECT 33.060 24.890 33.380 25.210 ;
        RECT 33.500 24.890 33.820 25.210 ;
        RECT 60.180 24.890 60.500 25.210 ;
        RECT 60.620 24.890 60.940 25.210 ;
        RECT 61.060 24.890 61.380 25.210 ;
        RECT 61.500 24.890 61.820 25.210 ;
      LAYER met3 ;
        RECT 4.000 87.000 118.000 89.000 ;
        RECT 32.000 56.610 34.000 57.090 ;
        RECT 60.000 56.610 62.000 57.090 ;
        RECT 88.000 56.610 90.000 57.090 ;
        RECT 116.000 49.960 118.000 50.440 ;
        RECT 4.000 48.560 6.000 49.040 ;
        RECT 32.000 24.810 34.000 25.290 ;
        RECT 60.000 24.810 62.000 25.290 ;
        RECT 4.000 -8.000 118.000 -6.000 ;
      LAYER via3 ;
        RECT 4.200 88.400 4.600 88.800 ;
        RECT 4.800 88.400 5.200 88.800 ;
        RECT 5.400 88.400 5.800 88.800 ;
        RECT 32.200 88.400 32.600 88.800 ;
        RECT 32.800 88.400 33.200 88.800 ;
        RECT 33.400 88.400 33.800 88.800 ;
        RECT 60.200 88.400 60.600 88.800 ;
        RECT 60.800 88.400 61.200 88.800 ;
        RECT 61.400 88.400 61.800 88.800 ;
        RECT 88.200 88.400 88.600 88.800 ;
        RECT 88.800 88.400 89.200 88.800 ;
        RECT 89.400 88.400 89.800 88.800 ;
        RECT 116.200 88.400 116.600 88.800 ;
        RECT 116.800 88.400 117.200 88.800 ;
        RECT 117.400 88.400 117.800 88.800 ;
        RECT 4.200 87.800 4.600 88.200 ;
        RECT 4.800 87.800 5.200 88.200 ;
        RECT 5.400 87.800 5.800 88.200 ;
        RECT 32.200 87.800 32.600 88.200 ;
        RECT 32.800 87.800 33.200 88.200 ;
        RECT 33.400 87.800 33.800 88.200 ;
        RECT 60.200 87.800 60.600 88.200 ;
        RECT 60.800 87.800 61.200 88.200 ;
        RECT 61.400 87.800 61.800 88.200 ;
        RECT 88.200 87.800 88.600 88.200 ;
        RECT 88.800 87.800 89.200 88.200 ;
        RECT 89.400 87.800 89.800 88.200 ;
        RECT 116.200 87.800 116.600 88.200 ;
        RECT 116.800 87.800 117.200 88.200 ;
        RECT 117.400 87.800 117.800 88.200 ;
        RECT 4.200 87.200 4.600 87.600 ;
        RECT 4.800 87.200 5.200 87.600 ;
        RECT 5.400 87.200 5.800 87.600 ;
        RECT 32.200 87.200 32.600 87.600 ;
        RECT 32.800 87.200 33.200 87.600 ;
        RECT 33.400 87.200 33.800 87.600 ;
        RECT 60.200 87.200 60.600 87.600 ;
        RECT 60.800 87.200 61.200 87.600 ;
        RECT 61.400 87.200 61.800 87.600 ;
        RECT 88.200 87.200 88.600 87.600 ;
        RECT 88.800 87.200 89.200 87.600 ;
        RECT 89.400 87.200 89.800 87.600 ;
        RECT 116.200 87.200 116.600 87.600 ;
        RECT 116.800 87.200 117.200 87.600 ;
        RECT 117.400 87.200 117.800 87.600 ;
        RECT 32.160 56.670 32.520 57.035 ;
        RECT 32.600 56.670 32.960 57.035 ;
        RECT 33.040 56.670 33.400 57.035 ;
        RECT 33.480 56.670 33.840 57.035 ;
        RECT 60.160 56.670 60.520 57.035 ;
        RECT 60.600 56.670 60.960 57.035 ;
        RECT 61.040 56.670 61.400 57.035 ;
        RECT 61.480 56.670 61.840 57.035 ;
        RECT 88.160 56.670 88.520 57.035 ;
        RECT 88.600 56.670 88.960 57.035 ;
        RECT 89.040 56.670 89.400 57.035 ;
        RECT 89.480 56.670 89.840 57.035 ;
        RECT 116.160 50.020 116.520 50.385 ;
        RECT 116.600 50.020 116.960 50.385 ;
        RECT 117.040 50.020 117.400 50.385 ;
        RECT 117.480 50.020 117.840 50.385 ;
        RECT 4.160 48.620 4.520 48.985 ;
        RECT 4.600 48.620 4.960 48.985 ;
        RECT 5.040 48.620 5.400 48.985 ;
        RECT 5.480 48.620 5.840 48.985 ;
        RECT 32.160 24.870 32.520 25.235 ;
        RECT 32.600 24.870 32.960 25.235 ;
        RECT 33.040 24.870 33.400 25.235 ;
        RECT 33.480 24.870 33.840 25.235 ;
        RECT 60.160 24.870 60.520 25.235 ;
        RECT 60.600 24.870 60.960 25.235 ;
        RECT 61.040 24.870 61.400 25.235 ;
        RECT 61.480 24.870 61.840 25.235 ;
        RECT 4.200 -6.600 4.600 -6.200 ;
        RECT 4.800 -6.600 5.200 -6.200 ;
        RECT 5.400 -6.600 5.800 -6.200 ;
        RECT 32.200 -6.600 32.600 -6.200 ;
        RECT 32.800 -6.600 33.200 -6.200 ;
        RECT 33.400 -6.600 33.800 -6.200 ;
        RECT 60.200 -6.600 60.600 -6.200 ;
        RECT 60.800 -6.600 61.200 -6.200 ;
        RECT 61.400 -6.600 61.800 -6.200 ;
        RECT 88.200 -6.600 88.600 -6.200 ;
        RECT 88.800 -6.600 89.200 -6.200 ;
        RECT 89.400 -6.600 89.800 -6.200 ;
        RECT 116.200 -6.600 116.600 -6.200 ;
        RECT 116.800 -6.600 117.200 -6.200 ;
        RECT 117.400 -6.600 117.800 -6.200 ;
        RECT 4.200 -7.200 4.600 -6.800 ;
        RECT 4.800 -7.200 5.200 -6.800 ;
        RECT 5.400 -7.200 5.800 -6.800 ;
        RECT 32.200 -7.200 32.600 -6.800 ;
        RECT 32.800 -7.200 33.200 -6.800 ;
        RECT 33.400 -7.200 33.800 -6.800 ;
        RECT 60.200 -7.200 60.600 -6.800 ;
        RECT 60.800 -7.200 61.200 -6.800 ;
        RECT 61.400 -7.200 61.800 -6.800 ;
        RECT 88.200 -7.200 88.600 -6.800 ;
        RECT 88.800 -7.200 89.200 -6.800 ;
        RECT 89.400 -7.200 89.800 -6.800 ;
        RECT 116.200 -7.200 116.600 -6.800 ;
        RECT 116.800 -7.200 117.200 -6.800 ;
        RECT 117.400 -7.200 117.800 -6.800 ;
        RECT 4.200 -7.800 4.600 -7.400 ;
        RECT 4.800 -7.800 5.200 -7.400 ;
        RECT 5.400 -7.800 5.800 -7.400 ;
        RECT 32.200 -7.800 32.600 -7.400 ;
        RECT 32.800 -7.800 33.200 -7.400 ;
        RECT 33.400 -7.800 33.800 -7.400 ;
        RECT 60.200 -7.800 60.600 -7.400 ;
        RECT 60.800 -7.800 61.200 -7.400 ;
        RECT 61.400 -7.800 61.800 -7.400 ;
        RECT 88.200 -7.800 88.600 -7.400 ;
        RECT 88.800 -7.800 89.200 -7.400 ;
        RECT 89.400 -7.800 89.800 -7.400 ;
        RECT 116.200 -7.800 116.600 -7.400 ;
        RECT 116.800 -7.800 117.200 -7.400 ;
        RECT 117.400 -7.800 117.800 -7.400 ;
      LAYER met4 ;
        RECT 4.000 -8.000 6.000 89.000 ;
        RECT 32.000 -8.000 34.000 89.000 ;
        RECT 60.000 -8.000 62.000 89.000 ;
        RECT 88.000 -8.000 90.000 89.000 ;
        RECT 116.000 -8.000 118.000 89.000 ;
    END
  END vssd2
  OBS
      LAYER pwell ;
        RECT 6.840 48.715 7.010 48.885 ;
        RECT 10.830 48.715 11.000 48.885 ;
        RECT 15.980 41.470 105.050 48.570 ;
        RECT 108.000 46.000 111.000 51.000 ;
        RECT 108.000 45.000 116.000 46.000 ;
        RECT 110.000 43.000 116.000 45.000 ;
        RECT 7.500 33.270 114.280 40.370 ;
      LAYER li1 ;
        RECT 6.775 50.865 7.035 51.265 ;
        RECT 6.775 50.695 8.140 50.865 ;
        RECT 7.405 49.625 8.140 50.695 ;
        RECT 8.665 50.750 8.905 50.755 ;
        RECT 9.180 50.750 10.505 50.960 ;
        RECT 8.665 50.740 10.505 50.750 ;
        RECT 8.665 50.530 9.400 50.740 ;
        RECT 10.285 50.535 10.505 50.740 ;
        RECT 10.770 50.535 11.290 50.540 ;
        RECT 8.665 49.775 8.905 50.530 ;
        RECT 10.285 50.315 11.290 50.535 ;
        RECT 6.775 49.455 8.140 49.625 ;
        RECT 6.775 49.055 7.035 49.455 ;
        RECT 10.770 49.055 11.290 50.315 ;
        RECT 11.460 49.715 11.980 51.265 ;
        RECT 23.400 48.950 23.780 49.000 ;
        RECT 22.450 48.590 23.780 48.950 ;
        RECT 23.400 48.540 23.780 48.590 ;
        RECT 16.670 42.090 16.960 47.540 ;
        RECT 21.050 42.090 21.340 47.540 ;
        RECT 22.190 42.090 22.480 47.540 ;
        RECT 24.375 42.500 24.675 55.090 ;
        RECT 25.270 48.950 25.650 49.000 ;
        RECT 25.270 48.590 26.600 48.950 ;
        RECT 25.270 48.540 25.650 48.590 ;
        RECT 26.570 42.090 26.860 47.540 ;
        RECT 27.710 42.090 28.000 47.540 ;
        RECT 29.900 42.500 30.200 55.090 ;
        RECT 32.250 48.950 32.630 49.000 ;
        RECT 41.110 48.950 41.490 49.000 ;
        RECT 31.300 48.590 32.630 48.950 ;
        RECT 40.160 48.590 41.490 48.950 ;
        RECT 32.250 48.540 32.630 48.590 ;
        RECT 41.110 48.540 41.490 48.590 ;
        RECT 31.040 42.090 31.330 47.540 ;
        RECT 34.380 42.090 34.670 47.540 ;
        RECT 38.760 42.090 39.050 47.540 ;
        RECT 39.900 42.090 40.190 47.540 ;
        RECT 42.085 42.500 42.385 55.090 ;
        RECT 42.980 48.950 43.360 49.000 ;
        RECT 42.980 48.590 44.310 48.950 ;
        RECT 42.980 48.540 43.360 48.590 ;
        RECT 44.280 42.090 44.570 47.540 ;
        RECT 45.420 42.090 45.710 47.540 ;
        RECT 47.610 42.500 47.910 55.090 ;
        RECT 49.960 48.950 50.340 49.000 ;
        RECT 58.820 48.950 59.200 49.000 ;
        RECT 49.010 48.590 50.340 48.950 ;
        RECT 57.870 48.590 59.200 48.950 ;
        RECT 49.960 48.540 50.340 48.590 ;
        RECT 58.820 48.540 59.200 48.590 ;
        RECT 48.750 42.090 49.040 47.540 ;
        RECT 52.090 42.090 52.380 47.540 ;
        RECT 56.470 42.090 56.760 47.540 ;
        RECT 57.610 42.090 57.900 47.540 ;
        RECT 59.795 42.500 60.095 55.090 ;
        RECT 60.690 48.950 61.070 49.000 ;
        RECT 60.690 48.590 62.020 48.950 ;
        RECT 60.690 48.540 61.070 48.590 ;
        RECT 61.990 42.090 62.280 47.540 ;
        RECT 63.130 42.090 63.420 47.540 ;
        RECT 65.320 42.500 65.620 55.090 ;
        RECT 67.670 48.950 68.050 49.000 ;
        RECT 76.530 48.950 76.910 49.000 ;
        RECT 66.720 48.590 68.050 48.950 ;
        RECT 75.580 48.590 76.910 48.950 ;
        RECT 67.670 48.540 68.050 48.590 ;
        RECT 76.530 48.540 76.910 48.590 ;
        RECT 66.460 42.090 66.750 47.540 ;
        RECT 69.800 42.090 70.090 47.540 ;
        RECT 74.180 42.090 74.470 47.540 ;
        RECT 75.320 42.090 75.610 47.540 ;
        RECT 77.505 42.500 77.805 55.090 ;
        RECT 78.400 48.950 78.780 49.000 ;
        RECT 78.400 48.590 79.730 48.950 ;
        RECT 78.400 48.540 78.780 48.590 ;
        RECT 79.700 42.090 79.990 47.540 ;
        RECT 80.840 42.090 81.130 47.540 ;
        RECT 83.030 42.500 83.330 55.090 ;
        RECT 85.380 48.950 85.760 49.000 ;
        RECT 94.240 48.950 94.620 49.000 ;
        RECT 84.430 48.590 85.760 48.950 ;
        RECT 93.290 48.590 94.620 48.950 ;
        RECT 85.380 48.540 85.760 48.590 ;
        RECT 94.240 48.540 94.620 48.590 ;
        RECT 84.170 42.090 84.460 47.540 ;
        RECT 87.510 42.090 87.800 47.540 ;
        RECT 91.890 42.090 92.180 47.540 ;
        RECT 93.030 42.090 93.320 47.540 ;
        RECT 95.215 42.500 95.515 55.090 ;
        RECT 96.110 48.950 96.490 49.000 ;
        RECT 96.110 48.590 97.440 48.950 ;
        RECT 96.110 48.540 96.490 48.590 ;
        RECT 97.410 42.090 97.700 47.540 ;
        RECT 98.550 42.090 98.840 47.540 ;
        RECT 100.740 42.500 101.040 55.090 ;
        RECT 103.090 48.950 103.470 49.000 ;
        RECT 102.140 48.590 103.470 48.950 ;
        RECT 103.090 48.540 103.470 48.590 ;
        RECT 101.880 42.090 102.170 47.540 ;
        RECT 108.500 45.500 110.500 45.865 ;
        RECT 109.500 44.500 110.865 45.500 ;
        RECT 110.500 43.500 110.865 44.500 ;
        RECT 16.160 41.730 18.050 42.090 ;
        RECT 19.840 41.730 23.690 42.090 ;
        RECT 25.350 41.730 29.200 42.090 ;
        RECT 31.040 41.730 32.440 42.090 ;
        RECT 33.870 41.730 35.760 42.090 ;
        RECT 37.550 41.730 41.400 42.090 ;
        RECT 43.060 41.730 46.910 42.090 ;
        RECT 48.750 41.730 50.150 42.090 ;
        RECT 51.580 41.730 53.470 42.090 ;
        RECT 55.260 41.730 59.110 42.090 ;
        RECT 60.770 41.730 64.620 42.090 ;
        RECT 66.460 41.730 67.860 42.090 ;
        RECT 69.290 41.730 71.180 42.090 ;
        RECT 72.970 41.730 76.820 42.090 ;
        RECT 78.480 41.730 82.330 42.090 ;
        RECT 84.170 41.730 85.570 42.090 ;
        RECT 87.000 41.730 88.890 42.090 ;
        RECT 90.680 41.730 94.530 42.090 ;
        RECT 96.190 41.730 100.040 42.090 ;
        RECT 101.880 41.730 103.280 42.090 ;
        RECT 9.270 39.750 10.670 40.110 ;
        RECT 12.510 39.750 16.360 40.110 ;
        RECT 18.020 39.750 21.870 40.110 ;
        RECT 23.660 39.750 25.550 40.110 ;
        RECT 26.980 39.750 28.380 40.110 ;
        RECT 30.220 39.750 34.070 40.110 ;
        RECT 35.730 39.750 39.580 40.110 ;
        RECT 41.370 39.750 43.260 40.110 ;
        RECT 44.690 39.750 46.090 40.110 ;
        RECT 47.930 39.750 51.780 40.110 ;
        RECT 53.440 39.750 57.290 40.110 ;
        RECT 59.080 39.750 60.970 40.110 ;
        RECT 62.400 39.750 63.800 40.110 ;
        RECT 65.640 39.750 69.490 40.110 ;
        RECT 71.150 39.750 75.000 40.110 ;
        RECT 76.790 39.750 78.680 40.110 ;
        RECT 80.110 39.750 81.510 40.110 ;
        RECT 83.350 39.750 87.200 40.110 ;
        RECT 88.860 39.750 92.710 40.110 ;
        RECT 94.500 39.750 96.390 40.110 ;
        RECT 97.820 39.750 99.220 40.110 ;
        RECT 101.060 39.750 104.910 40.110 ;
        RECT 106.570 39.750 110.420 40.110 ;
        RECT 112.210 39.750 114.100 40.110 ;
        RECT 10.380 34.300 10.670 39.750 ;
        RECT 9.080 33.250 9.460 33.300 ;
        RECT 9.080 32.890 10.410 33.250 ;
        RECT 9.080 32.840 9.460 32.890 ;
        RECT 11.510 26.750 11.810 39.340 ;
        RECT 13.710 34.300 14.000 39.750 ;
        RECT 14.850 34.300 15.140 39.750 ;
        RECT 16.060 33.250 16.440 33.300 ;
        RECT 15.110 32.890 16.440 33.250 ;
        RECT 16.060 32.840 16.440 32.890 ;
        RECT 17.035 26.750 17.335 39.340 ;
        RECT 19.230 34.300 19.520 39.750 ;
        RECT 20.370 34.300 20.660 39.750 ;
        RECT 24.750 34.300 25.040 39.750 ;
        RECT 28.090 34.300 28.380 39.750 ;
        RECT 17.930 33.250 18.310 33.300 ;
        RECT 26.790 33.250 27.170 33.300 ;
        RECT 17.930 32.890 19.260 33.250 ;
        RECT 26.790 32.890 28.120 33.250 ;
        RECT 17.930 32.840 18.310 32.890 ;
        RECT 26.790 32.840 27.170 32.890 ;
        RECT 29.220 26.750 29.520 39.340 ;
        RECT 31.420 34.300 31.710 39.750 ;
        RECT 32.560 34.300 32.850 39.750 ;
        RECT 33.770 33.250 34.150 33.300 ;
        RECT 32.820 32.890 34.150 33.250 ;
        RECT 33.770 32.840 34.150 32.890 ;
        RECT 34.745 26.750 35.045 39.340 ;
        RECT 36.940 34.300 37.230 39.750 ;
        RECT 38.080 34.300 38.370 39.750 ;
        RECT 42.460 34.300 42.750 39.750 ;
        RECT 45.800 34.300 46.090 39.750 ;
        RECT 35.640 33.250 36.020 33.300 ;
        RECT 44.500 33.250 44.880 33.300 ;
        RECT 35.640 32.890 36.970 33.250 ;
        RECT 44.500 32.890 45.830 33.250 ;
        RECT 35.640 32.840 36.020 32.890 ;
        RECT 44.500 32.840 44.880 32.890 ;
        RECT 46.930 26.750 47.230 39.340 ;
        RECT 49.130 34.300 49.420 39.750 ;
        RECT 50.270 34.300 50.560 39.750 ;
        RECT 51.480 33.250 51.860 33.300 ;
        RECT 50.530 32.890 51.860 33.250 ;
        RECT 51.480 32.840 51.860 32.890 ;
        RECT 52.455 26.750 52.755 39.340 ;
        RECT 54.650 34.300 54.940 39.750 ;
        RECT 55.790 34.300 56.080 39.750 ;
        RECT 60.170 34.300 60.460 39.750 ;
        RECT 63.510 34.300 63.800 39.750 ;
        RECT 53.350 33.250 53.730 33.300 ;
        RECT 62.210 33.250 62.590 33.300 ;
        RECT 53.350 32.890 54.680 33.250 ;
        RECT 62.210 32.890 63.540 33.250 ;
        RECT 53.350 32.840 53.730 32.890 ;
        RECT 62.210 32.840 62.590 32.890 ;
        RECT 64.640 26.750 64.940 39.340 ;
        RECT 66.840 34.300 67.130 39.750 ;
        RECT 67.980 34.300 68.270 39.750 ;
        RECT 69.190 33.250 69.570 33.300 ;
        RECT 68.240 32.890 69.570 33.250 ;
        RECT 69.190 32.840 69.570 32.890 ;
        RECT 70.165 26.750 70.465 39.340 ;
        RECT 72.360 34.300 72.650 39.750 ;
        RECT 73.500 34.300 73.790 39.750 ;
        RECT 77.880 34.300 78.170 39.750 ;
        RECT 81.220 34.300 81.510 39.750 ;
        RECT 71.060 33.250 71.440 33.300 ;
        RECT 79.920 33.250 80.300 33.300 ;
        RECT 71.060 32.890 72.390 33.250 ;
        RECT 79.920 32.890 81.250 33.250 ;
        RECT 71.060 32.840 71.440 32.890 ;
        RECT 79.920 32.840 80.300 32.890 ;
        RECT 82.350 26.750 82.650 39.340 ;
        RECT 84.550 34.300 84.840 39.750 ;
        RECT 85.690 34.300 85.980 39.750 ;
        RECT 86.900 33.250 87.280 33.300 ;
        RECT 85.950 32.890 87.280 33.250 ;
        RECT 86.900 32.840 87.280 32.890 ;
        RECT 87.875 26.750 88.175 39.340 ;
        RECT 90.070 34.300 90.360 39.750 ;
        RECT 91.210 34.300 91.500 39.750 ;
        RECT 95.590 34.300 95.880 39.750 ;
        RECT 98.930 34.300 99.220 39.750 ;
        RECT 88.770 33.250 89.150 33.300 ;
        RECT 97.630 33.250 98.010 33.300 ;
        RECT 88.770 32.890 90.100 33.250 ;
        RECT 97.630 32.890 98.960 33.250 ;
        RECT 88.770 32.840 89.150 32.890 ;
        RECT 97.630 32.840 98.010 32.890 ;
        RECT 100.060 26.750 100.360 39.340 ;
        RECT 102.260 34.300 102.550 39.750 ;
        RECT 103.400 34.300 103.690 39.750 ;
        RECT 104.610 33.250 104.990 33.300 ;
        RECT 103.660 32.890 104.990 33.250 ;
        RECT 104.610 32.840 104.990 32.890 ;
        RECT 105.585 26.750 105.885 39.340 ;
        RECT 107.780 34.300 108.070 39.750 ;
        RECT 108.920 34.300 109.210 39.750 ;
        RECT 113.300 34.300 113.590 39.750 ;
        RECT 106.480 33.250 106.860 33.300 ;
        RECT 106.480 32.890 107.810 33.250 ;
        RECT 106.480 32.840 106.860 32.890 ;
      LAYER mcon ;
        RECT 22.450 48.620 22.750 48.920 ;
        RECT 22.940 48.620 23.240 48.920 ;
        RECT 23.430 48.620 23.730 48.920 ;
        RECT 25.320 48.620 25.620 48.920 ;
        RECT 25.810 48.620 26.110 48.920 ;
        RECT 26.300 48.620 26.600 48.920 ;
        RECT 24.375 47.260 24.675 47.560 ;
        RECT 31.300 48.620 31.600 48.920 ;
        RECT 31.790 48.620 32.090 48.920 ;
        RECT 32.280 48.620 32.580 48.920 ;
        RECT 40.160 48.620 40.460 48.920 ;
        RECT 40.650 48.620 40.950 48.920 ;
        RECT 41.140 48.620 41.440 48.920 ;
        RECT 29.900 47.260 30.200 47.560 ;
        RECT 43.030 48.620 43.330 48.920 ;
        RECT 43.520 48.620 43.820 48.920 ;
        RECT 44.010 48.620 44.310 48.920 ;
        RECT 42.085 47.260 42.385 47.560 ;
        RECT 49.010 48.620 49.310 48.920 ;
        RECT 49.500 48.620 49.800 48.920 ;
        RECT 49.990 48.620 50.290 48.920 ;
        RECT 57.870 48.620 58.170 48.920 ;
        RECT 58.360 48.620 58.660 48.920 ;
        RECT 58.850 48.620 59.150 48.920 ;
        RECT 47.610 47.260 47.910 47.560 ;
        RECT 60.740 48.620 61.040 48.920 ;
        RECT 61.230 48.620 61.530 48.920 ;
        RECT 61.720 48.620 62.020 48.920 ;
        RECT 59.795 47.260 60.095 47.560 ;
        RECT 66.720 48.620 67.020 48.920 ;
        RECT 67.210 48.620 67.510 48.920 ;
        RECT 67.700 48.620 68.000 48.920 ;
        RECT 75.580 48.620 75.880 48.920 ;
        RECT 76.070 48.620 76.370 48.920 ;
        RECT 76.560 48.620 76.860 48.920 ;
        RECT 65.320 47.260 65.620 47.560 ;
        RECT 78.450 48.620 78.750 48.920 ;
        RECT 78.940 48.620 79.240 48.920 ;
        RECT 79.430 48.620 79.730 48.920 ;
        RECT 77.505 47.260 77.805 47.560 ;
        RECT 84.430 48.620 84.730 48.920 ;
        RECT 84.920 48.620 85.220 48.920 ;
        RECT 85.410 48.620 85.710 48.920 ;
        RECT 93.290 48.620 93.590 48.920 ;
        RECT 93.780 48.620 94.080 48.920 ;
        RECT 94.270 48.620 94.570 48.920 ;
        RECT 83.030 47.260 83.330 47.560 ;
        RECT 96.160 48.620 96.460 48.920 ;
        RECT 96.650 48.620 96.950 48.920 ;
        RECT 97.140 48.620 97.440 48.920 ;
        RECT 95.215 47.260 95.515 47.560 ;
        RECT 102.140 48.620 102.440 48.920 ;
        RECT 102.630 48.620 102.930 48.920 ;
        RECT 103.120 48.620 103.420 48.920 ;
        RECT 100.740 47.260 101.040 47.560 ;
        RECT 109.590 45.120 109.890 45.420 ;
        RECT 110.110 45.120 110.410 45.420 ;
        RECT 109.590 44.600 109.890 44.900 ;
        RECT 110.110 44.600 110.410 44.900 ;
        RECT 16.220 41.760 16.520 42.060 ;
        RECT 16.710 41.760 17.010 42.060 ;
        RECT 17.200 41.760 17.500 42.060 ;
        RECT 17.690 41.760 17.990 42.060 ;
        RECT 19.900 41.760 20.200 42.060 ;
        RECT 20.390 41.760 20.690 42.060 ;
        RECT 20.880 41.760 21.180 42.060 ;
        RECT 21.370 41.760 21.670 42.060 ;
        RECT 21.860 41.760 22.160 42.060 ;
        RECT 22.350 41.760 22.650 42.060 ;
        RECT 22.840 41.760 23.140 42.060 ;
        RECT 23.330 41.760 23.630 42.060 ;
        RECT 25.410 41.760 25.710 42.060 ;
        RECT 25.900 41.760 26.200 42.060 ;
        RECT 26.390 41.760 26.690 42.060 ;
        RECT 26.880 41.760 27.180 42.060 ;
        RECT 27.370 41.760 27.670 42.060 ;
        RECT 27.860 41.760 28.160 42.060 ;
        RECT 28.350 41.760 28.650 42.060 ;
        RECT 28.840 41.760 29.140 42.060 ;
        RECT 31.100 41.760 31.400 42.060 ;
        RECT 31.590 41.760 31.890 42.060 ;
        RECT 32.080 41.760 32.380 42.060 ;
        RECT 33.930 41.760 34.230 42.060 ;
        RECT 34.420 41.760 34.720 42.060 ;
        RECT 34.910 41.760 35.210 42.060 ;
        RECT 35.400 41.760 35.700 42.060 ;
        RECT 37.610 41.760 37.910 42.060 ;
        RECT 38.100 41.760 38.400 42.060 ;
        RECT 38.590 41.760 38.890 42.060 ;
        RECT 39.080 41.760 39.380 42.060 ;
        RECT 39.570 41.760 39.870 42.060 ;
        RECT 40.060 41.760 40.360 42.060 ;
        RECT 40.550 41.760 40.850 42.060 ;
        RECT 41.040 41.760 41.340 42.060 ;
        RECT 43.120 41.760 43.420 42.060 ;
        RECT 43.610 41.760 43.910 42.060 ;
        RECT 44.100 41.760 44.400 42.060 ;
        RECT 44.590 41.760 44.890 42.060 ;
        RECT 45.080 41.760 45.380 42.060 ;
        RECT 45.570 41.760 45.870 42.060 ;
        RECT 46.060 41.760 46.360 42.060 ;
        RECT 46.550 41.760 46.850 42.060 ;
        RECT 48.810 41.760 49.110 42.060 ;
        RECT 49.300 41.760 49.600 42.060 ;
        RECT 49.790 41.760 50.090 42.060 ;
        RECT 51.640 41.760 51.940 42.060 ;
        RECT 52.130 41.760 52.430 42.060 ;
        RECT 52.620 41.760 52.920 42.060 ;
        RECT 53.110 41.760 53.410 42.060 ;
        RECT 55.320 41.760 55.620 42.060 ;
        RECT 55.810 41.760 56.110 42.060 ;
        RECT 56.300 41.760 56.600 42.060 ;
        RECT 56.790 41.760 57.090 42.060 ;
        RECT 57.280 41.760 57.580 42.060 ;
        RECT 57.770 41.760 58.070 42.060 ;
        RECT 58.260 41.760 58.560 42.060 ;
        RECT 58.750 41.760 59.050 42.060 ;
        RECT 60.830 41.760 61.130 42.060 ;
        RECT 61.320 41.760 61.620 42.060 ;
        RECT 61.810 41.760 62.110 42.060 ;
        RECT 62.300 41.760 62.600 42.060 ;
        RECT 62.790 41.760 63.090 42.060 ;
        RECT 63.280 41.760 63.580 42.060 ;
        RECT 63.770 41.760 64.070 42.060 ;
        RECT 64.260 41.760 64.560 42.060 ;
        RECT 66.520 41.760 66.820 42.060 ;
        RECT 67.010 41.760 67.310 42.060 ;
        RECT 67.500 41.760 67.800 42.060 ;
        RECT 69.350 41.760 69.650 42.060 ;
        RECT 69.840 41.760 70.140 42.060 ;
        RECT 70.330 41.760 70.630 42.060 ;
        RECT 70.820 41.760 71.120 42.060 ;
        RECT 73.030 41.760 73.330 42.060 ;
        RECT 73.520 41.760 73.820 42.060 ;
        RECT 74.010 41.760 74.310 42.060 ;
        RECT 74.500 41.760 74.800 42.060 ;
        RECT 74.990 41.760 75.290 42.060 ;
        RECT 75.480 41.760 75.780 42.060 ;
        RECT 75.970 41.760 76.270 42.060 ;
        RECT 76.460 41.760 76.760 42.060 ;
        RECT 78.540 41.760 78.840 42.060 ;
        RECT 79.030 41.760 79.330 42.060 ;
        RECT 79.520 41.760 79.820 42.060 ;
        RECT 80.010 41.760 80.310 42.060 ;
        RECT 80.500 41.760 80.800 42.060 ;
        RECT 80.990 41.760 81.290 42.060 ;
        RECT 81.480 41.760 81.780 42.060 ;
        RECT 81.970 41.760 82.270 42.060 ;
        RECT 84.230 41.760 84.530 42.060 ;
        RECT 84.720 41.760 85.020 42.060 ;
        RECT 85.210 41.760 85.510 42.060 ;
        RECT 87.060 41.760 87.360 42.060 ;
        RECT 87.550 41.760 87.850 42.060 ;
        RECT 88.040 41.760 88.340 42.060 ;
        RECT 88.530 41.760 88.830 42.060 ;
        RECT 90.740 41.760 91.040 42.060 ;
        RECT 91.230 41.760 91.530 42.060 ;
        RECT 91.720 41.760 92.020 42.060 ;
        RECT 92.210 41.760 92.510 42.060 ;
        RECT 92.700 41.760 93.000 42.060 ;
        RECT 93.190 41.760 93.490 42.060 ;
        RECT 93.680 41.760 93.980 42.060 ;
        RECT 94.170 41.760 94.470 42.060 ;
        RECT 96.250 41.760 96.550 42.060 ;
        RECT 96.740 41.760 97.040 42.060 ;
        RECT 97.230 41.760 97.530 42.060 ;
        RECT 97.720 41.760 98.020 42.060 ;
        RECT 98.210 41.760 98.510 42.060 ;
        RECT 98.700 41.760 99.000 42.060 ;
        RECT 99.190 41.760 99.490 42.060 ;
        RECT 99.680 41.760 99.980 42.060 ;
        RECT 101.940 41.760 102.240 42.060 ;
        RECT 102.430 41.760 102.730 42.060 ;
        RECT 102.920 41.760 103.220 42.060 ;
        RECT 9.330 39.780 9.630 40.080 ;
        RECT 9.820 39.780 10.120 40.080 ;
        RECT 10.310 39.780 10.610 40.080 ;
        RECT 12.570 39.780 12.870 40.080 ;
        RECT 13.060 39.780 13.360 40.080 ;
        RECT 13.550 39.780 13.850 40.080 ;
        RECT 14.040 39.780 14.340 40.080 ;
        RECT 14.530 39.780 14.830 40.080 ;
        RECT 15.020 39.780 15.320 40.080 ;
        RECT 15.510 39.780 15.810 40.080 ;
        RECT 16.000 39.780 16.300 40.080 ;
        RECT 18.080 39.780 18.380 40.080 ;
        RECT 18.570 39.780 18.870 40.080 ;
        RECT 19.060 39.780 19.360 40.080 ;
        RECT 19.550 39.780 19.850 40.080 ;
        RECT 20.040 39.780 20.340 40.080 ;
        RECT 20.530 39.780 20.830 40.080 ;
        RECT 21.020 39.780 21.320 40.080 ;
        RECT 21.510 39.780 21.810 40.080 ;
        RECT 23.720 39.780 24.020 40.080 ;
        RECT 24.210 39.780 24.510 40.080 ;
        RECT 24.700 39.780 25.000 40.080 ;
        RECT 25.190 39.780 25.490 40.080 ;
        RECT 27.040 39.780 27.340 40.080 ;
        RECT 27.530 39.780 27.830 40.080 ;
        RECT 28.020 39.780 28.320 40.080 ;
        RECT 30.280 39.780 30.580 40.080 ;
        RECT 30.770 39.780 31.070 40.080 ;
        RECT 31.260 39.780 31.560 40.080 ;
        RECT 31.750 39.780 32.050 40.080 ;
        RECT 32.240 39.780 32.540 40.080 ;
        RECT 32.730 39.780 33.030 40.080 ;
        RECT 33.220 39.780 33.520 40.080 ;
        RECT 33.710 39.780 34.010 40.080 ;
        RECT 35.790 39.780 36.090 40.080 ;
        RECT 36.280 39.780 36.580 40.080 ;
        RECT 36.770 39.780 37.070 40.080 ;
        RECT 37.260 39.780 37.560 40.080 ;
        RECT 37.750 39.780 38.050 40.080 ;
        RECT 38.240 39.780 38.540 40.080 ;
        RECT 38.730 39.780 39.030 40.080 ;
        RECT 39.220 39.780 39.520 40.080 ;
        RECT 41.430 39.780 41.730 40.080 ;
        RECT 41.920 39.780 42.220 40.080 ;
        RECT 42.410 39.780 42.710 40.080 ;
        RECT 42.900 39.780 43.200 40.080 ;
        RECT 44.750 39.780 45.050 40.080 ;
        RECT 45.240 39.780 45.540 40.080 ;
        RECT 45.730 39.780 46.030 40.080 ;
        RECT 47.990 39.780 48.290 40.080 ;
        RECT 48.480 39.780 48.780 40.080 ;
        RECT 48.970 39.780 49.270 40.080 ;
        RECT 49.460 39.780 49.760 40.080 ;
        RECT 49.950 39.780 50.250 40.080 ;
        RECT 50.440 39.780 50.740 40.080 ;
        RECT 50.930 39.780 51.230 40.080 ;
        RECT 51.420 39.780 51.720 40.080 ;
        RECT 53.500 39.780 53.800 40.080 ;
        RECT 53.990 39.780 54.290 40.080 ;
        RECT 54.480 39.780 54.780 40.080 ;
        RECT 54.970 39.780 55.270 40.080 ;
        RECT 55.460 39.780 55.760 40.080 ;
        RECT 55.950 39.780 56.250 40.080 ;
        RECT 56.440 39.780 56.740 40.080 ;
        RECT 56.930 39.780 57.230 40.080 ;
        RECT 59.140 39.780 59.440 40.080 ;
        RECT 59.630 39.780 59.930 40.080 ;
        RECT 60.120 39.780 60.420 40.080 ;
        RECT 60.610 39.780 60.910 40.080 ;
        RECT 62.460 39.780 62.760 40.080 ;
        RECT 62.950 39.780 63.250 40.080 ;
        RECT 63.440 39.780 63.740 40.080 ;
        RECT 65.700 39.780 66.000 40.080 ;
        RECT 66.190 39.780 66.490 40.080 ;
        RECT 66.680 39.780 66.980 40.080 ;
        RECT 67.170 39.780 67.470 40.080 ;
        RECT 67.660 39.780 67.960 40.080 ;
        RECT 68.150 39.780 68.450 40.080 ;
        RECT 68.640 39.780 68.940 40.080 ;
        RECT 69.130 39.780 69.430 40.080 ;
        RECT 71.210 39.780 71.510 40.080 ;
        RECT 71.700 39.780 72.000 40.080 ;
        RECT 72.190 39.780 72.490 40.080 ;
        RECT 72.680 39.780 72.980 40.080 ;
        RECT 73.170 39.780 73.470 40.080 ;
        RECT 73.660 39.780 73.960 40.080 ;
        RECT 74.150 39.780 74.450 40.080 ;
        RECT 74.640 39.780 74.940 40.080 ;
        RECT 76.850 39.780 77.150 40.080 ;
        RECT 77.340 39.780 77.640 40.080 ;
        RECT 77.830 39.780 78.130 40.080 ;
        RECT 78.320 39.780 78.620 40.080 ;
        RECT 80.170 39.780 80.470 40.080 ;
        RECT 80.660 39.780 80.960 40.080 ;
        RECT 81.150 39.780 81.450 40.080 ;
        RECT 83.410 39.780 83.710 40.080 ;
        RECT 83.900 39.780 84.200 40.080 ;
        RECT 84.390 39.780 84.690 40.080 ;
        RECT 84.880 39.780 85.180 40.080 ;
        RECT 85.370 39.780 85.670 40.080 ;
        RECT 85.860 39.780 86.160 40.080 ;
        RECT 86.350 39.780 86.650 40.080 ;
        RECT 86.840 39.780 87.140 40.080 ;
        RECT 88.920 39.780 89.220 40.080 ;
        RECT 89.410 39.780 89.710 40.080 ;
        RECT 89.900 39.780 90.200 40.080 ;
        RECT 90.390 39.780 90.690 40.080 ;
        RECT 90.880 39.780 91.180 40.080 ;
        RECT 91.370 39.780 91.670 40.080 ;
        RECT 91.860 39.780 92.160 40.080 ;
        RECT 92.350 39.780 92.650 40.080 ;
        RECT 94.560 39.780 94.860 40.080 ;
        RECT 95.050 39.780 95.350 40.080 ;
        RECT 95.540 39.780 95.840 40.080 ;
        RECT 96.030 39.780 96.330 40.080 ;
        RECT 97.880 39.780 98.180 40.080 ;
        RECT 98.370 39.780 98.670 40.080 ;
        RECT 98.860 39.780 99.160 40.080 ;
        RECT 101.120 39.780 101.420 40.080 ;
        RECT 101.610 39.780 101.910 40.080 ;
        RECT 102.100 39.780 102.400 40.080 ;
        RECT 102.590 39.780 102.890 40.080 ;
        RECT 103.080 39.780 103.380 40.080 ;
        RECT 103.570 39.780 103.870 40.080 ;
        RECT 104.060 39.780 104.360 40.080 ;
        RECT 104.550 39.780 104.850 40.080 ;
        RECT 106.630 39.780 106.930 40.080 ;
        RECT 107.120 39.780 107.420 40.080 ;
        RECT 107.610 39.780 107.910 40.080 ;
        RECT 108.100 39.780 108.400 40.080 ;
        RECT 108.590 39.780 108.890 40.080 ;
        RECT 109.080 39.780 109.380 40.080 ;
        RECT 109.570 39.780 109.870 40.080 ;
        RECT 110.060 39.780 110.360 40.080 ;
        RECT 112.270 39.780 112.570 40.080 ;
        RECT 112.760 39.780 113.060 40.080 ;
        RECT 113.250 39.780 113.550 40.080 ;
        RECT 113.740 39.780 114.040 40.080 ;
        RECT 11.510 34.280 11.810 34.580 ;
        RECT 9.130 32.920 9.430 33.220 ;
        RECT 9.620 32.920 9.920 33.220 ;
        RECT 10.110 32.920 10.410 33.220 ;
        RECT 17.035 34.280 17.335 34.580 ;
        RECT 15.110 32.920 15.410 33.220 ;
        RECT 15.600 32.920 15.900 33.220 ;
        RECT 16.090 32.920 16.390 33.220 ;
        RECT 29.220 34.280 29.520 34.580 ;
        RECT 17.980 32.920 18.280 33.220 ;
        RECT 18.470 32.920 18.770 33.220 ;
        RECT 18.960 32.920 19.260 33.220 ;
        RECT 26.840 32.920 27.140 33.220 ;
        RECT 27.330 32.920 27.630 33.220 ;
        RECT 27.820 32.920 28.120 33.220 ;
        RECT 34.745 34.280 35.045 34.580 ;
        RECT 32.820 32.920 33.120 33.220 ;
        RECT 33.310 32.920 33.610 33.220 ;
        RECT 33.800 32.920 34.100 33.220 ;
        RECT 46.930 34.280 47.230 34.580 ;
        RECT 35.690 32.920 35.990 33.220 ;
        RECT 36.180 32.920 36.480 33.220 ;
        RECT 36.670 32.920 36.970 33.220 ;
        RECT 44.550 32.920 44.850 33.220 ;
        RECT 45.040 32.920 45.340 33.220 ;
        RECT 45.530 32.920 45.830 33.220 ;
        RECT 52.455 34.280 52.755 34.580 ;
        RECT 50.530 32.920 50.830 33.220 ;
        RECT 51.020 32.920 51.320 33.220 ;
        RECT 51.510 32.920 51.810 33.220 ;
        RECT 64.640 34.280 64.940 34.580 ;
        RECT 53.400 32.920 53.700 33.220 ;
        RECT 53.890 32.920 54.190 33.220 ;
        RECT 54.380 32.920 54.680 33.220 ;
        RECT 62.260 32.920 62.560 33.220 ;
        RECT 62.750 32.920 63.050 33.220 ;
        RECT 63.240 32.920 63.540 33.220 ;
        RECT 70.165 34.280 70.465 34.580 ;
        RECT 68.240 32.920 68.540 33.220 ;
        RECT 68.730 32.920 69.030 33.220 ;
        RECT 69.220 32.920 69.520 33.220 ;
        RECT 82.350 34.280 82.650 34.580 ;
        RECT 71.110 32.920 71.410 33.220 ;
        RECT 71.600 32.920 71.900 33.220 ;
        RECT 72.090 32.920 72.390 33.220 ;
        RECT 79.970 32.920 80.270 33.220 ;
        RECT 80.460 32.920 80.760 33.220 ;
        RECT 80.950 32.920 81.250 33.220 ;
        RECT 87.875 34.280 88.175 34.580 ;
        RECT 85.950 32.920 86.250 33.220 ;
        RECT 86.440 32.920 86.740 33.220 ;
        RECT 86.930 32.920 87.230 33.220 ;
        RECT 100.060 34.280 100.360 34.580 ;
        RECT 88.820 32.920 89.120 33.220 ;
        RECT 89.310 32.920 89.610 33.220 ;
        RECT 89.800 32.920 90.100 33.220 ;
        RECT 97.680 32.920 97.980 33.220 ;
        RECT 98.170 32.920 98.470 33.220 ;
        RECT 98.660 32.920 98.960 33.220 ;
        RECT 105.585 34.280 105.885 34.580 ;
        RECT 103.660 32.920 103.960 33.220 ;
        RECT 104.150 32.920 104.450 33.220 ;
        RECT 104.640 32.920 104.940 33.220 ;
        RECT 106.530 32.920 106.830 33.220 ;
        RECT 107.020 32.920 107.320 33.220 ;
        RECT 107.510 32.920 107.810 33.220 ;
      LAYER met1 ;
        RECT 22.390 48.590 26.660 48.950 ;
        RECT 31.240 48.590 32.740 48.950 ;
        RECT 40.100 48.590 44.370 48.950 ;
        RECT 48.950 48.590 50.450 48.950 ;
        RECT 57.810 48.590 62.080 48.950 ;
        RECT 66.660 48.590 68.160 48.950 ;
        RECT 75.520 48.590 79.790 48.950 ;
        RECT 84.370 48.590 85.870 48.950 ;
        RECT 93.230 48.590 97.500 48.950 ;
        RECT 102.080 48.590 103.580 48.950 ;
        RECT 23.005 47.590 23.365 48.590 ;
        RECT 31.790 47.590 32.150 48.590 ;
        RECT 40.715 47.590 41.075 48.590 ;
        RECT 49.500 47.590 49.860 48.590 ;
        RECT 58.425 47.590 58.785 48.590 ;
        RECT 67.210 47.590 67.570 48.590 ;
        RECT 76.135 47.590 76.495 48.590 ;
        RECT 84.920 47.590 85.280 48.590 ;
        RECT 93.845 47.590 94.205 48.590 ;
        RECT 102.630 47.590 102.990 48.590 ;
        RECT 14.620 47.230 23.365 47.590 ;
        RECT 24.315 47.230 41.075 47.590 ;
        RECT 42.025 47.230 58.785 47.590 ;
        RECT 59.735 47.230 76.495 47.590 ;
        RECT 77.445 47.230 94.205 47.590 ;
        RECT 95.155 47.230 106.360 47.590 ;
        RECT 14.620 42.000 14.980 47.230 ;
        RECT 6.350 41.640 14.980 42.000 ;
        RECT 15.980 41.670 105.050 42.150 ;
        RECT 106.000 42.000 106.360 47.230 ;
        RECT 109.500 44.500 110.500 45.515 ;
        RECT 106.000 41.640 115.500 42.000 ;
        RECT 6.350 34.610 6.710 41.640 ;
        RECT 7.500 39.690 114.280 40.170 ;
        RECT 115.140 34.610 115.500 41.640 ;
        RECT 6.350 34.250 17.395 34.610 ;
        RECT 18.345 34.250 35.105 34.610 ;
        RECT 36.055 34.250 52.815 34.610 ;
        RECT 53.765 34.250 70.525 34.610 ;
        RECT 71.475 34.250 88.235 34.610 ;
        RECT 89.185 34.250 105.945 34.610 ;
        RECT 106.895 34.250 115.500 34.610 ;
        RECT 9.560 33.250 9.920 34.250 ;
        RECT 18.345 33.250 18.705 34.250 ;
        RECT 27.270 33.250 27.630 34.250 ;
        RECT 36.055 33.250 36.415 34.250 ;
        RECT 44.980 33.250 45.340 34.250 ;
        RECT 53.765 33.250 54.125 34.250 ;
        RECT 62.690 33.250 63.050 34.250 ;
        RECT 71.475 33.250 71.835 34.250 ;
        RECT 80.400 33.250 80.760 34.250 ;
        RECT 89.185 33.250 89.545 34.250 ;
        RECT 98.110 33.250 98.470 34.250 ;
        RECT 106.895 33.250 107.255 34.250 ;
        RECT 8.970 32.890 10.470 33.250 ;
        RECT 15.050 32.890 19.320 33.250 ;
        RECT 26.680 32.890 28.180 33.250 ;
        RECT 32.760 32.890 37.030 33.250 ;
        RECT 44.390 32.890 45.890 33.250 ;
        RECT 50.470 32.890 54.740 33.250 ;
        RECT 62.100 32.890 63.600 33.250 ;
        RECT 68.180 32.890 72.450 33.250 ;
        RECT 79.810 32.890 81.310 33.250 ;
        RECT 85.890 32.890 90.160 33.250 ;
        RECT 97.520 32.890 99.020 33.250 ;
        RECT 103.600 32.890 107.870 33.250 ;
      LAYER via ;
        RECT 19.500 41.770 19.760 42.030 ;
        RECT 19.870 41.770 20.130 42.030 ;
        RECT 20.240 41.770 20.500 42.030 ;
        RECT 25.500 41.770 25.760 42.030 ;
        RECT 25.870 41.770 26.130 42.030 ;
        RECT 26.240 41.770 26.500 42.030 ;
        RECT 31.500 41.770 31.760 42.030 ;
        RECT 31.870 41.770 32.130 42.030 ;
        RECT 32.240 41.770 32.500 42.030 ;
        RECT 37.500 41.770 37.760 42.030 ;
        RECT 37.870 41.770 38.130 42.030 ;
        RECT 38.240 41.770 38.500 42.030 ;
        RECT 43.500 41.770 43.760 42.030 ;
        RECT 43.870 41.770 44.130 42.030 ;
        RECT 44.240 41.770 44.500 42.030 ;
        RECT 49.500 41.770 49.760 42.030 ;
        RECT 49.870 41.770 50.130 42.030 ;
        RECT 50.240 41.770 50.500 42.030 ;
        RECT 55.500 41.770 55.760 42.030 ;
        RECT 55.870 41.770 56.130 42.030 ;
        RECT 56.240 41.770 56.500 42.030 ;
        RECT 61.500 41.770 61.760 42.030 ;
        RECT 61.870 41.770 62.130 42.030 ;
        RECT 62.240 41.770 62.500 42.030 ;
        RECT 67.500 41.770 67.760 42.030 ;
        RECT 67.870 41.770 68.130 42.030 ;
        RECT 68.240 41.770 68.500 42.030 ;
        RECT 73.500 41.770 73.760 42.030 ;
        RECT 73.870 41.770 74.130 42.030 ;
        RECT 74.240 41.770 74.500 42.030 ;
        RECT 79.500 41.770 79.760 42.030 ;
        RECT 79.870 41.770 80.130 42.030 ;
        RECT 80.240 41.770 80.500 42.030 ;
        RECT 85.500 41.770 85.760 42.030 ;
        RECT 85.870 41.770 86.130 42.030 ;
        RECT 86.240 41.770 86.500 42.030 ;
        RECT 91.500 41.770 91.760 42.030 ;
        RECT 91.870 41.770 92.130 42.030 ;
        RECT 92.240 41.770 92.500 42.030 ;
        RECT 97.500 41.770 97.760 42.030 ;
        RECT 97.870 41.770 98.130 42.030 ;
        RECT 98.240 41.770 98.500 42.030 ;
        RECT 103.500 41.770 103.760 42.030 ;
        RECT 103.870 41.770 104.130 42.030 ;
        RECT 104.240 41.770 104.500 42.030 ;
        RECT 109.570 45.100 109.910 45.440 ;
        RECT 110.090 45.100 110.430 45.440 ;
        RECT 109.570 44.580 109.910 44.920 ;
        RECT 110.090 44.580 110.430 44.920 ;
        RECT 7.500 39.790 7.760 40.050 ;
        RECT 7.870 39.790 8.130 40.050 ;
        RECT 8.240 39.790 8.500 40.050 ;
        RECT 13.500 39.790 13.760 40.050 ;
        RECT 13.870 39.790 14.130 40.050 ;
        RECT 14.240 39.790 14.500 40.050 ;
        RECT 19.500 39.790 19.760 40.050 ;
        RECT 19.870 39.790 20.130 40.050 ;
        RECT 20.240 39.790 20.500 40.050 ;
        RECT 25.500 39.790 25.760 40.050 ;
        RECT 25.870 39.790 26.130 40.050 ;
        RECT 26.240 39.790 26.500 40.050 ;
        RECT 31.500 39.790 31.760 40.050 ;
        RECT 31.870 39.790 32.130 40.050 ;
        RECT 32.240 39.790 32.500 40.050 ;
        RECT 37.500 39.790 37.760 40.050 ;
        RECT 37.870 39.790 38.130 40.050 ;
        RECT 38.240 39.790 38.500 40.050 ;
        RECT 43.500 39.790 43.760 40.050 ;
        RECT 43.870 39.790 44.130 40.050 ;
        RECT 44.240 39.790 44.500 40.050 ;
        RECT 49.500 39.790 49.760 40.050 ;
        RECT 49.870 39.790 50.130 40.050 ;
        RECT 50.240 39.790 50.500 40.050 ;
        RECT 55.500 39.790 55.760 40.050 ;
        RECT 55.870 39.790 56.130 40.050 ;
        RECT 56.240 39.790 56.500 40.050 ;
        RECT 61.500 39.790 61.760 40.050 ;
        RECT 61.870 39.790 62.130 40.050 ;
        RECT 62.240 39.790 62.500 40.050 ;
        RECT 67.500 39.790 67.760 40.050 ;
        RECT 67.870 39.790 68.130 40.050 ;
        RECT 68.240 39.790 68.500 40.050 ;
        RECT 73.500 39.790 73.760 40.050 ;
        RECT 73.870 39.790 74.130 40.050 ;
        RECT 74.240 39.790 74.500 40.050 ;
        RECT 79.500 39.790 79.760 40.050 ;
        RECT 79.870 39.790 80.130 40.050 ;
        RECT 80.240 39.790 80.500 40.050 ;
        RECT 85.500 39.790 85.760 40.050 ;
        RECT 85.870 39.790 86.130 40.050 ;
        RECT 86.240 39.790 86.500 40.050 ;
        RECT 91.500 39.790 91.760 40.050 ;
        RECT 91.870 39.790 92.130 40.050 ;
        RECT 92.240 39.790 92.500 40.050 ;
        RECT 97.500 39.790 97.760 40.050 ;
        RECT 97.870 39.790 98.130 40.050 ;
        RECT 98.240 39.790 98.500 40.050 ;
        RECT 103.500 39.790 103.760 40.050 ;
        RECT 103.870 39.790 104.130 40.050 ;
        RECT 104.240 39.790 104.500 40.050 ;
        RECT 109.500 39.790 109.760 40.050 ;
        RECT 109.870 39.790 110.130 40.050 ;
        RECT 110.240 39.790 110.500 40.050 ;
        RECT 113.280 39.790 113.540 40.050 ;
        RECT 113.650 39.790 113.910 40.050 ;
        RECT 114.020 39.790 114.280 40.050 ;
      LAYER met2 ;
        RECT 109.500 44.500 110.500 45.515 ;
        RECT 19.500 41.700 20.500 42.100 ;
        RECT 25.500 41.700 26.500 42.100 ;
        RECT 31.500 41.700 32.500 42.100 ;
        RECT 37.500 41.700 38.500 42.100 ;
        RECT 43.500 41.700 44.500 42.100 ;
        RECT 49.500 41.700 50.500 42.100 ;
        RECT 55.500 41.700 56.500 42.100 ;
        RECT 61.500 41.700 62.500 42.100 ;
        RECT 67.500 41.700 68.500 42.100 ;
        RECT 73.500 41.700 74.500 42.100 ;
        RECT 79.500 41.700 80.500 42.100 ;
        RECT 85.500 41.700 86.500 42.100 ;
        RECT 91.500 41.700 92.500 42.100 ;
        RECT 97.500 41.700 98.500 42.100 ;
        RECT 103.500 41.700 104.500 42.100 ;
        RECT 7.500 39.720 8.500 40.120 ;
        RECT 13.500 39.720 14.500 40.120 ;
        RECT 19.500 39.720 20.500 40.120 ;
        RECT 25.500 39.720 26.500 40.120 ;
        RECT 31.500 39.720 32.500 40.120 ;
        RECT 37.500 39.720 38.500 40.120 ;
        RECT 43.500 39.720 44.500 40.120 ;
        RECT 49.500 39.720 50.500 40.120 ;
        RECT 55.500 39.720 56.500 40.120 ;
        RECT 61.500 39.720 62.500 40.120 ;
        RECT 67.500 39.720 68.500 40.120 ;
        RECT 73.500 39.720 74.500 40.120 ;
        RECT 79.500 39.720 80.500 40.120 ;
        RECT 85.500 39.720 86.500 40.120 ;
        RECT 91.500 39.720 92.500 40.120 ;
        RECT 97.500 39.720 98.500 40.120 ;
        RECT 103.500 39.720 104.500 40.120 ;
        RECT 109.500 39.720 110.500 40.120 ;
        RECT 113.280 39.720 114.280 40.120 ;
      LAYER via2 ;
        RECT 109.540 45.070 109.940 45.470 ;
        RECT 110.060 45.070 110.460 45.470 ;
        RECT 109.540 44.550 109.940 44.950 ;
        RECT 110.060 44.550 110.460 44.950 ;
        RECT 19.600 41.750 19.900 42.050 ;
        RECT 20.100 41.750 20.400 42.050 ;
        RECT 25.600 41.750 25.900 42.050 ;
        RECT 26.100 41.750 26.400 42.050 ;
        RECT 31.600 41.750 31.900 42.050 ;
        RECT 32.100 41.750 32.400 42.050 ;
        RECT 37.600 41.750 37.900 42.050 ;
        RECT 38.100 41.750 38.400 42.050 ;
        RECT 43.600 41.750 43.900 42.050 ;
        RECT 44.100 41.750 44.400 42.050 ;
        RECT 49.600 41.750 49.900 42.050 ;
        RECT 50.100 41.750 50.400 42.050 ;
        RECT 55.600 41.750 55.900 42.050 ;
        RECT 56.100 41.750 56.400 42.050 ;
        RECT 61.600 41.750 61.900 42.050 ;
        RECT 62.100 41.750 62.400 42.050 ;
        RECT 67.600 41.750 67.900 42.050 ;
        RECT 68.100 41.750 68.400 42.050 ;
        RECT 73.600 41.750 73.900 42.050 ;
        RECT 74.100 41.750 74.400 42.050 ;
        RECT 79.600 41.750 79.900 42.050 ;
        RECT 80.100 41.750 80.400 42.050 ;
        RECT 85.600 41.750 85.900 42.050 ;
        RECT 86.100 41.750 86.400 42.050 ;
        RECT 91.600 41.750 91.900 42.050 ;
        RECT 92.100 41.750 92.400 42.050 ;
        RECT 97.600 41.750 97.900 42.050 ;
        RECT 98.100 41.750 98.400 42.050 ;
        RECT 103.600 41.750 103.900 42.050 ;
        RECT 104.100 41.750 104.400 42.050 ;
        RECT 7.600 39.770 7.900 40.070 ;
        RECT 8.100 39.770 8.400 40.070 ;
        RECT 13.600 39.770 13.900 40.070 ;
        RECT 14.100 39.770 14.400 40.070 ;
        RECT 19.600 39.770 19.900 40.070 ;
        RECT 20.100 39.770 20.400 40.070 ;
        RECT 25.600 39.770 25.900 40.070 ;
        RECT 26.100 39.770 26.400 40.070 ;
        RECT 31.600 39.770 31.900 40.070 ;
        RECT 32.100 39.770 32.400 40.070 ;
        RECT 37.600 39.770 37.900 40.070 ;
        RECT 38.100 39.770 38.400 40.070 ;
        RECT 43.600 39.770 43.900 40.070 ;
        RECT 44.100 39.770 44.400 40.070 ;
        RECT 49.600 39.770 49.900 40.070 ;
        RECT 50.100 39.770 50.400 40.070 ;
        RECT 55.600 39.770 55.900 40.070 ;
        RECT 56.100 39.770 56.400 40.070 ;
        RECT 61.600 39.770 61.900 40.070 ;
        RECT 62.100 39.770 62.400 40.070 ;
        RECT 67.600 39.770 67.900 40.070 ;
        RECT 68.100 39.770 68.400 40.070 ;
        RECT 73.600 39.770 73.900 40.070 ;
        RECT 74.100 39.770 74.400 40.070 ;
        RECT 79.600 39.770 79.900 40.070 ;
        RECT 80.100 39.770 80.400 40.070 ;
        RECT 85.600 39.770 85.900 40.070 ;
        RECT 86.100 39.770 86.400 40.070 ;
        RECT 91.600 39.770 91.900 40.070 ;
        RECT 92.100 39.770 92.400 40.070 ;
        RECT 97.600 39.770 97.900 40.070 ;
        RECT 98.100 39.770 98.400 40.070 ;
        RECT 103.600 39.770 103.900 40.070 ;
        RECT 104.100 39.770 104.400 40.070 ;
        RECT 109.600 39.770 109.900 40.070 ;
        RECT 110.100 39.770 110.400 40.070 ;
        RECT 113.380 39.770 113.680 40.070 ;
        RECT 113.880 39.770 114.180 40.070 ;
      LAYER met3 ;
        RECT 19.500 41.670 20.500 42.150 ;
        RECT 25.500 41.670 26.500 42.150 ;
        RECT 31.500 41.670 32.500 42.150 ;
        RECT 37.500 41.670 38.500 42.150 ;
        RECT 43.500 41.670 44.500 42.150 ;
        RECT 49.500 41.670 50.500 42.150 ;
        RECT 55.500 41.670 56.500 42.150 ;
        RECT 61.500 41.670 62.500 42.150 ;
        RECT 67.500 41.670 68.500 42.150 ;
        RECT 73.500 41.670 74.500 42.150 ;
        RECT 79.500 41.670 80.500 42.150 ;
        RECT 85.500 41.670 86.500 42.150 ;
        RECT 91.500 41.670 92.500 42.150 ;
        RECT 97.500 41.670 98.500 42.150 ;
        RECT 103.500 41.670 104.500 42.150 ;
        RECT 109.500 41.670 110.500 45.515 ;
        RECT 7.500 40.170 114.280 41.670 ;
        RECT 7.500 39.690 8.500 40.170 ;
        RECT 13.500 39.690 14.500 40.170 ;
        RECT 19.500 39.690 20.500 40.170 ;
        RECT 25.500 39.690 26.500 40.170 ;
        RECT 31.500 39.690 32.500 40.170 ;
        RECT 37.500 39.690 38.500 40.170 ;
        RECT 43.500 39.690 44.500 40.170 ;
        RECT 49.500 39.690 50.500 40.170 ;
        RECT 55.500 39.690 56.500 40.170 ;
        RECT 61.500 39.690 62.500 40.170 ;
        RECT 67.500 39.690 68.500 40.170 ;
        RECT 73.500 39.690 74.500 40.170 ;
        RECT 79.500 39.690 80.500 40.170 ;
        RECT 85.500 39.690 86.500 40.170 ;
        RECT 91.500 39.690 92.500 40.170 ;
        RECT 97.500 39.690 98.500 40.170 ;
        RECT 103.500 39.690 104.500 40.170 ;
        RECT 109.500 39.690 110.500 40.170 ;
        RECT 113.280 39.690 114.280 40.170 ;
  END
END vco_w6_r100
END LIBRARY

