VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ring_osc_r100
  CLASS BLOCK ;
  FOREIGN ring_osc_r100 ;
  ORIGIN 0.000 1.290 ;
  SIZE 181.500 BY 40.660 ;
  OBS
      LAYER pwell ;
        RECT 18.390 32.310 28.420 38.370 ;
      LAYER nwell ;
        RECT 3.630 28.505 6.310 30.340 ;
        RECT 7.800 28.505 9.560 30.340 ;
      LAYER pwell ;
        RECT 4.310 27.985 6.115 28.215 ;
        RECT 3.825 27.305 6.115 27.985 ;
        RECT 3.970 27.115 4.140 27.305 ;
        RECT 8.135 27.115 8.305 27.285 ;
      LAYER nwell ;
        RECT 18.390 24.245 24.240 30.120 ;
        RECT 29.220 29.780 35.070 35.635 ;
      LAYER pwell ;
        RECT 36.365 32.270 42.215 38.370 ;
      LAYER nwell ;
        RECT 42.840 30.310 46.600 35.585 ;
      LAYER pwell ;
        RECT 47.890 32.310 57.920 38.370 ;
        RECT 25.040 21.460 35.070 27.860 ;
      LAYER nwell ;
        RECT 36.365 24.250 40.125 29.560 ;
      LAYER pwell ;
        RECT 40.745 26.625 46.595 27.565 ;
        RECT 40.745 26.575 46.600 26.625 ;
        RECT 40.750 21.465 46.600 26.575 ;
      LAYER nwell ;
        RECT 47.890 24.245 53.740 30.120 ;
        RECT 58.720 29.780 64.570 35.635 ;
      LAYER pwell ;
        RECT 65.865 32.270 71.715 38.370 ;
      LAYER nwell ;
        RECT 72.340 30.310 76.100 35.585 ;
      LAYER pwell ;
        RECT 77.390 32.310 87.420 38.370 ;
        RECT 54.540 21.460 64.570 27.860 ;
      LAYER nwell ;
        RECT 65.865 24.250 69.625 29.560 ;
      LAYER pwell ;
        RECT 70.245 26.625 76.095 27.565 ;
        RECT 70.245 26.575 76.100 26.625 ;
        RECT 70.250 21.465 76.100 26.575 ;
      LAYER nwell ;
        RECT 77.390 24.245 83.240 30.120 ;
        RECT 88.220 29.780 94.070 35.635 ;
      LAYER pwell ;
        RECT 95.365 32.270 101.215 38.370 ;
      LAYER nwell ;
        RECT 101.840 30.310 105.600 35.585 ;
      LAYER pwell ;
        RECT 106.890 32.310 116.920 38.370 ;
        RECT 84.040 21.460 94.070 27.860 ;
      LAYER nwell ;
        RECT 95.365 24.250 99.125 29.560 ;
      LAYER pwell ;
        RECT 99.745 26.625 105.595 27.565 ;
        RECT 99.745 26.575 105.600 26.625 ;
        RECT 99.750 21.465 105.600 26.575 ;
      LAYER nwell ;
        RECT 106.890 24.245 112.740 30.120 ;
        RECT 117.720 29.780 123.570 35.635 ;
      LAYER pwell ;
        RECT 124.865 32.270 130.715 38.370 ;
      LAYER nwell ;
        RECT 131.340 30.310 135.100 35.585 ;
      LAYER pwell ;
        RECT 136.390 32.310 146.420 38.370 ;
        RECT 113.540 21.460 123.570 27.860 ;
      LAYER nwell ;
        RECT 124.865 24.250 128.625 29.560 ;
      LAYER pwell ;
        RECT 129.245 26.625 135.095 27.565 ;
        RECT 129.245 26.575 135.100 26.625 ;
        RECT 129.250 21.465 135.100 26.575 ;
      LAYER nwell ;
        RECT 136.390 24.245 142.240 30.120 ;
        RECT 147.220 29.780 153.070 35.635 ;
      LAYER pwell ;
        RECT 154.365 32.270 160.215 38.370 ;
      LAYER nwell ;
        RECT 160.840 30.310 164.600 35.585 ;
      LAYER pwell ;
        RECT 143.040 21.460 153.070 27.860 ;
      LAYER nwell ;
        RECT 154.365 24.250 158.125 29.560 ;
      LAYER pwell ;
        RECT 158.745 26.625 164.595 27.565 ;
        RECT 158.745 26.575 164.600 26.625 ;
        RECT 158.750 21.465 164.600 26.575 ;
        RECT 171.590 20.280 178.380 27.280 ;
        RECT 2.790 11.505 8.640 16.615 ;
        RECT 2.790 11.455 8.645 11.505 ;
        RECT 2.795 10.515 8.645 11.455 ;
      LAYER nwell ;
        RECT 9.265 8.520 13.025 13.830 ;
      LAYER pwell ;
        RECT 14.320 10.220 24.350 16.620 ;
      LAYER nwell ;
        RECT 2.790 2.495 6.550 7.770 ;
      LAYER pwell ;
        RECT 7.175 -0.290 13.025 5.810 ;
      LAYER nwell ;
        RECT 14.320 2.445 20.170 8.300 ;
        RECT 25.150 7.960 31.000 13.835 ;
      LAYER pwell ;
        RECT 32.290 11.505 38.140 16.615 ;
        RECT 32.290 11.455 38.145 11.505 ;
        RECT 32.295 10.515 38.145 11.455 ;
      LAYER nwell ;
        RECT 38.765 8.520 42.525 13.830 ;
      LAYER pwell ;
        RECT 43.820 10.220 53.850 16.620 ;
        RECT 20.970 -0.290 31.000 5.770 ;
      LAYER nwell ;
        RECT 32.290 2.495 36.050 7.770 ;
      LAYER pwell ;
        RECT 36.675 -0.290 42.525 5.810 ;
      LAYER nwell ;
        RECT 43.820 2.445 49.670 8.300 ;
        RECT 54.650 7.960 60.500 13.835 ;
      LAYER pwell ;
        RECT 61.790 11.505 67.640 16.615 ;
        RECT 61.790 11.455 67.645 11.505 ;
        RECT 61.795 10.515 67.645 11.455 ;
      LAYER nwell ;
        RECT 68.265 8.520 72.025 13.830 ;
      LAYER pwell ;
        RECT 73.320 10.220 83.350 16.620 ;
        RECT 50.470 -0.290 60.500 5.770 ;
      LAYER nwell ;
        RECT 61.790 2.495 65.550 7.770 ;
      LAYER pwell ;
        RECT 66.175 -0.290 72.025 5.810 ;
      LAYER nwell ;
        RECT 73.320 2.445 79.170 8.300 ;
        RECT 84.150 7.960 90.000 13.835 ;
      LAYER pwell ;
        RECT 91.290 11.505 97.140 16.615 ;
        RECT 91.290 11.455 97.145 11.505 ;
        RECT 91.295 10.515 97.145 11.455 ;
      LAYER nwell ;
        RECT 97.765 8.520 101.525 13.830 ;
      LAYER pwell ;
        RECT 102.820 10.220 112.850 16.620 ;
        RECT 79.970 -0.290 90.000 5.770 ;
      LAYER nwell ;
        RECT 91.290 2.495 95.050 7.770 ;
      LAYER pwell ;
        RECT 95.675 -0.290 101.525 5.810 ;
      LAYER nwell ;
        RECT 102.820 2.445 108.670 8.300 ;
        RECT 113.650 7.960 119.500 13.835 ;
      LAYER pwell ;
        RECT 120.790 11.505 126.640 16.615 ;
        RECT 120.790 11.455 126.645 11.505 ;
        RECT 120.795 10.515 126.645 11.455 ;
      LAYER nwell ;
        RECT 127.265 8.520 131.025 13.830 ;
      LAYER pwell ;
        RECT 132.320 10.220 142.350 16.620 ;
        RECT 109.470 -0.290 119.500 5.770 ;
      LAYER nwell ;
        RECT 120.790 2.495 124.550 7.770 ;
      LAYER pwell ;
        RECT 125.175 -0.290 131.025 5.810 ;
      LAYER nwell ;
        RECT 132.320 2.445 138.170 8.300 ;
        RECT 143.150 7.960 149.000 13.835 ;
      LAYER pwell ;
        RECT 150.290 11.505 156.140 16.615 ;
        RECT 150.290 11.455 156.145 11.505 ;
        RECT 150.295 10.515 156.145 11.455 ;
      LAYER nwell ;
        RECT 156.765 8.520 160.525 13.830 ;
      LAYER pwell ;
        RECT 161.820 10.220 171.850 16.620 ;
        RECT 138.970 -0.290 149.000 5.770 ;
      LAYER nwell ;
        RECT 150.290 2.495 154.050 7.770 ;
      LAYER pwell ;
        RECT 154.675 -0.290 160.525 5.810 ;
      LAYER nwell ;
        RECT 161.820 2.445 167.670 8.300 ;
        RECT 172.650 7.960 178.500 13.835 ;
      LAYER pwell ;
        RECT 168.470 -0.290 178.500 5.770 ;
      LAYER li1 ;
        RECT 18.570 37.840 20.915 38.320 ;
        RECT 21.980 37.840 24.840 38.320 ;
        RECT 25.895 37.840 28.240 38.320 ;
        RECT 36.545 37.840 38.890 38.320 ;
        RECT 39.690 37.840 42.035 38.320 ;
        RECT 48.070 37.840 50.415 38.320 ;
        RECT 51.480 37.840 54.340 38.320 ;
        RECT 55.395 37.840 57.740 38.320 ;
        RECT 66.045 37.840 68.390 38.320 ;
        RECT 69.190 37.840 71.535 38.320 ;
        RECT 77.570 37.840 79.915 38.320 ;
        RECT 80.980 37.840 83.840 38.320 ;
        RECT 84.895 37.840 87.240 38.320 ;
        RECT 95.545 37.840 97.890 38.320 ;
        RECT 98.690 37.840 101.035 38.320 ;
        RECT 107.070 37.840 109.415 38.320 ;
        RECT 110.480 37.840 113.340 38.320 ;
        RECT 114.395 37.840 116.740 38.320 ;
        RECT 125.045 37.840 127.390 38.320 ;
        RECT 128.190 37.840 130.535 38.320 ;
        RECT 136.570 37.840 138.915 38.320 ;
        RECT 139.980 37.840 142.840 38.320 ;
        RECT 143.895 37.840 146.240 38.320 ;
        RECT 154.545 37.840 156.890 38.320 ;
        RECT 157.690 37.840 160.035 38.320 ;
        RECT 19.080 33.245 19.370 37.840 ;
        RECT 19.140 33.000 19.310 33.245 ;
        RECT 19.290 30.790 20.420 31.790 ;
        RECT 21.170 31.480 21.460 37.540 ;
        RECT 23.260 33.245 23.550 37.840 ;
        RECT 23.320 33.000 23.490 33.245 ;
        RECT 25.350 31.580 25.640 37.540 ;
        RECT 27.440 33.245 27.730 37.840 ;
        RECT 29.400 35.455 31.745 35.600 ;
        RECT 32.545 35.455 34.890 35.600 ;
        RECT 29.400 35.285 34.890 35.455 ;
        RECT 29.400 35.120 31.745 35.285 ;
        RECT 32.545 35.120 34.890 35.285 ;
        RECT 27.500 33.235 27.695 33.245 ;
        RECT 27.500 33.000 27.670 33.235 ;
        RECT 25.350 31.480 26.170 31.580 ;
        RECT 21.170 30.980 26.170 31.480 ;
        RECT 4.340 30.005 5.310 30.160 ;
        RECT 8.340 30.005 9.310 30.160 ;
        RECT 3.820 29.835 6.120 30.005 ;
        RECT 7.990 29.835 9.370 30.005 ;
        RECT 3.905 29.265 4.165 29.665 ;
        RECT 4.335 29.435 5.270 29.835 ;
        RECT 5.440 29.325 6.035 29.665 ;
        RECT 3.905 29.095 5.270 29.265 ;
        RECT 3.905 28.195 4.365 28.925 ;
        RECT 4.535 28.025 5.270 29.095 ;
        RECT 3.905 27.855 5.270 28.025 ;
        RECT 5.440 28.005 5.615 29.325 ;
        RECT 6.330 29.155 7.780 29.375 ;
        RECT 5.795 29.075 7.780 29.155 ;
        RECT 8.265 29.110 8.595 29.835 ;
        RECT 5.795 28.855 6.630 29.075 ;
        RECT 7.480 28.940 7.780 29.075 ;
        RECT 5.795 28.175 6.035 28.855 ;
        RECT 5.440 27.875 6.035 28.005 ;
        RECT 6.860 27.875 7.160 28.710 ;
        RECT 7.480 28.640 8.595 28.940 ;
        RECT 3.905 27.455 4.165 27.855 ;
        RECT 4.335 27.285 5.270 27.685 ;
        RECT 5.440 27.575 7.160 27.875 ;
        RECT 5.440 27.455 6.035 27.575 ;
        RECT 8.075 27.455 8.595 28.640 ;
        RECT 8.765 28.115 9.285 29.665 ;
        RECT 8.765 27.285 9.105 27.945 ;
        RECT 3.820 27.115 6.120 27.285 ;
        RECT 7.990 27.115 9.370 27.285 ;
        RECT 18.570 24.720 18.740 29.575 ;
        RECT 19.080 24.720 19.370 29.570 ;
        RECT 21.170 25.030 21.460 30.980 ;
        RECT 29.400 30.460 29.570 35.120 ;
        RECT 29.910 30.290 30.200 35.120 ;
        RECT 32.000 29.850 32.290 34.850 ;
        RECT 34.090 30.290 34.380 35.120 ;
        RECT 34.720 30.520 34.890 35.120 ;
        RECT 37.055 33.490 37.345 37.840 ;
        RECT 37.290 31.580 38.490 31.890 ;
        RECT 36.790 30.960 38.490 31.580 ;
        RECT 37.290 30.760 38.490 30.960 ;
        RECT 39.140 29.850 39.435 37.530 ;
        RECT 41.235 33.490 41.525 37.840 ;
        RECT 44.325 35.570 46.420 35.600 ;
        RECT 44.170 35.405 46.420 35.570 ;
        RECT 43.020 35.235 46.420 35.405 ;
        RECT 43.020 32.260 43.190 35.235 ;
        RECT 44.170 35.150 46.420 35.235 ;
        RECT 44.325 35.120 46.420 35.150 ;
        RECT 43.525 31.675 43.820 34.750 ;
        RECT 43.295 30.895 44.035 31.675 ;
        RECT 23.260 24.720 23.550 29.570 ;
        RECT 23.890 24.720 24.060 29.575 ;
        RECT 29.360 29.350 41.955 29.850 ;
        RECT 29.360 27.910 29.860 29.350 ;
        RECT 30.890 28.320 34.890 28.920 ;
        RECT 32.890 28.200 34.890 28.320 ;
        RECT 27.820 27.620 32.290 27.910 ;
        RECT 32.890 27.620 34.090 28.200 ;
        RECT 25.790 26.595 25.960 26.830 ;
        RECT 25.765 26.585 25.960 26.595 ;
        RECT 18.570 24.595 20.915 24.720 ;
        RECT 21.715 24.690 24.060 24.720 ;
        RECT 21.715 24.595 24.240 24.690 ;
        RECT 18.570 24.425 24.240 24.595 ;
        RECT 18.570 24.240 20.915 24.425 ;
        RECT 21.715 24.270 24.240 24.425 ;
        RECT 21.715 24.240 24.060 24.270 ;
        RECT 25.730 22.000 26.020 26.585 ;
        RECT 27.820 22.290 28.110 27.620 ;
        RECT 29.970 26.585 30.140 26.810 ;
        RECT 29.910 22.000 30.200 26.585 ;
        RECT 32.000 22.290 32.290 27.620 ;
        RECT 34.150 26.585 34.320 26.810 ;
        RECT 34.090 22.000 34.380 26.585 ;
        RECT 36.545 24.720 36.715 28.645 ;
        RECT 37.055 24.720 37.345 28.790 ;
        RECT 39.145 25.085 39.440 29.350 ;
        RECT 36.545 24.690 38.640 24.720 ;
        RECT 36.545 24.600 38.795 24.690 ;
        RECT 39.775 24.600 39.945 28.635 ;
        RECT 41.455 28.200 41.955 29.350 ;
        RECT 36.545 24.430 39.945 24.600 ;
        RECT 36.545 24.270 38.795 24.430 ;
        RECT 36.545 24.240 38.640 24.270 ;
        RECT 41.440 22.000 41.730 26.345 ;
        RECT 43.525 22.305 43.820 30.895 ;
        RECT 45.620 30.710 45.910 35.120 ;
        RECT 46.250 30.705 46.420 35.120 ;
        RECT 48.580 33.245 48.870 37.840 ;
        RECT 48.640 33.000 48.810 33.245 ;
        RECT 48.790 30.790 49.920 31.790 ;
        RECT 50.670 31.480 50.960 37.540 ;
        RECT 52.760 33.245 53.050 37.840 ;
        RECT 52.820 33.000 52.990 33.245 ;
        RECT 54.850 31.580 55.140 37.540 ;
        RECT 56.940 33.245 57.230 37.840 ;
        RECT 58.900 35.455 61.245 35.600 ;
        RECT 62.045 35.455 64.390 35.600 ;
        RECT 58.900 35.285 64.390 35.455 ;
        RECT 58.900 35.120 61.245 35.285 ;
        RECT 62.045 35.120 64.390 35.285 ;
        RECT 57.000 33.235 57.195 33.245 ;
        RECT 57.000 33.000 57.170 33.235 ;
        RECT 54.850 31.480 55.670 31.580 ;
        RECT 50.670 30.980 55.670 31.480 ;
        RECT 44.440 28.860 45.620 29.060 ;
        RECT 44.440 28.260 46.120 28.860 ;
        RECT 44.440 27.980 45.620 28.260 ;
        RECT 45.620 22.000 45.910 26.345 ;
        RECT 48.070 24.720 48.240 29.575 ;
        RECT 48.580 24.720 48.870 29.570 ;
        RECT 50.670 25.030 50.960 30.980 ;
        RECT 58.900 30.460 59.070 35.120 ;
        RECT 59.410 30.290 59.700 35.120 ;
        RECT 61.500 29.850 61.790 34.850 ;
        RECT 63.590 30.290 63.880 35.120 ;
        RECT 64.220 30.520 64.390 35.120 ;
        RECT 66.555 33.490 66.845 37.840 ;
        RECT 66.790 31.580 67.990 31.890 ;
        RECT 66.290 30.960 67.990 31.580 ;
        RECT 66.790 30.760 67.990 30.960 ;
        RECT 68.640 29.850 68.935 37.530 ;
        RECT 70.735 33.490 71.025 37.840 ;
        RECT 73.825 35.570 75.920 35.600 ;
        RECT 73.670 35.405 75.920 35.570 ;
        RECT 72.520 35.235 75.920 35.405 ;
        RECT 72.520 32.260 72.690 35.235 ;
        RECT 73.670 35.150 75.920 35.235 ;
        RECT 73.825 35.120 75.920 35.150 ;
        RECT 73.025 31.675 73.320 34.750 ;
        RECT 72.795 30.895 73.535 31.675 ;
        RECT 52.760 24.720 53.050 29.570 ;
        RECT 53.390 24.720 53.560 29.575 ;
        RECT 58.860 29.350 71.455 29.850 ;
        RECT 58.860 27.910 59.360 29.350 ;
        RECT 60.390 28.320 64.390 28.920 ;
        RECT 62.390 28.200 64.390 28.320 ;
        RECT 57.320 27.620 61.790 27.910 ;
        RECT 62.390 27.620 63.590 28.200 ;
        RECT 55.290 26.595 55.460 26.830 ;
        RECT 55.265 26.585 55.460 26.595 ;
        RECT 48.070 24.595 50.415 24.720 ;
        RECT 51.215 24.690 53.560 24.720 ;
        RECT 51.215 24.595 53.740 24.690 ;
        RECT 48.070 24.425 53.740 24.595 ;
        RECT 48.070 24.240 50.415 24.425 ;
        RECT 51.215 24.270 53.740 24.425 ;
        RECT 51.215 24.240 53.560 24.270 ;
        RECT 55.230 22.000 55.520 26.585 ;
        RECT 57.320 22.290 57.610 27.620 ;
        RECT 59.470 26.585 59.640 26.810 ;
        RECT 59.410 22.000 59.700 26.585 ;
        RECT 61.500 22.290 61.790 27.620 ;
        RECT 63.650 26.585 63.820 26.810 ;
        RECT 63.590 22.000 63.880 26.585 ;
        RECT 66.045 24.720 66.215 28.645 ;
        RECT 66.555 24.720 66.845 28.790 ;
        RECT 68.645 25.085 68.940 29.350 ;
        RECT 66.045 24.690 68.140 24.720 ;
        RECT 66.045 24.600 68.295 24.690 ;
        RECT 69.275 24.600 69.445 28.635 ;
        RECT 70.955 28.200 71.455 29.350 ;
        RECT 66.045 24.430 69.445 24.600 ;
        RECT 66.045 24.270 68.295 24.430 ;
        RECT 66.045 24.240 68.140 24.270 ;
        RECT 70.940 22.000 71.230 26.345 ;
        RECT 73.025 22.305 73.320 30.895 ;
        RECT 75.120 30.710 75.410 35.120 ;
        RECT 75.750 30.705 75.920 35.120 ;
        RECT 78.080 33.245 78.370 37.840 ;
        RECT 78.140 33.000 78.310 33.245 ;
        RECT 78.290 30.790 79.420 31.790 ;
        RECT 80.170 31.480 80.460 37.540 ;
        RECT 82.260 33.245 82.550 37.840 ;
        RECT 82.320 33.000 82.490 33.245 ;
        RECT 84.350 31.580 84.640 37.540 ;
        RECT 86.440 33.245 86.730 37.840 ;
        RECT 88.400 35.455 90.745 35.600 ;
        RECT 91.545 35.455 93.890 35.600 ;
        RECT 88.400 35.285 93.890 35.455 ;
        RECT 88.400 35.120 90.745 35.285 ;
        RECT 91.545 35.120 93.890 35.285 ;
        RECT 86.500 33.235 86.695 33.245 ;
        RECT 86.500 33.000 86.670 33.235 ;
        RECT 84.350 31.480 85.170 31.580 ;
        RECT 80.170 30.980 85.170 31.480 ;
        RECT 73.940 28.860 75.120 29.060 ;
        RECT 73.940 28.260 75.620 28.860 ;
        RECT 73.940 27.980 75.120 28.260 ;
        RECT 75.120 22.000 75.410 26.345 ;
        RECT 77.570 24.720 77.740 29.575 ;
        RECT 78.080 24.720 78.370 29.570 ;
        RECT 80.170 25.030 80.460 30.980 ;
        RECT 88.400 30.460 88.570 35.120 ;
        RECT 88.910 30.290 89.200 35.120 ;
        RECT 91.000 29.850 91.290 34.850 ;
        RECT 93.090 30.290 93.380 35.120 ;
        RECT 93.720 30.520 93.890 35.120 ;
        RECT 96.055 33.490 96.345 37.840 ;
        RECT 96.290 31.580 97.490 31.890 ;
        RECT 95.790 30.960 97.490 31.580 ;
        RECT 96.290 30.760 97.490 30.960 ;
        RECT 98.140 29.850 98.435 37.530 ;
        RECT 100.235 33.490 100.525 37.840 ;
        RECT 103.325 35.570 105.420 35.600 ;
        RECT 103.170 35.405 105.420 35.570 ;
        RECT 102.020 35.235 105.420 35.405 ;
        RECT 102.020 32.260 102.190 35.235 ;
        RECT 103.170 35.150 105.420 35.235 ;
        RECT 103.325 35.120 105.420 35.150 ;
        RECT 102.525 31.675 102.820 34.750 ;
        RECT 102.295 30.895 103.035 31.675 ;
        RECT 82.260 24.720 82.550 29.570 ;
        RECT 82.890 24.720 83.060 29.575 ;
        RECT 88.360 29.350 100.955 29.850 ;
        RECT 88.360 27.910 88.860 29.350 ;
        RECT 89.890 28.320 93.890 28.920 ;
        RECT 91.890 28.200 93.890 28.320 ;
        RECT 86.820 27.620 91.290 27.910 ;
        RECT 91.890 27.620 93.090 28.200 ;
        RECT 84.790 26.595 84.960 26.830 ;
        RECT 84.765 26.585 84.960 26.595 ;
        RECT 77.570 24.595 79.915 24.720 ;
        RECT 80.715 24.690 83.060 24.720 ;
        RECT 80.715 24.595 83.240 24.690 ;
        RECT 77.570 24.425 83.240 24.595 ;
        RECT 77.570 24.240 79.915 24.425 ;
        RECT 80.715 24.270 83.240 24.425 ;
        RECT 80.715 24.240 83.060 24.270 ;
        RECT 84.730 22.000 85.020 26.585 ;
        RECT 86.820 22.290 87.110 27.620 ;
        RECT 88.970 26.585 89.140 26.810 ;
        RECT 88.910 22.000 89.200 26.585 ;
        RECT 91.000 22.290 91.290 27.620 ;
        RECT 93.150 26.585 93.320 26.810 ;
        RECT 93.090 22.000 93.380 26.585 ;
        RECT 95.545 24.720 95.715 28.645 ;
        RECT 96.055 24.720 96.345 28.790 ;
        RECT 98.145 25.085 98.440 29.350 ;
        RECT 95.545 24.690 97.640 24.720 ;
        RECT 95.545 24.600 97.795 24.690 ;
        RECT 98.775 24.600 98.945 28.635 ;
        RECT 100.455 28.200 100.955 29.350 ;
        RECT 95.545 24.430 98.945 24.600 ;
        RECT 95.545 24.270 97.795 24.430 ;
        RECT 95.545 24.240 97.640 24.270 ;
        RECT 100.440 22.000 100.730 26.345 ;
        RECT 102.525 22.305 102.820 30.895 ;
        RECT 104.620 30.710 104.910 35.120 ;
        RECT 105.250 30.705 105.420 35.120 ;
        RECT 107.580 33.245 107.870 37.840 ;
        RECT 107.640 33.000 107.810 33.245 ;
        RECT 107.790 30.790 108.920 31.790 ;
        RECT 109.670 31.480 109.960 37.540 ;
        RECT 111.760 33.245 112.050 37.840 ;
        RECT 111.820 33.000 111.990 33.245 ;
        RECT 113.850 31.580 114.140 37.540 ;
        RECT 115.940 33.245 116.230 37.840 ;
        RECT 117.900 35.455 120.245 35.600 ;
        RECT 121.045 35.455 123.390 35.600 ;
        RECT 117.900 35.285 123.390 35.455 ;
        RECT 117.900 35.120 120.245 35.285 ;
        RECT 121.045 35.120 123.390 35.285 ;
        RECT 116.000 33.235 116.195 33.245 ;
        RECT 116.000 33.000 116.170 33.235 ;
        RECT 113.850 31.480 114.670 31.580 ;
        RECT 109.670 30.980 114.670 31.480 ;
        RECT 103.440 28.860 104.620 29.060 ;
        RECT 103.440 28.260 105.120 28.860 ;
        RECT 103.440 27.980 104.620 28.260 ;
        RECT 104.620 22.000 104.910 26.345 ;
        RECT 107.070 24.720 107.240 29.575 ;
        RECT 107.580 24.720 107.870 29.570 ;
        RECT 109.670 25.030 109.960 30.980 ;
        RECT 117.900 30.460 118.070 35.120 ;
        RECT 118.410 30.290 118.700 35.120 ;
        RECT 120.500 29.850 120.790 34.850 ;
        RECT 122.590 30.290 122.880 35.120 ;
        RECT 123.220 30.520 123.390 35.120 ;
        RECT 125.555 33.490 125.845 37.840 ;
        RECT 125.790 31.580 126.990 31.890 ;
        RECT 125.290 30.960 126.990 31.580 ;
        RECT 125.790 30.760 126.990 30.960 ;
        RECT 127.640 29.850 127.935 37.530 ;
        RECT 129.735 33.490 130.025 37.840 ;
        RECT 132.825 35.570 134.920 35.600 ;
        RECT 132.670 35.405 134.920 35.570 ;
        RECT 131.520 35.235 134.920 35.405 ;
        RECT 131.520 32.260 131.690 35.235 ;
        RECT 132.670 35.150 134.920 35.235 ;
        RECT 132.825 35.120 134.920 35.150 ;
        RECT 132.025 31.675 132.320 34.750 ;
        RECT 131.795 30.895 132.535 31.675 ;
        RECT 111.760 24.720 112.050 29.570 ;
        RECT 112.390 24.720 112.560 29.575 ;
        RECT 117.860 29.350 130.455 29.850 ;
        RECT 117.860 27.910 118.360 29.350 ;
        RECT 119.390 28.320 123.390 28.920 ;
        RECT 121.390 28.200 123.390 28.320 ;
        RECT 116.320 27.620 120.790 27.910 ;
        RECT 121.390 27.620 122.590 28.200 ;
        RECT 114.290 26.595 114.460 26.830 ;
        RECT 114.265 26.585 114.460 26.595 ;
        RECT 107.070 24.595 109.415 24.720 ;
        RECT 110.215 24.690 112.560 24.720 ;
        RECT 110.215 24.595 112.740 24.690 ;
        RECT 107.070 24.425 112.740 24.595 ;
        RECT 107.070 24.240 109.415 24.425 ;
        RECT 110.215 24.270 112.740 24.425 ;
        RECT 110.215 24.240 112.560 24.270 ;
        RECT 114.230 22.000 114.520 26.585 ;
        RECT 116.320 22.290 116.610 27.620 ;
        RECT 118.470 26.585 118.640 26.810 ;
        RECT 118.410 22.000 118.700 26.585 ;
        RECT 120.500 22.290 120.790 27.620 ;
        RECT 122.650 26.585 122.820 26.810 ;
        RECT 122.590 22.000 122.880 26.585 ;
        RECT 125.045 24.720 125.215 28.645 ;
        RECT 125.555 24.720 125.845 28.790 ;
        RECT 127.645 25.085 127.940 29.350 ;
        RECT 125.045 24.690 127.140 24.720 ;
        RECT 125.045 24.600 127.295 24.690 ;
        RECT 128.275 24.600 128.445 28.635 ;
        RECT 129.955 28.200 130.455 29.350 ;
        RECT 125.045 24.430 128.445 24.600 ;
        RECT 125.045 24.270 127.295 24.430 ;
        RECT 125.045 24.240 127.140 24.270 ;
        RECT 129.940 22.000 130.230 26.345 ;
        RECT 132.025 22.305 132.320 30.895 ;
        RECT 134.120 30.710 134.410 35.120 ;
        RECT 134.750 30.705 134.920 35.120 ;
        RECT 137.080 33.245 137.370 37.840 ;
        RECT 137.140 33.000 137.310 33.245 ;
        RECT 137.290 30.790 138.420 31.790 ;
        RECT 139.170 31.480 139.460 37.540 ;
        RECT 141.260 33.245 141.550 37.840 ;
        RECT 141.320 33.000 141.490 33.245 ;
        RECT 143.350 31.580 143.640 37.540 ;
        RECT 145.440 33.245 145.730 37.840 ;
        RECT 147.400 35.455 149.745 35.600 ;
        RECT 150.545 35.455 152.890 35.600 ;
        RECT 147.400 35.285 152.890 35.455 ;
        RECT 147.400 35.120 149.745 35.285 ;
        RECT 150.545 35.120 152.890 35.285 ;
        RECT 145.500 33.235 145.695 33.245 ;
        RECT 145.500 33.000 145.670 33.235 ;
        RECT 143.350 31.480 144.170 31.580 ;
        RECT 139.170 30.980 144.170 31.480 ;
        RECT 132.940 28.860 134.120 29.060 ;
        RECT 132.940 28.260 134.620 28.860 ;
        RECT 132.940 27.980 134.120 28.260 ;
        RECT 134.120 22.000 134.410 26.345 ;
        RECT 136.570 24.720 136.740 29.575 ;
        RECT 137.080 24.720 137.370 29.570 ;
        RECT 139.170 25.030 139.460 30.980 ;
        RECT 147.400 30.460 147.570 35.120 ;
        RECT 147.910 30.290 148.200 35.120 ;
        RECT 150.000 29.850 150.290 34.850 ;
        RECT 152.090 30.290 152.380 35.120 ;
        RECT 152.720 30.520 152.890 35.120 ;
        RECT 155.055 33.490 155.345 37.840 ;
        RECT 155.290 31.580 156.490 31.890 ;
        RECT 154.790 30.960 156.490 31.580 ;
        RECT 155.290 30.760 156.490 30.960 ;
        RECT 157.140 29.850 157.435 37.530 ;
        RECT 159.235 33.490 159.525 37.840 ;
        RECT 162.325 35.570 164.420 35.600 ;
        RECT 162.170 35.405 164.420 35.570 ;
        RECT 161.020 35.235 164.420 35.405 ;
        RECT 161.020 32.260 161.190 35.235 ;
        RECT 162.170 35.150 164.420 35.235 ;
        RECT 162.325 35.120 164.420 35.150 ;
        RECT 161.525 31.675 161.820 34.750 ;
        RECT 161.295 30.895 162.035 31.675 ;
        RECT 141.260 24.720 141.550 29.570 ;
        RECT 141.890 24.720 142.060 29.575 ;
        RECT 147.360 29.350 159.955 29.850 ;
        RECT 147.360 27.910 147.860 29.350 ;
        RECT 148.890 28.320 152.890 28.920 ;
        RECT 150.890 28.200 152.890 28.320 ;
        RECT 145.820 27.620 150.290 27.910 ;
        RECT 150.890 27.620 152.090 28.200 ;
        RECT 143.790 26.595 143.960 26.830 ;
        RECT 143.765 26.585 143.960 26.595 ;
        RECT 136.570 24.595 138.915 24.720 ;
        RECT 139.715 24.690 142.060 24.720 ;
        RECT 139.715 24.595 142.240 24.690 ;
        RECT 136.570 24.425 142.240 24.595 ;
        RECT 136.570 24.240 138.915 24.425 ;
        RECT 139.715 24.270 142.240 24.425 ;
        RECT 139.715 24.240 142.060 24.270 ;
        RECT 143.730 22.000 144.020 26.585 ;
        RECT 145.820 22.290 146.110 27.620 ;
        RECT 147.970 26.585 148.140 26.810 ;
        RECT 147.910 22.000 148.200 26.585 ;
        RECT 150.000 22.290 150.290 27.620 ;
        RECT 152.150 26.585 152.320 26.810 ;
        RECT 152.090 22.000 152.380 26.585 ;
        RECT 154.545 24.720 154.715 28.645 ;
        RECT 155.055 24.720 155.345 28.790 ;
        RECT 157.145 25.085 157.440 29.350 ;
        RECT 154.545 24.690 156.640 24.720 ;
        RECT 154.545 24.600 156.795 24.690 ;
        RECT 157.775 24.600 157.945 28.635 ;
        RECT 159.455 28.200 159.955 29.350 ;
        RECT 154.545 24.430 157.945 24.600 ;
        RECT 154.545 24.270 156.795 24.430 ;
        RECT 154.545 24.240 156.640 24.270 ;
        RECT 159.440 22.000 159.730 26.345 ;
        RECT 161.525 22.305 161.820 30.895 ;
        RECT 163.620 30.710 163.910 35.120 ;
        RECT 164.250 30.705 164.420 35.120 ;
        RECT 162.440 28.860 163.620 29.060 ;
        RECT 162.440 28.260 164.120 28.860 ;
        RECT 162.440 27.980 163.620 28.260 ;
        RECT 163.620 22.000 163.910 26.345 ;
        RECT 172.420 26.200 174.420 26.370 ;
        RECT 172.500 26.170 174.340 26.200 ;
        RECT 175.550 25.740 177.550 25.910 ;
        RECT 175.630 25.710 177.470 25.740 ;
        RECT 25.220 21.520 27.570 22.000 ;
        RECT 28.620 21.520 31.480 22.000 ;
        RECT 32.545 21.520 34.890 22.000 ;
        RECT 40.930 21.970 43.270 22.000 ;
        RECT 44.080 21.970 46.420 22.000 ;
        RECT 40.930 21.550 43.275 21.970 ;
        RECT 44.075 21.550 46.420 21.970 ;
        RECT 40.930 21.520 43.270 21.550 ;
        RECT 44.080 21.520 46.420 21.550 ;
        RECT 54.720 21.520 57.070 22.000 ;
        RECT 58.120 21.520 60.980 22.000 ;
        RECT 62.045 21.520 64.390 22.000 ;
        RECT 70.430 21.970 72.770 22.000 ;
        RECT 73.580 21.970 75.920 22.000 ;
        RECT 70.430 21.550 72.775 21.970 ;
        RECT 73.575 21.550 75.920 21.970 ;
        RECT 70.430 21.520 72.770 21.550 ;
        RECT 73.580 21.520 75.920 21.550 ;
        RECT 84.220 21.520 86.570 22.000 ;
        RECT 87.620 21.520 90.480 22.000 ;
        RECT 91.545 21.520 93.890 22.000 ;
        RECT 99.930 21.970 102.270 22.000 ;
        RECT 103.080 21.970 105.420 22.000 ;
        RECT 99.930 21.550 102.275 21.970 ;
        RECT 103.075 21.550 105.420 21.970 ;
        RECT 99.930 21.520 102.270 21.550 ;
        RECT 103.080 21.520 105.420 21.550 ;
        RECT 113.720 21.520 116.070 22.000 ;
        RECT 117.120 21.520 119.980 22.000 ;
        RECT 121.045 21.520 123.390 22.000 ;
        RECT 129.430 21.970 131.770 22.000 ;
        RECT 132.580 21.970 134.920 22.000 ;
        RECT 129.430 21.550 131.775 21.970 ;
        RECT 132.575 21.550 134.920 21.970 ;
        RECT 129.430 21.520 131.770 21.550 ;
        RECT 132.580 21.520 134.920 21.550 ;
        RECT 143.220 21.520 145.570 22.000 ;
        RECT 146.620 21.520 149.480 22.000 ;
        RECT 150.545 21.520 152.890 22.000 ;
        RECT 158.930 21.970 161.270 22.000 ;
        RECT 162.080 21.970 164.420 22.000 ;
        RECT 158.930 21.550 161.275 21.970 ;
        RECT 162.075 21.550 164.420 21.970 ;
        RECT 172.500 21.820 174.340 21.850 ;
        RECT 172.420 21.650 174.420 21.820 ;
        RECT 158.930 21.520 161.270 21.550 ;
        RECT 162.080 21.520 164.420 21.550 ;
        RECT 175.630 21.360 177.470 21.390 ;
        RECT 175.550 21.190 177.550 21.360 ;
        RECT 2.970 16.530 5.310 16.560 ;
        RECT 6.120 16.530 8.460 16.560 ;
        RECT 2.970 16.110 5.315 16.530 ;
        RECT 6.115 16.110 8.460 16.530 ;
        RECT 2.970 16.080 5.310 16.110 ;
        RECT 6.120 16.080 8.460 16.110 ;
        RECT 14.500 16.080 16.845 16.560 ;
        RECT 17.910 16.080 20.770 16.560 ;
        RECT 21.820 16.080 24.170 16.560 ;
        RECT 32.470 16.530 34.810 16.560 ;
        RECT 35.620 16.530 37.960 16.560 ;
        RECT 32.470 16.110 34.815 16.530 ;
        RECT 35.615 16.110 37.960 16.530 ;
        RECT 32.470 16.080 34.810 16.110 ;
        RECT 35.620 16.080 37.960 16.110 ;
        RECT 44.000 16.080 46.345 16.560 ;
        RECT 47.410 16.080 50.270 16.560 ;
        RECT 51.320 16.080 53.670 16.560 ;
        RECT 61.970 16.530 64.310 16.560 ;
        RECT 65.120 16.530 67.460 16.560 ;
        RECT 61.970 16.110 64.315 16.530 ;
        RECT 65.115 16.110 67.460 16.530 ;
        RECT 61.970 16.080 64.310 16.110 ;
        RECT 65.120 16.080 67.460 16.110 ;
        RECT 73.500 16.080 75.845 16.560 ;
        RECT 76.910 16.080 79.770 16.560 ;
        RECT 80.820 16.080 83.170 16.560 ;
        RECT 91.470 16.530 93.810 16.560 ;
        RECT 94.620 16.530 96.960 16.560 ;
        RECT 91.470 16.110 93.815 16.530 ;
        RECT 94.615 16.110 96.960 16.530 ;
        RECT 91.470 16.080 93.810 16.110 ;
        RECT 94.620 16.080 96.960 16.110 ;
        RECT 103.000 16.080 105.345 16.560 ;
        RECT 106.410 16.080 109.270 16.560 ;
        RECT 110.320 16.080 112.670 16.560 ;
        RECT 120.970 16.530 123.310 16.560 ;
        RECT 124.120 16.530 126.460 16.560 ;
        RECT 120.970 16.110 123.315 16.530 ;
        RECT 124.115 16.110 126.460 16.530 ;
        RECT 120.970 16.080 123.310 16.110 ;
        RECT 124.120 16.080 126.460 16.110 ;
        RECT 132.500 16.080 134.845 16.560 ;
        RECT 135.910 16.080 138.770 16.560 ;
        RECT 139.820 16.080 142.170 16.560 ;
        RECT 150.470 16.530 152.810 16.560 ;
        RECT 153.620 16.530 155.960 16.560 ;
        RECT 150.470 16.110 152.815 16.530 ;
        RECT 153.615 16.110 155.960 16.530 ;
        RECT 150.470 16.080 152.810 16.110 ;
        RECT 153.620 16.080 155.960 16.110 ;
        RECT 162.000 16.080 164.345 16.560 ;
        RECT 165.410 16.080 168.270 16.560 ;
        RECT 169.320 16.080 171.670 16.560 ;
        RECT 3.480 11.735 3.770 16.080 ;
        RECT 3.770 9.820 4.950 10.100 ;
        RECT 3.270 9.220 4.950 9.820 ;
        RECT 3.770 9.020 4.950 9.220 ;
        RECT 2.970 2.960 3.140 7.375 ;
        RECT 3.480 2.960 3.770 7.370 ;
        RECT 5.570 7.185 5.865 15.775 ;
        RECT 7.660 11.735 7.950 16.080 ;
        RECT 10.750 13.810 12.845 13.840 ;
        RECT 10.595 13.650 12.845 13.810 ;
        RECT 9.445 13.480 12.845 13.650 ;
        RECT 7.435 8.730 7.935 9.880 ;
        RECT 9.445 9.445 9.615 13.480 ;
        RECT 10.595 13.390 12.845 13.480 ;
        RECT 10.750 13.360 12.845 13.390 ;
        RECT 9.950 8.730 10.245 12.995 ;
        RECT 12.045 9.290 12.335 13.360 ;
        RECT 12.675 9.435 12.845 13.360 ;
        RECT 15.010 11.495 15.300 16.080 ;
        RECT 15.070 11.270 15.240 11.495 ;
        RECT 17.100 10.460 17.390 15.790 ;
        RECT 19.190 11.495 19.480 16.080 ;
        RECT 19.250 11.270 19.420 11.495 ;
        RECT 21.280 10.460 21.570 15.790 ;
        RECT 23.370 11.495 23.660 16.080 ;
        RECT 25.330 13.810 27.675 13.840 ;
        RECT 25.150 13.655 27.675 13.810 ;
        RECT 28.475 13.655 30.820 13.840 ;
        RECT 25.150 13.485 30.820 13.655 ;
        RECT 25.150 13.390 27.675 13.485 ;
        RECT 25.330 13.360 27.675 13.390 ;
        RECT 28.475 13.360 30.820 13.485 ;
        RECT 23.430 11.485 23.625 11.495 ;
        RECT 23.430 11.250 23.600 11.485 ;
        RECT 15.300 9.880 16.500 10.460 ;
        RECT 17.100 10.170 21.570 10.460 ;
        RECT 14.500 9.760 16.500 9.880 ;
        RECT 14.500 9.160 18.500 9.760 ;
        RECT 19.530 8.730 20.030 10.170 ;
        RECT 7.435 8.230 20.030 8.730 ;
        RECT 25.330 8.505 25.500 13.360 ;
        RECT 25.840 8.510 26.130 13.360 ;
        RECT 5.355 6.405 6.095 7.185 ;
        RECT 5.570 3.330 5.865 6.405 ;
        RECT 2.970 2.930 5.065 2.960 ;
        RECT 2.970 2.845 5.220 2.930 ;
        RECT 6.200 2.845 6.370 5.820 ;
        RECT 2.970 2.675 6.370 2.845 ;
        RECT 2.970 2.510 5.220 2.675 ;
        RECT 2.970 2.480 5.065 2.510 ;
        RECT 7.865 0.240 8.155 4.590 ;
        RECT 9.955 0.550 10.250 8.230 ;
        RECT 10.900 7.120 12.100 7.320 ;
        RECT 10.900 6.500 12.600 7.120 ;
        RECT 10.900 6.190 12.100 6.500 ;
        RECT 12.045 0.240 12.335 4.590 ;
        RECT 14.500 2.960 14.670 7.560 ;
        RECT 15.010 2.960 15.300 7.790 ;
        RECT 17.100 3.230 17.390 8.230 ;
        RECT 19.190 2.960 19.480 7.790 ;
        RECT 19.820 2.960 19.990 7.620 ;
        RECT 27.930 7.100 28.220 13.050 ;
        RECT 30.020 8.510 30.310 13.360 ;
        RECT 30.650 8.505 30.820 13.360 ;
        RECT 32.980 11.735 33.270 16.080 ;
        RECT 33.270 9.820 34.450 10.100 ;
        RECT 32.770 9.220 34.450 9.820 ;
        RECT 33.270 9.020 34.450 9.220 ;
        RECT 23.220 6.600 28.220 7.100 ;
        RECT 23.220 6.500 24.040 6.600 ;
        RECT 21.720 4.845 21.890 5.080 ;
        RECT 21.695 4.835 21.890 4.845 ;
        RECT 14.500 2.795 16.845 2.960 ;
        RECT 17.645 2.795 19.990 2.960 ;
        RECT 14.500 2.625 19.990 2.795 ;
        RECT 14.500 2.480 16.845 2.625 ;
        RECT 17.645 2.480 19.990 2.625 ;
        RECT 21.660 0.240 21.950 4.835 ;
        RECT 23.750 0.540 24.040 6.500 ;
        RECT 25.900 4.835 26.070 5.080 ;
        RECT 25.840 0.240 26.130 4.835 ;
        RECT 27.930 0.540 28.220 6.600 ;
        RECT 28.970 6.290 30.100 7.290 ;
        RECT 30.080 4.835 30.250 5.080 ;
        RECT 30.020 0.240 30.310 4.835 ;
        RECT 32.470 2.960 32.640 7.375 ;
        RECT 32.980 2.960 33.270 7.370 ;
        RECT 35.070 7.185 35.365 15.775 ;
        RECT 37.160 11.735 37.450 16.080 ;
        RECT 40.250 13.810 42.345 13.840 ;
        RECT 40.095 13.650 42.345 13.810 ;
        RECT 38.945 13.480 42.345 13.650 ;
        RECT 36.935 8.730 37.435 9.880 ;
        RECT 38.945 9.445 39.115 13.480 ;
        RECT 40.095 13.390 42.345 13.480 ;
        RECT 40.250 13.360 42.345 13.390 ;
        RECT 39.450 8.730 39.745 12.995 ;
        RECT 41.545 9.290 41.835 13.360 ;
        RECT 42.175 9.435 42.345 13.360 ;
        RECT 44.510 11.495 44.800 16.080 ;
        RECT 44.570 11.270 44.740 11.495 ;
        RECT 46.600 10.460 46.890 15.790 ;
        RECT 48.690 11.495 48.980 16.080 ;
        RECT 48.750 11.270 48.920 11.495 ;
        RECT 50.780 10.460 51.070 15.790 ;
        RECT 52.870 11.495 53.160 16.080 ;
        RECT 54.830 13.810 57.175 13.840 ;
        RECT 54.650 13.655 57.175 13.810 ;
        RECT 57.975 13.655 60.320 13.840 ;
        RECT 54.650 13.485 60.320 13.655 ;
        RECT 54.650 13.390 57.175 13.485 ;
        RECT 54.830 13.360 57.175 13.390 ;
        RECT 57.975 13.360 60.320 13.485 ;
        RECT 52.930 11.485 53.125 11.495 ;
        RECT 52.930 11.250 53.100 11.485 ;
        RECT 44.800 9.880 46.000 10.460 ;
        RECT 46.600 10.170 51.070 10.460 ;
        RECT 44.000 9.760 46.000 9.880 ;
        RECT 44.000 9.160 48.000 9.760 ;
        RECT 49.030 8.730 49.530 10.170 ;
        RECT 36.935 8.230 49.530 8.730 ;
        RECT 54.830 8.505 55.000 13.360 ;
        RECT 55.340 8.510 55.630 13.360 ;
        RECT 34.855 6.405 35.595 7.185 ;
        RECT 35.070 3.330 35.365 6.405 ;
        RECT 32.470 2.930 34.565 2.960 ;
        RECT 32.470 2.845 34.720 2.930 ;
        RECT 35.700 2.845 35.870 5.820 ;
        RECT 32.470 2.675 35.870 2.845 ;
        RECT 32.470 2.510 34.720 2.675 ;
        RECT 32.470 2.480 34.565 2.510 ;
        RECT 37.365 0.240 37.655 4.590 ;
        RECT 39.455 0.550 39.750 8.230 ;
        RECT 40.400 7.120 41.600 7.320 ;
        RECT 40.400 6.500 42.100 7.120 ;
        RECT 40.400 6.190 41.600 6.500 ;
        RECT 41.545 0.240 41.835 4.590 ;
        RECT 44.000 2.960 44.170 7.560 ;
        RECT 44.510 2.960 44.800 7.790 ;
        RECT 46.600 3.230 46.890 8.230 ;
        RECT 48.690 2.960 48.980 7.790 ;
        RECT 49.320 2.960 49.490 7.620 ;
        RECT 57.430 7.100 57.720 13.050 ;
        RECT 59.520 8.510 59.810 13.360 ;
        RECT 60.150 8.505 60.320 13.360 ;
        RECT 62.480 11.735 62.770 16.080 ;
        RECT 62.770 9.820 63.950 10.100 ;
        RECT 62.270 9.220 63.950 9.820 ;
        RECT 62.770 9.020 63.950 9.220 ;
        RECT 52.720 6.600 57.720 7.100 ;
        RECT 52.720 6.500 53.540 6.600 ;
        RECT 51.220 4.845 51.390 5.080 ;
        RECT 51.195 4.835 51.390 4.845 ;
        RECT 44.000 2.795 46.345 2.960 ;
        RECT 47.145 2.795 49.490 2.960 ;
        RECT 44.000 2.625 49.490 2.795 ;
        RECT 44.000 2.480 46.345 2.625 ;
        RECT 47.145 2.480 49.490 2.625 ;
        RECT 51.160 0.240 51.450 4.835 ;
        RECT 53.250 0.540 53.540 6.500 ;
        RECT 55.400 4.835 55.570 5.080 ;
        RECT 55.340 0.240 55.630 4.835 ;
        RECT 57.430 0.540 57.720 6.600 ;
        RECT 58.470 6.290 59.600 7.290 ;
        RECT 59.580 4.835 59.750 5.080 ;
        RECT 59.520 0.240 59.810 4.835 ;
        RECT 61.970 2.960 62.140 7.375 ;
        RECT 62.480 2.960 62.770 7.370 ;
        RECT 64.570 7.185 64.865 15.775 ;
        RECT 66.660 11.735 66.950 16.080 ;
        RECT 69.750 13.810 71.845 13.840 ;
        RECT 69.595 13.650 71.845 13.810 ;
        RECT 68.445 13.480 71.845 13.650 ;
        RECT 66.435 8.730 66.935 9.880 ;
        RECT 68.445 9.445 68.615 13.480 ;
        RECT 69.595 13.390 71.845 13.480 ;
        RECT 69.750 13.360 71.845 13.390 ;
        RECT 68.950 8.730 69.245 12.995 ;
        RECT 71.045 9.290 71.335 13.360 ;
        RECT 71.675 9.435 71.845 13.360 ;
        RECT 74.010 11.495 74.300 16.080 ;
        RECT 74.070 11.270 74.240 11.495 ;
        RECT 76.100 10.460 76.390 15.790 ;
        RECT 78.190 11.495 78.480 16.080 ;
        RECT 78.250 11.270 78.420 11.495 ;
        RECT 80.280 10.460 80.570 15.790 ;
        RECT 82.370 11.495 82.660 16.080 ;
        RECT 84.330 13.810 86.675 13.840 ;
        RECT 84.150 13.655 86.675 13.810 ;
        RECT 87.475 13.655 89.820 13.840 ;
        RECT 84.150 13.485 89.820 13.655 ;
        RECT 84.150 13.390 86.675 13.485 ;
        RECT 84.330 13.360 86.675 13.390 ;
        RECT 87.475 13.360 89.820 13.485 ;
        RECT 82.430 11.485 82.625 11.495 ;
        RECT 82.430 11.250 82.600 11.485 ;
        RECT 74.300 9.880 75.500 10.460 ;
        RECT 76.100 10.170 80.570 10.460 ;
        RECT 73.500 9.760 75.500 9.880 ;
        RECT 73.500 9.160 77.500 9.760 ;
        RECT 78.530 8.730 79.030 10.170 ;
        RECT 66.435 8.230 79.030 8.730 ;
        RECT 84.330 8.505 84.500 13.360 ;
        RECT 84.840 8.510 85.130 13.360 ;
        RECT 64.355 6.405 65.095 7.185 ;
        RECT 64.570 3.330 64.865 6.405 ;
        RECT 61.970 2.930 64.065 2.960 ;
        RECT 61.970 2.845 64.220 2.930 ;
        RECT 65.200 2.845 65.370 5.820 ;
        RECT 61.970 2.675 65.370 2.845 ;
        RECT 61.970 2.510 64.220 2.675 ;
        RECT 61.970 2.480 64.065 2.510 ;
        RECT 66.865 0.240 67.155 4.590 ;
        RECT 68.955 0.550 69.250 8.230 ;
        RECT 69.900 7.120 71.100 7.320 ;
        RECT 69.900 6.500 71.600 7.120 ;
        RECT 69.900 6.190 71.100 6.500 ;
        RECT 71.045 0.240 71.335 4.590 ;
        RECT 73.500 2.960 73.670 7.560 ;
        RECT 74.010 2.960 74.300 7.790 ;
        RECT 76.100 3.230 76.390 8.230 ;
        RECT 78.190 2.960 78.480 7.790 ;
        RECT 78.820 2.960 78.990 7.620 ;
        RECT 86.930 7.100 87.220 13.050 ;
        RECT 89.020 8.510 89.310 13.360 ;
        RECT 89.650 8.505 89.820 13.360 ;
        RECT 91.980 11.735 92.270 16.080 ;
        RECT 92.270 9.820 93.450 10.100 ;
        RECT 91.770 9.220 93.450 9.820 ;
        RECT 92.270 9.020 93.450 9.220 ;
        RECT 82.220 6.600 87.220 7.100 ;
        RECT 82.220 6.500 83.040 6.600 ;
        RECT 80.720 4.845 80.890 5.080 ;
        RECT 80.695 4.835 80.890 4.845 ;
        RECT 73.500 2.795 75.845 2.960 ;
        RECT 76.645 2.795 78.990 2.960 ;
        RECT 73.500 2.625 78.990 2.795 ;
        RECT 73.500 2.480 75.845 2.625 ;
        RECT 76.645 2.480 78.990 2.625 ;
        RECT 80.660 0.240 80.950 4.835 ;
        RECT 82.750 0.540 83.040 6.500 ;
        RECT 84.900 4.835 85.070 5.080 ;
        RECT 84.840 0.240 85.130 4.835 ;
        RECT 86.930 0.540 87.220 6.600 ;
        RECT 87.970 6.290 89.100 7.290 ;
        RECT 89.080 4.835 89.250 5.080 ;
        RECT 89.020 0.240 89.310 4.835 ;
        RECT 91.470 2.960 91.640 7.375 ;
        RECT 91.980 2.960 92.270 7.370 ;
        RECT 94.070 7.185 94.365 15.775 ;
        RECT 96.160 11.735 96.450 16.080 ;
        RECT 99.250 13.810 101.345 13.840 ;
        RECT 99.095 13.650 101.345 13.810 ;
        RECT 97.945 13.480 101.345 13.650 ;
        RECT 95.935 8.730 96.435 9.880 ;
        RECT 97.945 9.445 98.115 13.480 ;
        RECT 99.095 13.390 101.345 13.480 ;
        RECT 99.250 13.360 101.345 13.390 ;
        RECT 98.450 8.730 98.745 12.995 ;
        RECT 100.545 9.290 100.835 13.360 ;
        RECT 101.175 9.435 101.345 13.360 ;
        RECT 103.510 11.495 103.800 16.080 ;
        RECT 103.570 11.270 103.740 11.495 ;
        RECT 105.600 10.460 105.890 15.790 ;
        RECT 107.690 11.495 107.980 16.080 ;
        RECT 107.750 11.270 107.920 11.495 ;
        RECT 109.780 10.460 110.070 15.790 ;
        RECT 111.870 11.495 112.160 16.080 ;
        RECT 113.830 13.810 116.175 13.840 ;
        RECT 113.650 13.655 116.175 13.810 ;
        RECT 116.975 13.655 119.320 13.840 ;
        RECT 113.650 13.485 119.320 13.655 ;
        RECT 113.650 13.390 116.175 13.485 ;
        RECT 113.830 13.360 116.175 13.390 ;
        RECT 116.975 13.360 119.320 13.485 ;
        RECT 111.930 11.485 112.125 11.495 ;
        RECT 111.930 11.250 112.100 11.485 ;
        RECT 103.800 9.880 105.000 10.460 ;
        RECT 105.600 10.170 110.070 10.460 ;
        RECT 103.000 9.760 105.000 9.880 ;
        RECT 103.000 9.160 107.000 9.760 ;
        RECT 108.030 8.730 108.530 10.170 ;
        RECT 95.935 8.230 108.530 8.730 ;
        RECT 113.830 8.505 114.000 13.360 ;
        RECT 114.340 8.510 114.630 13.360 ;
        RECT 93.855 6.405 94.595 7.185 ;
        RECT 94.070 3.330 94.365 6.405 ;
        RECT 91.470 2.930 93.565 2.960 ;
        RECT 91.470 2.845 93.720 2.930 ;
        RECT 94.700 2.845 94.870 5.820 ;
        RECT 91.470 2.675 94.870 2.845 ;
        RECT 91.470 2.510 93.720 2.675 ;
        RECT 91.470 2.480 93.565 2.510 ;
        RECT 96.365 0.240 96.655 4.590 ;
        RECT 98.455 0.550 98.750 8.230 ;
        RECT 99.400 7.120 100.600 7.320 ;
        RECT 99.400 6.500 101.100 7.120 ;
        RECT 99.400 6.190 100.600 6.500 ;
        RECT 100.545 0.240 100.835 4.590 ;
        RECT 103.000 2.960 103.170 7.560 ;
        RECT 103.510 2.960 103.800 7.790 ;
        RECT 105.600 3.230 105.890 8.230 ;
        RECT 107.690 2.960 107.980 7.790 ;
        RECT 108.320 2.960 108.490 7.620 ;
        RECT 116.430 7.100 116.720 13.050 ;
        RECT 118.520 8.510 118.810 13.360 ;
        RECT 119.150 8.505 119.320 13.360 ;
        RECT 121.480 11.735 121.770 16.080 ;
        RECT 121.770 9.820 122.950 10.100 ;
        RECT 121.270 9.220 122.950 9.820 ;
        RECT 121.770 9.020 122.950 9.220 ;
        RECT 111.720 6.600 116.720 7.100 ;
        RECT 111.720 6.500 112.540 6.600 ;
        RECT 110.220 4.845 110.390 5.080 ;
        RECT 110.195 4.835 110.390 4.845 ;
        RECT 103.000 2.795 105.345 2.960 ;
        RECT 106.145 2.795 108.490 2.960 ;
        RECT 103.000 2.625 108.490 2.795 ;
        RECT 103.000 2.480 105.345 2.625 ;
        RECT 106.145 2.480 108.490 2.625 ;
        RECT 110.160 0.240 110.450 4.835 ;
        RECT 112.250 0.540 112.540 6.500 ;
        RECT 114.400 4.835 114.570 5.080 ;
        RECT 114.340 0.240 114.630 4.835 ;
        RECT 116.430 0.540 116.720 6.600 ;
        RECT 117.470 6.290 118.600 7.290 ;
        RECT 118.580 4.835 118.750 5.080 ;
        RECT 118.520 0.240 118.810 4.835 ;
        RECT 120.970 2.960 121.140 7.375 ;
        RECT 121.480 2.960 121.770 7.370 ;
        RECT 123.570 7.185 123.865 15.775 ;
        RECT 125.660 11.735 125.950 16.080 ;
        RECT 128.750 13.810 130.845 13.840 ;
        RECT 128.595 13.650 130.845 13.810 ;
        RECT 127.445 13.480 130.845 13.650 ;
        RECT 125.435 8.730 125.935 9.880 ;
        RECT 127.445 9.445 127.615 13.480 ;
        RECT 128.595 13.390 130.845 13.480 ;
        RECT 128.750 13.360 130.845 13.390 ;
        RECT 127.950 8.730 128.245 12.995 ;
        RECT 130.045 9.290 130.335 13.360 ;
        RECT 130.675 9.435 130.845 13.360 ;
        RECT 133.010 11.495 133.300 16.080 ;
        RECT 133.070 11.270 133.240 11.495 ;
        RECT 135.100 10.460 135.390 15.790 ;
        RECT 137.190 11.495 137.480 16.080 ;
        RECT 137.250 11.270 137.420 11.495 ;
        RECT 139.280 10.460 139.570 15.790 ;
        RECT 141.370 11.495 141.660 16.080 ;
        RECT 143.330 13.810 145.675 13.840 ;
        RECT 143.150 13.655 145.675 13.810 ;
        RECT 146.475 13.655 148.820 13.840 ;
        RECT 143.150 13.485 148.820 13.655 ;
        RECT 143.150 13.390 145.675 13.485 ;
        RECT 143.330 13.360 145.675 13.390 ;
        RECT 146.475 13.360 148.820 13.485 ;
        RECT 141.430 11.485 141.625 11.495 ;
        RECT 141.430 11.250 141.600 11.485 ;
        RECT 133.300 9.880 134.500 10.460 ;
        RECT 135.100 10.170 139.570 10.460 ;
        RECT 132.500 9.760 134.500 9.880 ;
        RECT 132.500 9.160 136.500 9.760 ;
        RECT 137.530 8.730 138.030 10.170 ;
        RECT 125.435 8.230 138.030 8.730 ;
        RECT 143.330 8.505 143.500 13.360 ;
        RECT 143.840 8.510 144.130 13.360 ;
        RECT 123.355 6.405 124.095 7.185 ;
        RECT 123.570 3.330 123.865 6.405 ;
        RECT 120.970 2.930 123.065 2.960 ;
        RECT 120.970 2.845 123.220 2.930 ;
        RECT 124.200 2.845 124.370 5.820 ;
        RECT 120.970 2.675 124.370 2.845 ;
        RECT 120.970 2.510 123.220 2.675 ;
        RECT 120.970 2.480 123.065 2.510 ;
        RECT 125.865 0.240 126.155 4.590 ;
        RECT 127.955 0.550 128.250 8.230 ;
        RECT 128.900 7.120 130.100 7.320 ;
        RECT 128.900 6.500 130.600 7.120 ;
        RECT 128.900 6.190 130.100 6.500 ;
        RECT 130.045 0.240 130.335 4.590 ;
        RECT 132.500 2.960 132.670 7.560 ;
        RECT 133.010 2.960 133.300 7.790 ;
        RECT 135.100 3.230 135.390 8.230 ;
        RECT 137.190 2.960 137.480 7.790 ;
        RECT 137.820 2.960 137.990 7.620 ;
        RECT 145.930 7.100 146.220 13.050 ;
        RECT 148.020 8.510 148.310 13.360 ;
        RECT 148.650 8.505 148.820 13.360 ;
        RECT 150.980 11.735 151.270 16.080 ;
        RECT 151.270 9.820 152.450 10.100 ;
        RECT 150.770 9.220 152.450 9.820 ;
        RECT 151.270 9.020 152.450 9.220 ;
        RECT 141.220 6.600 146.220 7.100 ;
        RECT 141.220 6.500 142.040 6.600 ;
        RECT 139.720 4.845 139.890 5.080 ;
        RECT 139.695 4.835 139.890 4.845 ;
        RECT 132.500 2.795 134.845 2.960 ;
        RECT 135.645 2.795 137.990 2.960 ;
        RECT 132.500 2.625 137.990 2.795 ;
        RECT 132.500 2.480 134.845 2.625 ;
        RECT 135.645 2.480 137.990 2.625 ;
        RECT 139.660 0.240 139.950 4.835 ;
        RECT 141.750 0.540 142.040 6.500 ;
        RECT 143.900 4.835 144.070 5.080 ;
        RECT 143.840 0.240 144.130 4.835 ;
        RECT 145.930 0.540 146.220 6.600 ;
        RECT 146.970 6.290 148.100 7.290 ;
        RECT 148.080 4.835 148.250 5.080 ;
        RECT 148.020 0.240 148.310 4.835 ;
        RECT 150.470 2.960 150.640 7.375 ;
        RECT 150.980 2.960 151.270 7.370 ;
        RECT 153.070 7.185 153.365 15.775 ;
        RECT 155.160 11.735 155.450 16.080 ;
        RECT 158.250 13.810 160.345 13.840 ;
        RECT 158.095 13.650 160.345 13.810 ;
        RECT 156.945 13.480 160.345 13.650 ;
        RECT 154.935 8.730 155.435 9.880 ;
        RECT 156.945 9.445 157.115 13.480 ;
        RECT 158.095 13.390 160.345 13.480 ;
        RECT 158.250 13.360 160.345 13.390 ;
        RECT 157.450 8.730 157.745 12.995 ;
        RECT 159.545 9.290 159.835 13.360 ;
        RECT 160.175 9.435 160.345 13.360 ;
        RECT 162.510 11.495 162.800 16.080 ;
        RECT 162.570 11.270 162.740 11.495 ;
        RECT 164.600 10.460 164.890 15.790 ;
        RECT 166.690 11.495 166.980 16.080 ;
        RECT 166.750 11.270 166.920 11.495 ;
        RECT 168.780 10.460 169.070 15.790 ;
        RECT 170.870 11.495 171.160 16.080 ;
        RECT 172.830 13.810 175.175 13.840 ;
        RECT 172.650 13.655 175.175 13.810 ;
        RECT 175.975 13.655 178.320 13.840 ;
        RECT 172.650 13.485 178.320 13.655 ;
        RECT 172.650 13.390 175.175 13.485 ;
        RECT 172.830 13.360 175.175 13.390 ;
        RECT 175.975 13.360 178.320 13.485 ;
        RECT 170.930 11.485 171.125 11.495 ;
        RECT 170.930 11.250 171.100 11.485 ;
        RECT 162.800 9.880 164.000 10.460 ;
        RECT 164.600 10.170 169.070 10.460 ;
        RECT 162.000 9.760 164.000 9.880 ;
        RECT 162.000 9.160 166.000 9.760 ;
        RECT 167.030 8.730 167.530 10.170 ;
        RECT 154.935 8.230 167.530 8.730 ;
        RECT 172.830 8.505 173.000 13.360 ;
        RECT 173.340 8.510 173.630 13.360 ;
        RECT 152.855 6.405 153.595 7.185 ;
        RECT 153.070 3.330 153.365 6.405 ;
        RECT 150.470 2.930 152.565 2.960 ;
        RECT 150.470 2.845 152.720 2.930 ;
        RECT 153.700 2.845 153.870 5.820 ;
        RECT 150.470 2.675 153.870 2.845 ;
        RECT 150.470 2.510 152.720 2.675 ;
        RECT 150.470 2.480 152.565 2.510 ;
        RECT 155.365 0.240 155.655 4.590 ;
        RECT 157.455 0.550 157.750 8.230 ;
        RECT 158.400 7.120 159.600 7.320 ;
        RECT 158.400 6.500 160.100 7.120 ;
        RECT 158.400 6.190 159.600 6.500 ;
        RECT 159.545 0.240 159.835 4.590 ;
        RECT 162.000 2.960 162.170 7.560 ;
        RECT 162.510 2.960 162.800 7.790 ;
        RECT 164.600 3.230 164.890 8.230 ;
        RECT 166.690 2.960 166.980 7.790 ;
        RECT 167.320 2.960 167.490 7.620 ;
        RECT 175.430 7.100 175.720 13.050 ;
        RECT 177.520 8.510 177.810 13.360 ;
        RECT 178.150 8.505 178.320 13.360 ;
        RECT 170.720 6.600 175.720 7.100 ;
        RECT 170.720 6.500 171.540 6.600 ;
        RECT 169.220 4.845 169.390 5.080 ;
        RECT 169.195 4.835 169.390 4.845 ;
        RECT 162.000 2.795 164.345 2.960 ;
        RECT 165.145 2.795 167.490 2.960 ;
        RECT 162.000 2.625 167.490 2.795 ;
        RECT 162.000 2.480 164.345 2.625 ;
        RECT 165.145 2.480 167.490 2.625 ;
        RECT 169.160 0.240 169.450 4.835 ;
        RECT 171.250 0.540 171.540 6.500 ;
        RECT 173.400 4.835 173.570 5.080 ;
        RECT 173.340 0.240 173.630 4.835 ;
        RECT 175.430 0.540 175.720 6.600 ;
        RECT 176.470 6.290 177.600 7.290 ;
        RECT 177.580 4.835 177.750 5.080 ;
        RECT 177.520 0.240 177.810 4.835 ;
        RECT 7.355 -0.240 9.700 0.240 ;
        RECT 10.500 -0.240 12.845 0.240 ;
        RECT 21.150 -0.240 23.495 0.240 ;
        RECT 24.550 -0.240 27.410 0.240 ;
        RECT 28.475 -0.240 30.820 0.240 ;
        RECT 36.855 -0.240 39.200 0.240 ;
        RECT 40.000 -0.240 42.345 0.240 ;
        RECT 50.650 -0.240 52.995 0.240 ;
        RECT 54.050 -0.240 56.910 0.240 ;
        RECT 57.975 -0.240 60.320 0.240 ;
        RECT 66.355 -0.240 68.700 0.240 ;
        RECT 69.500 -0.240 71.845 0.240 ;
        RECT 80.150 -0.240 82.495 0.240 ;
        RECT 83.550 -0.240 86.410 0.240 ;
        RECT 87.475 -0.240 89.820 0.240 ;
        RECT 95.855 -0.240 98.200 0.240 ;
        RECT 99.000 -0.240 101.345 0.240 ;
        RECT 109.650 -0.240 111.995 0.240 ;
        RECT 113.050 -0.240 115.910 0.240 ;
        RECT 116.975 -0.240 119.320 0.240 ;
        RECT 125.355 -0.240 127.700 0.240 ;
        RECT 128.500 -0.240 130.845 0.240 ;
        RECT 139.150 -0.240 141.495 0.240 ;
        RECT 142.550 -0.240 145.410 0.240 ;
        RECT 146.475 -0.240 148.820 0.240 ;
        RECT 154.855 -0.240 157.200 0.240 ;
        RECT 158.000 -0.240 160.345 0.240 ;
        RECT 168.650 -0.240 170.995 0.240 ;
        RECT 172.050 -0.240 174.910 0.240 ;
        RECT 175.975 -0.240 178.320 0.240 ;
      LAYER mcon ;
        RECT 18.570 37.870 19.085 38.290 ;
        RECT 19.275 37.870 19.695 38.290 ;
        RECT 19.885 37.870 20.305 38.290 ;
        RECT 20.495 37.870 20.915 38.290 ;
        RECT 21.980 37.870 22.400 38.290 ;
        RECT 22.590 37.870 23.010 38.290 ;
        RECT 23.200 37.870 23.620 38.290 ;
        RECT 23.810 37.870 24.230 38.290 ;
        RECT 24.420 37.870 24.840 38.290 ;
        RECT 25.895 37.870 26.315 38.290 ;
        RECT 26.505 37.870 26.925 38.290 ;
        RECT 27.115 37.870 27.535 38.290 ;
        RECT 27.725 37.870 28.240 38.290 ;
        RECT 36.545 37.870 36.965 38.290 ;
        RECT 37.155 37.870 37.575 38.290 ;
        RECT 37.765 37.870 38.185 38.290 ;
        RECT 38.375 37.870 38.890 38.290 ;
        RECT 39.690 37.870 40.205 38.290 ;
        RECT 40.395 37.870 40.815 38.290 ;
        RECT 41.005 37.870 41.425 38.290 ;
        RECT 41.615 37.870 42.035 38.290 ;
        RECT 48.070 37.870 48.585 38.290 ;
        RECT 48.775 37.870 49.195 38.290 ;
        RECT 49.385 37.870 49.805 38.290 ;
        RECT 49.995 37.870 50.415 38.290 ;
        RECT 51.480 37.870 51.900 38.290 ;
        RECT 52.090 37.870 52.510 38.290 ;
        RECT 52.700 37.870 53.120 38.290 ;
        RECT 53.310 37.870 53.730 38.290 ;
        RECT 53.920 37.870 54.340 38.290 ;
        RECT 55.395 37.870 55.815 38.290 ;
        RECT 56.005 37.870 56.425 38.290 ;
        RECT 56.615 37.870 57.035 38.290 ;
        RECT 57.225 37.870 57.740 38.290 ;
        RECT 66.045 37.870 66.465 38.290 ;
        RECT 66.655 37.870 67.075 38.290 ;
        RECT 67.265 37.870 67.685 38.290 ;
        RECT 67.875 37.870 68.390 38.290 ;
        RECT 69.190 37.870 69.705 38.290 ;
        RECT 69.895 37.870 70.315 38.290 ;
        RECT 70.505 37.870 70.925 38.290 ;
        RECT 71.115 37.870 71.535 38.290 ;
        RECT 77.570 37.870 78.085 38.290 ;
        RECT 78.275 37.870 78.695 38.290 ;
        RECT 78.885 37.870 79.305 38.290 ;
        RECT 79.495 37.870 79.915 38.290 ;
        RECT 80.980 37.870 81.400 38.290 ;
        RECT 81.590 37.870 82.010 38.290 ;
        RECT 82.200 37.870 82.620 38.290 ;
        RECT 82.810 37.870 83.230 38.290 ;
        RECT 83.420 37.870 83.840 38.290 ;
        RECT 84.895 37.870 85.315 38.290 ;
        RECT 85.505 37.870 85.925 38.290 ;
        RECT 86.115 37.870 86.535 38.290 ;
        RECT 86.725 37.870 87.240 38.290 ;
        RECT 95.545 37.870 95.965 38.290 ;
        RECT 96.155 37.870 96.575 38.290 ;
        RECT 96.765 37.870 97.185 38.290 ;
        RECT 97.375 37.870 97.890 38.290 ;
        RECT 98.690 37.870 99.205 38.290 ;
        RECT 99.395 37.870 99.815 38.290 ;
        RECT 100.005 37.870 100.425 38.290 ;
        RECT 100.615 37.870 101.035 38.290 ;
        RECT 107.070 37.870 107.585 38.290 ;
        RECT 107.775 37.870 108.195 38.290 ;
        RECT 108.385 37.870 108.805 38.290 ;
        RECT 108.995 37.870 109.415 38.290 ;
        RECT 110.480 37.870 110.900 38.290 ;
        RECT 111.090 37.870 111.510 38.290 ;
        RECT 111.700 37.870 112.120 38.290 ;
        RECT 112.310 37.870 112.730 38.290 ;
        RECT 112.920 37.870 113.340 38.290 ;
        RECT 114.395 37.870 114.815 38.290 ;
        RECT 115.005 37.870 115.425 38.290 ;
        RECT 115.615 37.870 116.035 38.290 ;
        RECT 116.225 37.870 116.740 38.290 ;
        RECT 125.045 37.870 125.465 38.290 ;
        RECT 125.655 37.870 126.075 38.290 ;
        RECT 126.265 37.870 126.685 38.290 ;
        RECT 126.875 37.870 127.390 38.290 ;
        RECT 128.190 37.870 128.705 38.290 ;
        RECT 128.895 37.870 129.315 38.290 ;
        RECT 129.505 37.870 129.925 38.290 ;
        RECT 130.115 37.870 130.535 38.290 ;
        RECT 136.570 37.870 137.085 38.290 ;
        RECT 137.275 37.870 137.695 38.290 ;
        RECT 137.885 37.870 138.305 38.290 ;
        RECT 138.495 37.870 138.915 38.290 ;
        RECT 139.980 37.870 140.400 38.290 ;
        RECT 140.590 37.870 141.010 38.290 ;
        RECT 141.200 37.870 141.620 38.290 ;
        RECT 141.810 37.870 142.230 38.290 ;
        RECT 142.420 37.870 142.840 38.290 ;
        RECT 143.895 37.870 144.315 38.290 ;
        RECT 144.505 37.870 144.925 38.290 ;
        RECT 145.115 37.870 145.535 38.290 ;
        RECT 145.725 37.870 146.240 38.290 ;
        RECT 154.545 37.870 154.965 38.290 ;
        RECT 155.155 37.870 155.575 38.290 ;
        RECT 155.765 37.870 156.185 38.290 ;
        RECT 156.375 37.870 156.890 38.290 ;
        RECT 157.690 37.870 158.205 38.290 ;
        RECT 158.395 37.870 158.815 38.290 ;
        RECT 159.005 37.870 159.425 38.290 ;
        RECT 159.615 37.870 160.035 38.290 ;
        RECT 19.320 30.820 20.330 31.760 ;
        RECT 29.400 35.150 29.915 35.570 ;
        RECT 30.105 35.150 30.525 35.570 ;
        RECT 30.715 35.150 31.135 35.570 ;
        RECT 31.325 35.150 31.745 35.570 ;
        RECT 32.545 35.150 32.965 35.570 ;
        RECT 33.155 35.150 33.575 35.570 ;
        RECT 33.765 35.150 34.185 35.570 ;
        RECT 34.375 35.150 34.890 35.570 ;
        RECT 25.350 30.980 26.170 31.580 ;
        RECT 3.965 29.835 4.135 30.005 ;
        RECT 4.425 29.835 4.595 30.005 ;
        RECT 4.885 29.835 5.055 30.005 ;
        RECT 5.345 29.835 5.515 30.005 ;
        RECT 5.805 29.835 5.975 30.005 ;
        RECT 8.135 29.835 8.305 30.005 ;
        RECT 8.595 29.835 8.765 30.005 ;
        RECT 9.055 29.835 9.225 30.005 ;
        RECT 6.925 28.475 7.095 28.645 ;
        RECT 3.965 27.115 4.135 27.285 ;
        RECT 4.425 27.115 4.595 27.285 ;
        RECT 4.885 27.115 5.055 27.285 ;
        RECT 5.345 27.115 5.515 27.285 ;
        RECT 5.805 27.115 5.975 27.285 ;
        RECT 8.135 27.115 8.305 27.285 ;
        RECT 8.595 27.115 8.765 27.285 ;
        RECT 9.055 27.115 9.225 27.285 ;
        RECT 36.820 30.990 37.270 31.580 ;
        RECT 37.460 30.990 38.490 31.580 ;
        RECT 44.780 35.150 45.200 35.570 ;
        RECT 45.390 35.150 45.810 35.570 ;
        RECT 46.000 35.150 46.420 35.570 ;
        RECT 43.355 30.925 43.975 31.645 ;
        RECT 30.890 28.320 31.490 28.920 ;
        RECT 31.690 28.320 32.290 28.920 ;
        RECT 32.490 28.320 33.090 28.920 ;
        RECT 33.290 28.230 33.990 28.920 ;
        RECT 34.190 28.230 34.830 28.860 ;
        RECT 18.570 24.270 19.085 24.690 ;
        RECT 19.275 24.270 19.695 24.690 ;
        RECT 19.885 24.270 20.305 24.690 ;
        RECT 20.495 24.270 20.915 24.690 ;
        RECT 21.895 24.270 22.315 24.690 ;
        RECT 22.505 24.270 22.925 24.690 ;
        RECT 23.115 24.270 23.535 24.690 ;
        RECT 23.725 24.270 24.240 24.690 ;
        RECT 37.155 24.270 37.575 24.690 ;
        RECT 37.765 24.270 38.185 24.690 ;
        RECT 38.375 24.270 38.795 24.690 ;
        RECT 41.455 28.260 41.955 28.860 ;
        RECT 48.820 30.820 49.830 31.760 ;
        RECT 58.900 35.150 59.415 35.570 ;
        RECT 59.605 35.150 60.025 35.570 ;
        RECT 60.215 35.150 60.635 35.570 ;
        RECT 60.825 35.150 61.245 35.570 ;
        RECT 62.045 35.150 62.465 35.570 ;
        RECT 62.655 35.150 63.075 35.570 ;
        RECT 63.265 35.150 63.685 35.570 ;
        RECT 63.875 35.150 64.390 35.570 ;
        RECT 54.850 30.980 55.670 31.580 ;
        RECT 44.520 28.310 45.470 28.810 ;
        RECT 45.670 28.310 46.070 28.810 ;
        RECT 66.320 30.990 66.770 31.580 ;
        RECT 66.960 30.990 67.990 31.580 ;
        RECT 74.280 35.150 74.700 35.570 ;
        RECT 74.890 35.150 75.310 35.570 ;
        RECT 75.500 35.150 75.920 35.570 ;
        RECT 72.855 30.925 73.475 31.645 ;
        RECT 60.390 28.320 60.990 28.920 ;
        RECT 61.190 28.320 61.790 28.920 ;
        RECT 61.990 28.320 62.590 28.920 ;
        RECT 62.790 28.230 63.490 28.920 ;
        RECT 63.690 28.230 64.330 28.860 ;
        RECT 48.070 24.270 48.585 24.690 ;
        RECT 48.775 24.270 49.195 24.690 ;
        RECT 49.385 24.270 49.805 24.690 ;
        RECT 49.995 24.270 50.415 24.690 ;
        RECT 51.395 24.270 51.815 24.690 ;
        RECT 52.005 24.270 52.425 24.690 ;
        RECT 52.615 24.270 53.035 24.690 ;
        RECT 53.225 24.270 53.740 24.690 ;
        RECT 66.655 24.270 67.075 24.690 ;
        RECT 67.265 24.270 67.685 24.690 ;
        RECT 67.875 24.270 68.295 24.690 ;
        RECT 70.955 28.260 71.455 28.860 ;
        RECT 78.320 30.820 79.330 31.760 ;
        RECT 88.400 35.150 88.915 35.570 ;
        RECT 89.105 35.150 89.525 35.570 ;
        RECT 89.715 35.150 90.135 35.570 ;
        RECT 90.325 35.150 90.745 35.570 ;
        RECT 91.545 35.150 91.965 35.570 ;
        RECT 92.155 35.150 92.575 35.570 ;
        RECT 92.765 35.150 93.185 35.570 ;
        RECT 93.375 35.150 93.890 35.570 ;
        RECT 84.350 30.980 85.170 31.580 ;
        RECT 74.020 28.310 74.970 28.810 ;
        RECT 75.170 28.310 75.570 28.810 ;
        RECT 95.820 30.990 96.270 31.580 ;
        RECT 96.460 30.990 97.490 31.580 ;
        RECT 103.780 35.150 104.200 35.570 ;
        RECT 104.390 35.150 104.810 35.570 ;
        RECT 105.000 35.150 105.420 35.570 ;
        RECT 102.355 30.925 102.975 31.645 ;
        RECT 89.890 28.320 90.490 28.920 ;
        RECT 90.690 28.320 91.290 28.920 ;
        RECT 91.490 28.320 92.090 28.920 ;
        RECT 92.290 28.230 92.990 28.920 ;
        RECT 93.190 28.230 93.830 28.860 ;
        RECT 77.570 24.270 78.085 24.690 ;
        RECT 78.275 24.270 78.695 24.690 ;
        RECT 78.885 24.270 79.305 24.690 ;
        RECT 79.495 24.270 79.915 24.690 ;
        RECT 80.895 24.270 81.315 24.690 ;
        RECT 81.505 24.270 81.925 24.690 ;
        RECT 82.115 24.270 82.535 24.690 ;
        RECT 82.725 24.270 83.240 24.690 ;
        RECT 96.155 24.270 96.575 24.690 ;
        RECT 96.765 24.270 97.185 24.690 ;
        RECT 97.375 24.270 97.795 24.690 ;
        RECT 100.455 28.260 100.955 28.860 ;
        RECT 107.820 30.820 108.830 31.760 ;
        RECT 117.900 35.150 118.415 35.570 ;
        RECT 118.605 35.150 119.025 35.570 ;
        RECT 119.215 35.150 119.635 35.570 ;
        RECT 119.825 35.150 120.245 35.570 ;
        RECT 121.045 35.150 121.465 35.570 ;
        RECT 121.655 35.150 122.075 35.570 ;
        RECT 122.265 35.150 122.685 35.570 ;
        RECT 122.875 35.150 123.390 35.570 ;
        RECT 113.850 30.980 114.670 31.580 ;
        RECT 103.520 28.310 104.470 28.810 ;
        RECT 104.670 28.310 105.070 28.810 ;
        RECT 125.320 30.990 125.770 31.580 ;
        RECT 125.960 30.990 126.990 31.580 ;
        RECT 133.280 35.150 133.700 35.570 ;
        RECT 133.890 35.150 134.310 35.570 ;
        RECT 134.500 35.150 134.920 35.570 ;
        RECT 131.855 30.925 132.475 31.645 ;
        RECT 119.390 28.320 119.990 28.920 ;
        RECT 120.190 28.320 120.790 28.920 ;
        RECT 120.990 28.320 121.590 28.920 ;
        RECT 121.790 28.230 122.490 28.920 ;
        RECT 122.690 28.230 123.330 28.860 ;
        RECT 107.070 24.270 107.585 24.690 ;
        RECT 107.775 24.270 108.195 24.690 ;
        RECT 108.385 24.270 108.805 24.690 ;
        RECT 108.995 24.270 109.415 24.690 ;
        RECT 110.395 24.270 110.815 24.690 ;
        RECT 111.005 24.270 111.425 24.690 ;
        RECT 111.615 24.270 112.035 24.690 ;
        RECT 112.225 24.270 112.740 24.690 ;
        RECT 125.655 24.270 126.075 24.690 ;
        RECT 126.265 24.270 126.685 24.690 ;
        RECT 126.875 24.270 127.295 24.690 ;
        RECT 129.955 28.260 130.455 28.860 ;
        RECT 137.320 30.820 138.330 31.760 ;
        RECT 147.400 35.150 147.915 35.570 ;
        RECT 148.105 35.150 148.525 35.570 ;
        RECT 148.715 35.150 149.135 35.570 ;
        RECT 149.325 35.150 149.745 35.570 ;
        RECT 150.545 35.150 150.965 35.570 ;
        RECT 151.155 35.150 151.575 35.570 ;
        RECT 151.765 35.150 152.185 35.570 ;
        RECT 152.375 35.150 152.890 35.570 ;
        RECT 143.350 30.980 144.170 31.580 ;
        RECT 133.020 28.310 133.970 28.810 ;
        RECT 134.170 28.310 134.570 28.810 ;
        RECT 154.820 30.990 155.270 31.580 ;
        RECT 155.460 30.990 156.490 31.580 ;
        RECT 162.780 35.150 163.200 35.570 ;
        RECT 163.390 35.150 163.810 35.570 ;
        RECT 164.000 35.150 164.420 35.570 ;
        RECT 161.355 30.925 161.975 31.645 ;
        RECT 148.890 28.320 149.490 28.920 ;
        RECT 149.690 28.320 150.290 28.920 ;
        RECT 150.490 28.320 151.090 28.920 ;
        RECT 151.290 28.230 151.990 28.920 ;
        RECT 152.190 28.230 152.830 28.860 ;
        RECT 136.570 24.270 137.085 24.690 ;
        RECT 137.275 24.270 137.695 24.690 ;
        RECT 137.885 24.270 138.305 24.690 ;
        RECT 138.495 24.270 138.915 24.690 ;
        RECT 139.895 24.270 140.315 24.690 ;
        RECT 140.505 24.270 140.925 24.690 ;
        RECT 141.115 24.270 141.535 24.690 ;
        RECT 141.725 24.270 142.240 24.690 ;
        RECT 155.155 24.270 155.575 24.690 ;
        RECT 155.765 24.270 156.185 24.690 ;
        RECT 156.375 24.270 156.795 24.690 ;
        RECT 159.455 28.260 159.955 28.860 ;
        RECT 162.520 28.310 163.470 28.810 ;
        RECT 163.670 28.310 164.070 28.810 ;
        RECT 172.615 26.185 172.785 26.355 ;
        RECT 172.975 26.185 173.145 26.355 ;
        RECT 173.335 26.185 173.505 26.355 ;
        RECT 173.695 26.185 173.865 26.355 ;
        RECT 174.055 26.185 174.225 26.355 ;
        RECT 175.745 25.725 175.915 25.895 ;
        RECT 176.105 25.725 176.275 25.895 ;
        RECT 176.465 25.725 176.635 25.895 ;
        RECT 176.825 25.725 176.995 25.895 ;
        RECT 177.185 25.725 177.355 25.895 ;
        RECT 25.220 21.550 25.735 21.970 ;
        RECT 25.925 21.550 26.345 21.970 ;
        RECT 26.535 21.550 26.955 21.970 ;
        RECT 27.145 21.550 27.565 21.970 ;
        RECT 28.620 21.550 29.040 21.970 ;
        RECT 29.230 21.550 29.650 21.970 ;
        RECT 29.840 21.550 30.260 21.970 ;
        RECT 30.450 21.550 30.870 21.970 ;
        RECT 31.060 21.550 31.480 21.970 ;
        RECT 32.545 21.550 32.965 21.970 ;
        RECT 33.155 21.550 33.575 21.970 ;
        RECT 33.765 21.550 34.185 21.970 ;
        RECT 34.375 21.550 34.890 21.970 ;
        RECT 41.640 21.550 42.050 21.970 ;
        RECT 42.250 21.550 42.660 21.970 ;
        RECT 42.860 21.550 43.275 21.970 ;
        RECT 44.685 21.550 45.105 21.970 ;
        RECT 45.295 21.550 45.715 21.970 ;
        RECT 45.905 21.550 46.420 21.970 ;
        RECT 54.720 21.550 55.235 21.970 ;
        RECT 55.425 21.550 55.845 21.970 ;
        RECT 56.035 21.550 56.455 21.970 ;
        RECT 56.645 21.550 57.065 21.970 ;
        RECT 58.120 21.550 58.540 21.970 ;
        RECT 58.730 21.550 59.150 21.970 ;
        RECT 59.340 21.550 59.760 21.970 ;
        RECT 59.950 21.550 60.370 21.970 ;
        RECT 60.560 21.550 60.980 21.970 ;
        RECT 62.045 21.550 62.465 21.970 ;
        RECT 62.655 21.550 63.075 21.970 ;
        RECT 63.265 21.550 63.685 21.970 ;
        RECT 63.875 21.550 64.390 21.970 ;
        RECT 71.140 21.550 71.550 21.970 ;
        RECT 71.750 21.550 72.160 21.970 ;
        RECT 72.360 21.550 72.775 21.970 ;
        RECT 74.185 21.550 74.605 21.970 ;
        RECT 74.795 21.550 75.215 21.970 ;
        RECT 75.405 21.550 75.920 21.970 ;
        RECT 84.220 21.550 84.735 21.970 ;
        RECT 84.925 21.550 85.345 21.970 ;
        RECT 85.535 21.550 85.955 21.970 ;
        RECT 86.145 21.550 86.565 21.970 ;
        RECT 87.620 21.550 88.040 21.970 ;
        RECT 88.230 21.550 88.650 21.970 ;
        RECT 88.840 21.550 89.260 21.970 ;
        RECT 89.450 21.550 89.870 21.970 ;
        RECT 90.060 21.550 90.480 21.970 ;
        RECT 91.545 21.550 91.965 21.970 ;
        RECT 92.155 21.550 92.575 21.970 ;
        RECT 92.765 21.550 93.185 21.970 ;
        RECT 93.375 21.550 93.890 21.970 ;
        RECT 100.640 21.550 101.050 21.970 ;
        RECT 101.250 21.550 101.660 21.970 ;
        RECT 101.860 21.550 102.275 21.970 ;
        RECT 103.685 21.550 104.105 21.970 ;
        RECT 104.295 21.550 104.715 21.970 ;
        RECT 104.905 21.550 105.420 21.970 ;
        RECT 113.720 21.550 114.235 21.970 ;
        RECT 114.425 21.550 114.845 21.970 ;
        RECT 115.035 21.550 115.455 21.970 ;
        RECT 115.645 21.550 116.065 21.970 ;
        RECT 117.120 21.550 117.540 21.970 ;
        RECT 117.730 21.550 118.150 21.970 ;
        RECT 118.340 21.550 118.760 21.970 ;
        RECT 118.950 21.550 119.370 21.970 ;
        RECT 119.560 21.550 119.980 21.970 ;
        RECT 121.045 21.550 121.465 21.970 ;
        RECT 121.655 21.550 122.075 21.970 ;
        RECT 122.265 21.550 122.685 21.970 ;
        RECT 122.875 21.550 123.390 21.970 ;
        RECT 130.140 21.550 130.550 21.970 ;
        RECT 130.750 21.550 131.160 21.970 ;
        RECT 131.360 21.550 131.775 21.970 ;
        RECT 133.185 21.550 133.605 21.970 ;
        RECT 133.795 21.550 134.215 21.970 ;
        RECT 134.405 21.550 134.920 21.970 ;
        RECT 143.220 21.550 143.735 21.970 ;
        RECT 143.925 21.550 144.345 21.970 ;
        RECT 144.535 21.550 144.955 21.970 ;
        RECT 145.145 21.550 145.565 21.970 ;
        RECT 146.620 21.550 147.040 21.970 ;
        RECT 147.230 21.550 147.650 21.970 ;
        RECT 147.840 21.550 148.260 21.970 ;
        RECT 148.450 21.550 148.870 21.970 ;
        RECT 149.060 21.550 149.480 21.970 ;
        RECT 150.545 21.550 150.965 21.970 ;
        RECT 151.155 21.550 151.575 21.970 ;
        RECT 151.765 21.550 152.185 21.970 ;
        RECT 152.375 21.550 152.890 21.970 ;
        RECT 159.640 21.550 160.050 21.970 ;
        RECT 160.250 21.550 160.660 21.970 ;
        RECT 160.860 21.550 161.275 21.970 ;
        RECT 162.685 21.550 163.105 21.970 ;
        RECT 163.295 21.550 163.715 21.970 ;
        RECT 163.905 21.550 164.420 21.970 ;
        RECT 172.615 21.665 172.785 21.835 ;
        RECT 172.975 21.665 173.145 21.835 ;
        RECT 173.335 21.665 173.505 21.835 ;
        RECT 173.695 21.665 173.865 21.835 ;
        RECT 174.055 21.665 174.225 21.835 ;
        RECT 175.745 21.205 175.915 21.375 ;
        RECT 176.105 21.205 176.275 21.375 ;
        RECT 176.465 21.205 176.635 21.375 ;
        RECT 176.825 21.205 176.995 21.375 ;
        RECT 177.185 21.205 177.355 21.375 ;
        RECT 3.675 16.110 4.095 16.530 ;
        RECT 4.285 16.110 4.705 16.530 ;
        RECT 4.895 16.110 5.315 16.530 ;
        RECT 6.730 16.110 7.140 16.530 ;
        RECT 7.340 16.110 7.750 16.530 ;
        RECT 7.950 16.110 8.460 16.530 ;
        RECT 14.500 16.110 15.015 16.530 ;
        RECT 15.205 16.110 15.625 16.530 ;
        RECT 15.815 16.110 16.235 16.530 ;
        RECT 16.425 16.110 16.845 16.530 ;
        RECT 17.910 16.110 18.330 16.530 ;
        RECT 18.520 16.110 18.940 16.530 ;
        RECT 19.130 16.110 19.550 16.530 ;
        RECT 19.740 16.110 20.160 16.530 ;
        RECT 20.350 16.110 20.770 16.530 ;
        RECT 21.825 16.110 22.245 16.530 ;
        RECT 22.435 16.110 22.855 16.530 ;
        RECT 23.045 16.110 23.465 16.530 ;
        RECT 23.655 16.110 24.170 16.530 ;
        RECT 33.175 16.110 33.595 16.530 ;
        RECT 33.785 16.110 34.205 16.530 ;
        RECT 34.395 16.110 34.815 16.530 ;
        RECT 36.230 16.110 36.640 16.530 ;
        RECT 36.840 16.110 37.250 16.530 ;
        RECT 37.450 16.110 37.960 16.530 ;
        RECT 44.000 16.110 44.515 16.530 ;
        RECT 44.705 16.110 45.125 16.530 ;
        RECT 45.315 16.110 45.735 16.530 ;
        RECT 45.925 16.110 46.345 16.530 ;
        RECT 47.410 16.110 47.830 16.530 ;
        RECT 48.020 16.110 48.440 16.530 ;
        RECT 48.630 16.110 49.050 16.530 ;
        RECT 49.240 16.110 49.660 16.530 ;
        RECT 49.850 16.110 50.270 16.530 ;
        RECT 51.325 16.110 51.745 16.530 ;
        RECT 51.935 16.110 52.355 16.530 ;
        RECT 52.545 16.110 52.965 16.530 ;
        RECT 53.155 16.110 53.670 16.530 ;
        RECT 62.675 16.110 63.095 16.530 ;
        RECT 63.285 16.110 63.705 16.530 ;
        RECT 63.895 16.110 64.315 16.530 ;
        RECT 65.730 16.110 66.140 16.530 ;
        RECT 66.340 16.110 66.750 16.530 ;
        RECT 66.950 16.110 67.460 16.530 ;
        RECT 73.500 16.110 74.015 16.530 ;
        RECT 74.205 16.110 74.625 16.530 ;
        RECT 74.815 16.110 75.235 16.530 ;
        RECT 75.425 16.110 75.845 16.530 ;
        RECT 76.910 16.110 77.330 16.530 ;
        RECT 77.520 16.110 77.940 16.530 ;
        RECT 78.130 16.110 78.550 16.530 ;
        RECT 78.740 16.110 79.160 16.530 ;
        RECT 79.350 16.110 79.770 16.530 ;
        RECT 80.825 16.110 81.245 16.530 ;
        RECT 81.435 16.110 81.855 16.530 ;
        RECT 82.045 16.110 82.465 16.530 ;
        RECT 82.655 16.110 83.170 16.530 ;
        RECT 92.175 16.110 92.595 16.530 ;
        RECT 92.785 16.110 93.205 16.530 ;
        RECT 93.395 16.110 93.815 16.530 ;
        RECT 95.230 16.110 95.640 16.530 ;
        RECT 95.840 16.110 96.250 16.530 ;
        RECT 96.450 16.110 96.960 16.530 ;
        RECT 103.000 16.110 103.515 16.530 ;
        RECT 103.705 16.110 104.125 16.530 ;
        RECT 104.315 16.110 104.735 16.530 ;
        RECT 104.925 16.110 105.345 16.530 ;
        RECT 106.410 16.110 106.830 16.530 ;
        RECT 107.020 16.110 107.440 16.530 ;
        RECT 107.630 16.110 108.050 16.530 ;
        RECT 108.240 16.110 108.660 16.530 ;
        RECT 108.850 16.110 109.270 16.530 ;
        RECT 110.325 16.110 110.745 16.530 ;
        RECT 110.935 16.110 111.355 16.530 ;
        RECT 111.545 16.110 111.965 16.530 ;
        RECT 112.155 16.110 112.670 16.530 ;
        RECT 121.675 16.110 122.095 16.530 ;
        RECT 122.285 16.110 122.705 16.530 ;
        RECT 122.895 16.110 123.315 16.530 ;
        RECT 124.730 16.110 125.140 16.530 ;
        RECT 125.340 16.110 125.750 16.530 ;
        RECT 125.950 16.110 126.460 16.530 ;
        RECT 132.500 16.110 133.015 16.530 ;
        RECT 133.205 16.110 133.625 16.530 ;
        RECT 133.815 16.110 134.235 16.530 ;
        RECT 134.425 16.110 134.845 16.530 ;
        RECT 135.910 16.110 136.330 16.530 ;
        RECT 136.520 16.110 136.940 16.530 ;
        RECT 137.130 16.110 137.550 16.530 ;
        RECT 137.740 16.110 138.160 16.530 ;
        RECT 138.350 16.110 138.770 16.530 ;
        RECT 139.825 16.110 140.245 16.530 ;
        RECT 140.435 16.110 140.855 16.530 ;
        RECT 141.045 16.110 141.465 16.530 ;
        RECT 141.655 16.110 142.170 16.530 ;
        RECT 151.175 16.110 151.595 16.530 ;
        RECT 151.785 16.110 152.205 16.530 ;
        RECT 152.395 16.110 152.815 16.530 ;
        RECT 154.230 16.110 154.640 16.530 ;
        RECT 154.840 16.110 155.250 16.530 ;
        RECT 155.450 16.110 155.960 16.530 ;
        RECT 162.000 16.110 162.515 16.530 ;
        RECT 162.705 16.110 163.125 16.530 ;
        RECT 163.315 16.110 163.735 16.530 ;
        RECT 163.925 16.110 164.345 16.530 ;
        RECT 165.410 16.110 165.830 16.530 ;
        RECT 166.020 16.110 166.440 16.530 ;
        RECT 166.630 16.110 167.050 16.530 ;
        RECT 167.240 16.110 167.660 16.530 ;
        RECT 167.850 16.110 168.270 16.530 ;
        RECT 169.325 16.110 169.745 16.530 ;
        RECT 169.935 16.110 170.355 16.530 ;
        RECT 170.545 16.110 170.965 16.530 ;
        RECT 171.155 16.110 171.670 16.530 ;
        RECT 3.320 9.270 3.720 9.770 ;
        RECT 3.920 9.270 4.870 9.770 ;
        RECT 7.435 9.220 7.935 9.820 ;
        RECT 11.205 13.390 11.625 13.810 ;
        RECT 11.815 13.390 12.235 13.810 ;
        RECT 12.425 13.390 12.845 13.810 ;
        RECT 25.855 13.390 26.275 13.810 ;
        RECT 26.465 13.390 26.885 13.810 ;
        RECT 27.075 13.390 27.495 13.810 ;
        RECT 28.475 13.390 28.895 13.810 ;
        RECT 29.085 13.390 29.505 13.810 ;
        RECT 29.695 13.390 30.115 13.810 ;
        RECT 30.305 13.390 30.820 13.810 ;
        RECT 14.560 9.220 15.200 9.850 ;
        RECT 15.400 9.160 16.100 9.850 ;
        RECT 16.300 9.160 16.900 9.760 ;
        RECT 17.100 9.160 17.700 9.760 ;
        RECT 17.900 9.160 18.500 9.760 ;
        RECT 5.415 6.435 6.035 7.155 ;
        RECT 3.580 2.510 4.000 2.930 ;
        RECT 4.190 2.510 4.610 2.930 ;
        RECT 4.800 2.510 5.220 2.930 ;
        RECT 10.900 6.500 11.930 7.090 ;
        RECT 12.120 6.500 12.570 7.090 ;
        RECT 32.820 9.270 33.220 9.770 ;
        RECT 33.420 9.270 34.370 9.770 ;
        RECT 14.500 2.510 15.015 2.930 ;
        RECT 15.205 2.510 15.625 2.930 ;
        RECT 15.815 2.510 16.235 2.930 ;
        RECT 16.425 2.510 16.845 2.930 ;
        RECT 17.645 2.510 18.065 2.930 ;
        RECT 18.255 2.510 18.675 2.930 ;
        RECT 18.865 2.510 19.285 2.930 ;
        RECT 19.475 2.510 19.990 2.930 ;
        RECT 29.060 6.320 30.070 7.260 ;
        RECT 36.935 9.220 37.435 9.820 ;
        RECT 40.705 13.390 41.125 13.810 ;
        RECT 41.315 13.390 41.735 13.810 ;
        RECT 41.925 13.390 42.345 13.810 ;
        RECT 55.355 13.390 55.775 13.810 ;
        RECT 55.965 13.390 56.385 13.810 ;
        RECT 56.575 13.390 56.995 13.810 ;
        RECT 57.975 13.390 58.395 13.810 ;
        RECT 58.585 13.390 59.005 13.810 ;
        RECT 59.195 13.390 59.615 13.810 ;
        RECT 59.805 13.390 60.320 13.810 ;
        RECT 44.060 9.220 44.700 9.850 ;
        RECT 44.900 9.160 45.600 9.850 ;
        RECT 45.800 9.160 46.400 9.760 ;
        RECT 46.600 9.160 47.200 9.760 ;
        RECT 47.400 9.160 48.000 9.760 ;
        RECT 34.915 6.435 35.535 7.155 ;
        RECT 33.080 2.510 33.500 2.930 ;
        RECT 33.690 2.510 34.110 2.930 ;
        RECT 34.300 2.510 34.720 2.930 ;
        RECT 40.400 6.500 41.430 7.090 ;
        RECT 41.620 6.500 42.070 7.090 ;
        RECT 62.320 9.270 62.720 9.770 ;
        RECT 62.920 9.270 63.870 9.770 ;
        RECT 44.000 2.510 44.515 2.930 ;
        RECT 44.705 2.510 45.125 2.930 ;
        RECT 45.315 2.510 45.735 2.930 ;
        RECT 45.925 2.510 46.345 2.930 ;
        RECT 47.145 2.510 47.565 2.930 ;
        RECT 47.755 2.510 48.175 2.930 ;
        RECT 48.365 2.510 48.785 2.930 ;
        RECT 48.975 2.510 49.490 2.930 ;
        RECT 58.560 6.320 59.570 7.260 ;
        RECT 66.435 9.220 66.935 9.820 ;
        RECT 70.205 13.390 70.625 13.810 ;
        RECT 70.815 13.390 71.235 13.810 ;
        RECT 71.425 13.390 71.845 13.810 ;
        RECT 84.855 13.390 85.275 13.810 ;
        RECT 85.465 13.390 85.885 13.810 ;
        RECT 86.075 13.390 86.495 13.810 ;
        RECT 87.475 13.390 87.895 13.810 ;
        RECT 88.085 13.390 88.505 13.810 ;
        RECT 88.695 13.390 89.115 13.810 ;
        RECT 89.305 13.390 89.820 13.810 ;
        RECT 73.560 9.220 74.200 9.850 ;
        RECT 74.400 9.160 75.100 9.850 ;
        RECT 75.300 9.160 75.900 9.760 ;
        RECT 76.100 9.160 76.700 9.760 ;
        RECT 76.900 9.160 77.500 9.760 ;
        RECT 64.415 6.435 65.035 7.155 ;
        RECT 62.580 2.510 63.000 2.930 ;
        RECT 63.190 2.510 63.610 2.930 ;
        RECT 63.800 2.510 64.220 2.930 ;
        RECT 69.900 6.500 70.930 7.090 ;
        RECT 71.120 6.500 71.570 7.090 ;
        RECT 91.820 9.270 92.220 9.770 ;
        RECT 92.420 9.270 93.370 9.770 ;
        RECT 73.500 2.510 74.015 2.930 ;
        RECT 74.205 2.510 74.625 2.930 ;
        RECT 74.815 2.510 75.235 2.930 ;
        RECT 75.425 2.510 75.845 2.930 ;
        RECT 76.645 2.510 77.065 2.930 ;
        RECT 77.255 2.510 77.675 2.930 ;
        RECT 77.865 2.510 78.285 2.930 ;
        RECT 78.475 2.510 78.990 2.930 ;
        RECT 88.060 6.320 89.070 7.260 ;
        RECT 95.935 9.220 96.435 9.820 ;
        RECT 99.705 13.390 100.125 13.810 ;
        RECT 100.315 13.390 100.735 13.810 ;
        RECT 100.925 13.390 101.345 13.810 ;
        RECT 114.355 13.390 114.775 13.810 ;
        RECT 114.965 13.390 115.385 13.810 ;
        RECT 115.575 13.390 115.995 13.810 ;
        RECT 116.975 13.390 117.395 13.810 ;
        RECT 117.585 13.390 118.005 13.810 ;
        RECT 118.195 13.390 118.615 13.810 ;
        RECT 118.805 13.390 119.320 13.810 ;
        RECT 103.060 9.220 103.700 9.850 ;
        RECT 103.900 9.160 104.600 9.850 ;
        RECT 104.800 9.160 105.400 9.760 ;
        RECT 105.600 9.160 106.200 9.760 ;
        RECT 106.400 9.160 107.000 9.760 ;
        RECT 93.915 6.435 94.535 7.155 ;
        RECT 92.080 2.510 92.500 2.930 ;
        RECT 92.690 2.510 93.110 2.930 ;
        RECT 93.300 2.510 93.720 2.930 ;
        RECT 99.400 6.500 100.430 7.090 ;
        RECT 100.620 6.500 101.070 7.090 ;
        RECT 121.320 9.270 121.720 9.770 ;
        RECT 121.920 9.270 122.870 9.770 ;
        RECT 103.000 2.510 103.515 2.930 ;
        RECT 103.705 2.510 104.125 2.930 ;
        RECT 104.315 2.510 104.735 2.930 ;
        RECT 104.925 2.510 105.345 2.930 ;
        RECT 106.145 2.510 106.565 2.930 ;
        RECT 106.755 2.510 107.175 2.930 ;
        RECT 107.365 2.510 107.785 2.930 ;
        RECT 107.975 2.510 108.490 2.930 ;
        RECT 117.560 6.320 118.570 7.260 ;
        RECT 125.435 9.220 125.935 9.820 ;
        RECT 129.205 13.390 129.625 13.810 ;
        RECT 129.815 13.390 130.235 13.810 ;
        RECT 130.425 13.390 130.845 13.810 ;
        RECT 143.855 13.390 144.275 13.810 ;
        RECT 144.465 13.390 144.885 13.810 ;
        RECT 145.075 13.390 145.495 13.810 ;
        RECT 146.475 13.390 146.895 13.810 ;
        RECT 147.085 13.390 147.505 13.810 ;
        RECT 147.695 13.390 148.115 13.810 ;
        RECT 148.305 13.390 148.820 13.810 ;
        RECT 132.560 9.220 133.200 9.850 ;
        RECT 133.400 9.160 134.100 9.850 ;
        RECT 134.300 9.160 134.900 9.760 ;
        RECT 135.100 9.160 135.700 9.760 ;
        RECT 135.900 9.160 136.500 9.760 ;
        RECT 123.415 6.435 124.035 7.155 ;
        RECT 121.580 2.510 122.000 2.930 ;
        RECT 122.190 2.510 122.610 2.930 ;
        RECT 122.800 2.510 123.220 2.930 ;
        RECT 128.900 6.500 129.930 7.090 ;
        RECT 130.120 6.500 130.570 7.090 ;
        RECT 150.820 9.270 151.220 9.770 ;
        RECT 151.420 9.270 152.370 9.770 ;
        RECT 132.500 2.510 133.015 2.930 ;
        RECT 133.205 2.510 133.625 2.930 ;
        RECT 133.815 2.510 134.235 2.930 ;
        RECT 134.425 2.510 134.845 2.930 ;
        RECT 135.645 2.510 136.065 2.930 ;
        RECT 136.255 2.510 136.675 2.930 ;
        RECT 136.865 2.510 137.285 2.930 ;
        RECT 137.475 2.510 137.990 2.930 ;
        RECT 147.060 6.320 148.070 7.260 ;
        RECT 154.935 9.220 155.435 9.820 ;
        RECT 158.705 13.390 159.125 13.810 ;
        RECT 159.315 13.390 159.735 13.810 ;
        RECT 159.925 13.390 160.345 13.810 ;
        RECT 173.355 13.390 173.775 13.810 ;
        RECT 173.965 13.390 174.385 13.810 ;
        RECT 174.575 13.390 174.995 13.810 ;
        RECT 175.975 13.390 176.395 13.810 ;
        RECT 176.585 13.390 177.005 13.810 ;
        RECT 177.195 13.390 177.615 13.810 ;
        RECT 177.805 13.390 178.320 13.810 ;
        RECT 162.060 9.220 162.700 9.850 ;
        RECT 162.900 9.160 163.600 9.850 ;
        RECT 163.800 9.160 164.400 9.760 ;
        RECT 164.600 9.160 165.200 9.760 ;
        RECT 165.400 9.160 166.000 9.760 ;
        RECT 152.915 6.435 153.535 7.155 ;
        RECT 151.080 2.510 151.500 2.930 ;
        RECT 151.690 2.510 152.110 2.930 ;
        RECT 152.300 2.510 152.720 2.930 ;
        RECT 158.400 6.500 159.430 7.090 ;
        RECT 159.620 6.500 160.070 7.090 ;
        RECT 162.000 2.510 162.515 2.930 ;
        RECT 162.705 2.510 163.125 2.930 ;
        RECT 163.315 2.510 163.735 2.930 ;
        RECT 163.925 2.510 164.345 2.930 ;
        RECT 165.145 2.510 165.565 2.930 ;
        RECT 165.755 2.510 166.175 2.930 ;
        RECT 166.365 2.510 166.785 2.930 ;
        RECT 166.975 2.510 167.490 2.930 ;
        RECT 176.560 6.320 177.570 7.260 ;
        RECT 7.355 -0.210 7.775 0.210 ;
        RECT 7.965 -0.210 8.385 0.210 ;
        RECT 8.575 -0.210 8.995 0.210 ;
        RECT 9.185 -0.210 9.700 0.210 ;
        RECT 10.500 -0.210 11.015 0.210 ;
        RECT 11.205 -0.210 11.625 0.210 ;
        RECT 11.815 -0.210 12.235 0.210 ;
        RECT 12.425 -0.210 12.845 0.210 ;
        RECT 21.150 -0.210 21.665 0.210 ;
        RECT 21.855 -0.210 22.275 0.210 ;
        RECT 22.465 -0.210 22.885 0.210 ;
        RECT 23.075 -0.210 23.495 0.210 ;
        RECT 24.550 -0.210 24.970 0.210 ;
        RECT 25.160 -0.210 25.580 0.210 ;
        RECT 25.770 -0.210 26.190 0.210 ;
        RECT 26.380 -0.210 26.800 0.210 ;
        RECT 26.990 -0.210 27.410 0.210 ;
        RECT 28.475 -0.210 28.895 0.210 ;
        RECT 29.085 -0.210 29.505 0.210 ;
        RECT 29.695 -0.210 30.115 0.210 ;
        RECT 30.305 -0.210 30.820 0.210 ;
        RECT 36.855 -0.210 37.275 0.210 ;
        RECT 37.465 -0.210 37.885 0.210 ;
        RECT 38.075 -0.210 38.495 0.210 ;
        RECT 38.685 -0.210 39.200 0.210 ;
        RECT 40.000 -0.210 40.515 0.210 ;
        RECT 40.705 -0.210 41.125 0.210 ;
        RECT 41.315 -0.210 41.735 0.210 ;
        RECT 41.925 -0.210 42.345 0.210 ;
        RECT 50.650 -0.210 51.165 0.210 ;
        RECT 51.355 -0.210 51.775 0.210 ;
        RECT 51.965 -0.210 52.385 0.210 ;
        RECT 52.575 -0.210 52.995 0.210 ;
        RECT 54.050 -0.210 54.470 0.210 ;
        RECT 54.660 -0.210 55.080 0.210 ;
        RECT 55.270 -0.210 55.690 0.210 ;
        RECT 55.880 -0.210 56.300 0.210 ;
        RECT 56.490 -0.210 56.910 0.210 ;
        RECT 57.975 -0.210 58.395 0.210 ;
        RECT 58.585 -0.210 59.005 0.210 ;
        RECT 59.195 -0.210 59.615 0.210 ;
        RECT 59.805 -0.210 60.320 0.210 ;
        RECT 66.355 -0.210 66.775 0.210 ;
        RECT 66.965 -0.210 67.385 0.210 ;
        RECT 67.575 -0.210 67.995 0.210 ;
        RECT 68.185 -0.210 68.700 0.210 ;
        RECT 69.500 -0.210 70.015 0.210 ;
        RECT 70.205 -0.210 70.625 0.210 ;
        RECT 70.815 -0.210 71.235 0.210 ;
        RECT 71.425 -0.210 71.845 0.210 ;
        RECT 80.150 -0.210 80.665 0.210 ;
        RECT 80.855 -0.210 81.275 0.210 ;
        RECT 81.465 -0.210 81.885 0.210 ;
        RECT 82.075 -0.210 82.495 0.210 ;
        RECT 83.550 -0.210 83.970 0.210 ;
        RECT 84.160 -0.210 84.580 0.210 ;
        RECT 84.770 -0.210 85.190 0.210 ;
        RECT 85.380 -0.210 85.800 0.210 ;
        RECT 85.990 -0.210 86.410 0.210 ;
        RECT 87.475 -0.210 87.895 0.210 ;
        RECT 88.085 -0.210 88.505 0.210 ;
        RECT 88.695 -0.210 89.115 0.210 ;
        RECT 89.305 -0.210 89.820 0.210 ;
        RECT 95.855 -0.210 96.275 0.210 ;
        RECT 96.465 -0.210 96.885 0.210 ;
        RECT 97.075 -0.210 97.495 0.210 ;
        RECT 97.685 -0.210 98.200 0.210 ;
        RECT 99.000 -0.210 99.515 0.210 ;
        RECT 99.705 -0.210 100.125 0.210 ;
        RECT 100.315 -0.210 100.735 0.210 ;
        RECT 100.925 -0.210 101.345 0.210 ;
        RECT 109.650 -0.210 110.165 0.210 ;
        RECT 110.355 -0.210 110.775 0.210 ;
        RECT 110.965 -0.210 111.385 0.210 ;
        RECT 111.575 -0.210 111.995 0.210 ;
        RECT 113.050 -0.210 113.470 0.210 ;
        RECT 113.660 -0.210 114.080 0.210 ;
        RECT 114.270 -0.210 114.690 0.210 ;
        RECT 114.880 -0.210 115.300 0.210 ;
        RECT 115.490 -0.210 115.910 0.210 ;
        RECT 116.975 -0.210 117.395 0.210 ;
        RECT 117.585 -0.210 118.005 0.210 ;
        RECT 118.195 -0.210 118.615 0.210 ;
        RECT 118.805 -0.210 119.320 0.210 ;
        RECT 125.355 -0.210 125.775 0.210 ;
        RECT 125.965 -0.210 126.385 0.210 ;
        RECT 126.575 -0.210 126.995 0.210 ;
        RECT 127.185 -0.210 127.700 0.210 ;
        RECT 128.500 -0.210 129.015 0.210 ;
        RECT 129.205 -0.210 129.625 0.210 ;
        RECT 129.815 -0.210 130.235 0.210 ;
        RECT 130.425 -0.210 130.845 0.210 ;
        RECT 139.150 -0.210 139.665 0.210 ;
        RECT 139.855 -0.210 140.275 0.210 ;
        RECT 140.465 -0.210 140.885 0.210 ;
        RECT 141.075 -0.210 141.495 0.210 ;
        RECT 142.550 -0.210 142.970 0.210 ;
        RECT 143.160 -0.210 143.580 0.210 ;
        RECT 143.770 -0.210 144.190 0.210 ;
        RECT 144.380 -0.210 144.800 0.210 ;
        RECT 144.990 -0.210 145.410 0.210 ;
        RECT 146.475 -0.210 146.895 0.210 ;
        RECT 147.085 -0.210 147.505 0.210 ;
        RECT 147.695 -0.210 148.115 0.210 ;
        RECT 148.305 -0.210 148.820 0.210 ;
        RECT 154.855 -0.210 155.275 0.210 ;
        RECT 155.465 -0.210 155.885 0.210 ;
        RECT 156.075 -0.210 156.495 0.210 ;
        RECT 156.685 -0.210 157.200 0.210 ;
        RECT 158.000 -0.210 158.515 0.210 ;
        RECT 158.705 -0.210 159.125 0.210 ;
        RECT 159.315 -0.210 159.735 0.210 ;
        RECT 159.925 -0.210 160.345 0.210 ;
        RECT 168.650 -0.210 169.165 0.210 ;
        RECT 169.355 -0.210 169.775 0.210 ;
        RECT 169.965 -0.210 170.385 0.210 ;
        RECT 170.575 -0.210 170.995 0.210 ;
        RECT 172.050 -0.210 172.470 0.210 ;
        RECT 172.660 -0.210 173.080 0.210 ;
        RECT 173.270 -0.210 173.690 0.210 ;
        RECT 173.880 -0.210 174.300 0.210 ;
        RECT 174.490 -0.210 174.910 0.210 ;
        RECT 175.975 -0.210 176.395 0.210 ;
        RECT 176.585 -0.210 177.005 0.210 ;
        RECT 177.195 -0.210 177.615 0.210 ;
        RECT 177.805 -0.210 178.320 0.210 ;
      LAYER met1 ;
        RECT 16.280 37.840 173.490 38.320 ;
        RECT 16.000 35.120 165.390 35.600 ;
        RECT 19.290 31.615 20.420 31.840 ;
        RECT 43.295 31.615 44.035 31.675 ;
        RECT 48.790 31.615 49.920 31.840 ;
        RECT 72.795 31.615 73.535 31.675 ;
        RECT 78.290 31.615 79.420 31.840 ;
        RECT 102.295 31.615 103.035 31.675 ;
        RECT 107.790 31.615 108.920 31.840 ;
        RECT 131.795 31.615 132.535 31.675 ;
        RECT 137.290 31.615 138.420 31.840 ;
        RECT 161.295 31.615 162.035 31.675 ;
        RECT 17.840 30.955 20.420 31.615 ;
        RECT 35.060 31.610 49.920 31.615 ;
        RECT 64.560 31.610 79.420 31.615 ;
        RECT 94.060 31.610 108.920 31.615 ;
        RECT 123.560 31.610 138.420 31.615 ;
        RECT 153.060 31.610 165.440 31.615 ;
        RECT 19.290 30.740 20.420 30.955 ;
        RECT 25.290 30.955 49.920 31.610 ;
        RECT 25.290 30.950 38.550 30.955 ;
        RECT 43.295 30.895 44.035 30.955 ;
        RECT 48.790 30.740 49.920 30.955 ;
        RECT 54.790 30.955 79.420 31.610 ;
        RECT 54.790 30.950 68.050 30.955 ;
        RECT 72.795 30.895 73.535 30.955 ;
        RECT 78.290 30.740 79.420 30.955 ;
        RECT 84.290 30.955 108.920 31.610 ;
        RECT 84.290 30.950 97.550 30.955 ;
        RECT 102.295 30.895 103.035 30.955 ;
        RECT 107.790 30.740 108.920 30.955 ;
        RECT 113.790 30.955 138.420 31.610 ;
        RECT 113.790 30.950 127.050 30.955 ;
        RECT 131.795 30.895 132.535 30.955 ;
        RECT 137.290 30.740 138.420 30.955 ;
        RECT 143.290 30.955 165.440 31.610 ;
        RECT 143.290 30.950 156.550 30.955 ;
        RECT 161.295 30.895 162.035 30.955 ;
        RECT 3.820 29.680 20.290 30.160 ;
        RECT 30.790 28.920 34.090 28.950 ;
        RECT 60.290 28.920 63.590 28.950 ;
        RECT 89.790 28.920 93.090 28.950 ;
        RECT 119.290 28.920 122.590 28.950 ;
        RECT 148.790 28.920 152.090 28.950 ;
        RECT 30.790 28.860 34.890 28.920 ;
        RECT 6.800 28.710 7.220 28.740 ;
        RECT 17.000 28.710 34.890 28.860 ;
        RECT 6.800 28.410 34.890 28.710 ;
        RECT 6.800 28.380 7.220 28.410 ;
        RECT 17.000 28.260 34.890 28.410 ;
        RECT 30.790 28.200 34.890 28.260 ;
        RECT 41.425 28.860 41.985 28.920 ;
        RECT 60.290 28.860 64.390 28.920 ;
        RECT 41.425 28.260 64.390 28.860 ;
        RECT 41.425 28.200 41.985 28.260 ;
        RECT 60.290 28.200 64.390 28.260 ;
        RECT 70.925 28.860 71.485 28.920 ;
        RECT 89.790 28.860 93.890 28.920 ;
        RECT 70.925 28.260 93.890 28.860 ;
        RECT 70.925 28.200 71.485 28.260 ;
        RECT 89.790 28.200 93.890 28.260 ;
        RECT 100.425 28.860 100.985 28.920 ;
        RECT 119.290 28.860 123.390 28.920 ;
        RECT 100.425 28.260 123.390 28.860 ;
        RECT 100.425 28.200 100.985 28.260 ;
        RECT 119.290 28.200 123.390 28.260 ;
        RECT 129.925 28.860 130.485 28.920 ;
        RECT 148.790 28.860 152.890 28.920 ;
        RECT 129.925 28.260 152.890 28.860 ;
        RECT 129.925 28.200 130.485 28.260 ;
        RECT 148.790 28.200 152.890 28.260 ;
        RECT 159.425 28.860 159.985 28.920 ;
        RECT 159.425 28.260 165.440 28.860 ;
        RECT 159.425 28.200 159.985 28.260 ;
        RECT 0.000 26.960 9.965 27.440 ;
        RECT 171.590 26.960 178.550 27.440 ;
        RECT 172.440 26.140 174.400 26.960 ;
        RECT 175.520 25.680 177.580 25.940 ;
        RECT 15.005 24.240 172.440 24.720 ;
        RECT 17.890 21.990 165.390 22.000 ;
        RECT 17.000 21.510 177.530 21.990 ;
        RECT 175.570 21.160 177.530 21.510 ;
        RECT 2.000 16.080 180.440 16.560 ;
        RECT 0.000 13.360 179.440 13.840 ;
        RECT 7.405 9.820 7.965 9.880 ;
        RECT 2.000 9.220 7.965 9.820 ;
        RECT 7.405 9.160 7.965 9.220 ;
        RECT 14.500 9.820 18.600 9.880 ;
        RECT 36.905 9.820 37.465 9.880 ;
        RECT 14.500 9.220 37.465 9.820 ;
        RECT 14.500 9.160 18.600 9.220 ;
        RECT 36.905 9.160 37.465 9.220 ;
        RECT 44.000 9.820 48.100 9.880 ;
        RECT 66.405 9.820 66.965 9.880 ;
        RECT 44.000 9.220 66.965 9.820 ;
        RECT 44.000 9.160 48.100 9.220 ;
        RECT 66.405 9.160 66.965 9.220 ;
        RECT 73.500 9.820 77.600 9.880 ;
        RECT 95.905 9.820 96.465 9.880 ;
        RECT 73.500 9.220 96.465 9.820 ;
        RECT 73.500 9.160 77.600 9.220 ;
        RECT 95.905 9.160 96.465 9.220 ;
        RECT 103.000 9.820 107.100 9.880 ;
        RECT 125.405 9.820 125.965 9.880 ;
        RECT 103.000 9.220 125.965 9.820 ;
        RECT 103.000 9.160 107.100 9.220 ;
        RECT 125.405 9.160 125.965 9.220 ;
        RECT 132.500 9.820 136.600 9.880 ;
        RECT 154.905 9.820 155.465 9.880 ;
        RECT 132.500 9.220 155.465 9.820 ;
        RECT 132.500 9.160 136.600 9.220 ;
        RECT 154.905 9.160 155.465 9.220 ;
        RECT 162.000 9.820 166.100 9.880 ;
        RECT 162.000 9.220 179.000 9.820 ;
        RECT 162.000 9.160 166.100 9.220 ;
        RECT 15.300 9.130 18.600 9.160 ;
        RECT 44.800 9.130 48.100 9.160 ;
        RECT 74.300 9.130 77.600 9.160 ;
        RECT 103.800 9.130 107.100 9.160 ;
        RECT 133.300 9.130 136.600 9.160 ;
        RECT 162.800 9.130 166.100 9.160 ;
        RECT 5.355 7.125 6.095 7.185 ;
        RECT 10.840 7.125 24.100 7.130 ;
        RECT 2.000 6.470 24.100 7.125 ;
        RECT 28.970 7.125 30.100 7.340 ;
        RECT 34.855 7.125 35.595 7.185 ;
        RECT 40.340 7.125 53.600 7.130 ;
        RECT 28.970 6.470 53.600 7.125 ;
        RECT 58.470 7.125 59.600 7.340 ;
        RECT 64.355 7.125 65.095 7.185 ;
        RECT 69.840 7.125 83.100 7.130 ;
        RECT 58.470 6.470 83.100 7.125 ;
        RECT 87.970 7.125 89.100 7.340 ;
        RECT 93.855 7.125 94.595 7.185 ;
        RECT 99.340 7.125 112.600 7.130 ;
        RECT 87.970 6.470 112.600 7.125 ;
        RECT 117.470 7.125 118.600 7.340 ;
        RECT 123.355 7.125 124.095 7.185 ;
        RECT 128.840 7.125 142.100 7.130 ;
        RECT 117.470 6.470 142.100 7.125 ;
        RECT 146.970 7.125 148.100 7.340 ;
        RECT 152.855 7.125 153.595 7.185 ;
        RECT 158.340 7.125 171.600 7.130 ;
        RECT 146.970 6.470 171.600 7.125 ;
        RECT 176.470 7.125 177.600 7.340 ;
        RECT 176.470 7.095 179.000 7.125 ;
        RECT 172.640 6.495 179.000 7.095 ;
        RECT 2.000 6.465 14.330 6.470 ;
        RECT 28.970 6.465 43.830 6.470 ;
        RECT 58.470 6.465 73.330 6.470 ;
        RECT 87.970 6.465 102.830 6.470 ;
        RECT 117.470 6.465 132.330 6.470 ;
        RECT 146.970 6.465 161.830 6.470 ;
        RECT 176.470 6.465 179.000 6.495 ;
        RECT 5.355 6.405 6.095 6.465 ;
        RECT 28.970 6.240 30.100 6.465 ;
        RECT 34.855 6.405 35.595 6.465 ;
        RECT 58.470 6.240 59.600 6.465 ;
        RECT 64.355 6.405 65.095 6.465 ;
        RECT 87.970 6.240 89.100 6.465 ;
        RECT 93.855 6.405 94.595 6.465 ;
        RECT 117.470 6.240 118.600 6.465 ;
        RECT 123.355 6.405 124.095 6.465 ;
        RECT 146.970 6.240 148.100 6.465 ;
        RECT 152.855 6.405 153.595 6.465 ;
        RECT 176.470 6.240 177.600 6.465 ;
        RECT 0.000 2.480 179.440 2.960 ;
        RECT 2.000 -0.240 180.440 0.240 ;
      LAYER via ;
        RECT 39.000 37.940 39.260 38.200 ;
        RECT 39.370 37.940 39.630 38.200 ;
        RECT 39.740 37.940 40.000 38.200 ;
        RECT 70.000 37.940 70.260 38.200 ;
        RECT 70.370 37.940 70.630 38.200 ;
        RECT 70.740 37.940 71.000 38.200 ;
        RECT 112.000 37.940 112.260 38.200 ;
        RECT 112.370 37.940 112.630 38.200 ;
        RECT 112.740 37.940 113.000 38.200 ;
        RECT 143.000 37.940 143.260 38.200 ;
        RECT 143.370 37.940 143.630 38.200 ;
        RECT 143.740 37.940 144.000 38.200 ;
        RECT 172.490 37.950 172.750 38.210 ;
        RECT 172.810 37.950 173.070 38.210 ;
        RECT 173.130 37.950 173.390 38.210 ;
        RECT 18.045 30.995 18.625 31.575 ;
        RECT 164.480 30.995 165.380 31.575 ;
        RECT 17.925 28.270 18.825 28.850 ;
        RECT 46.560 28.270 47.140 28.850 ;
        RECT 47.300 28.270 47.880 28.850 ;
        RECT 76.060 28.270 76.640 28.850 ;
        RECT 76.800 28.270 77.380 28.850 ;
        RECT 105.560 28.270 106.140 28.850 ;
        RECT 106.300 28.270 106.880 28.850 ;
        RECT 135.060 28.270 135.640 28.850 ;
        RECT 135.800 28.270 136.380 28.850 ;
        RECT 164.470 28.270 165.370 28.850 ;
        RECT 175.620 25.680 175.880 25.940 ;
        RECT 175.940 25.680 176.200 25.940 ;
        RECT 176.260 25.680 176.520 25.940 ;
        RECT 176.580 25.680 176.840 25.940 ;
        RECT 176.900 25.680 177.160 25.940 ;
        RECT 177.220 25.680 177.480 25.940 ;
        RECT 39.000 21.620 39.260 21.880 ;
        RECT 39.370 21.620 39.630 21.880 ;
        RECT 39.740 21.620 40.000 21.880 ;
        RECT 70.000 21.620 70.260 21.880 ;
        RECT 70.370 21.620 70.630 21.880 ;
        RECT 70.740 21.620 71.000 21.880 ;
        RECT 112.000 21.620 112.260 21.880 ;
        RECT 112.370 21.620 112.630 21.880 ;
        RECT 112.740 21.620 113.000 21.880 ;
        RECT 143.000 21.620 143.260 21.880 ;
        RECT 143.370 21.620 143.630 21.880 ;
        RECT 143.740 21.620 144.000 21.880 ;
        RECT 172.470 21.650 172.730 21.910 ;
        RECT 172.830 21.650 173.090 21.910 ;
        RECT 173.190 21.650 173.450 21.910 ;
        RECT 173.550 21.650 173.810 21.910 ;
        RECT 173.920 21.650 174.180 21.910 ;
        RECT 174.280 21.650 174.540 21.910 ;
        RECT 174.660 21.650 174.920 21.910 ;
        RECT 175.035 21.650 175.295 21.910 ;
        RECT 175.415 21.650 175.675 21.910 ;
        RECT 175.790 21.650 176.050 21.910 ;
        RECT 176.165 21.650 176.425 21.910 ;
        RECT 176.535 21.650 176.795 21.910 ;
        RECT 176.915 21.650 177.175 21.910 ;
        RECT 39.000 16.180 39.260 16.440 ;
        RECT 39.370 16.180 39.630 16.440 ;
        RECT 39.740 16.180 40.000 16.440 ;
        RECT 70.000 16.180 70.260 16.440 ;
        RECT 70.370 16.180 70.630 16.440 ;
        RECT 70.740 16.180 71.000 16.440 ;
        RECT 112.000 16.180 112.260 16.440 ;
        RECT 112.370 16.180 112.630 16.440 ;
        RECT 112.740 16.180 113.000 16.440 ;
        RECT 143.000 16.180 143.260 16.440 ;
        RECT 143.370 16.180 143.630 16.440 ;
        RECT 143.740 16.180 144.000 16.440 ;
        RECT 179.465 16.190 179.725 16.450 ;
        RECT 179.785 16.190 180.045 16.450 ;
        RECT 180.105 16.190 180.365 16.450 ;
        RECT 6.765 9.230 7.345 9.810 ;
        RECT 31.010 9.230 31.590 9.810 ;
        RECT 31.750 9.230 32.330 9.810 ;
        RECT 60.510 9.230 61.090 9.810 ;
        RECT 61.250 9.230 61.830 9.810 ;
        RECT 90.010 9.230 90.590 9.810 ;
        RECT 90.750 9.230 91.330 9.810 ;
        RECT 119.510 9.230 120.090 9.810 ;
        RECT 120.250 9.230 120.830 9.810 ;
        RECT 149.010 9.230 149.590 9.810 ;
        RECT 149.750 9.230 150.330 9.810 ;
        RECT 166.150 9.230 166.730 9.810 ;
        RECT 166.870 9.230 167.450 9.810 ;
        RECT 4.055 6.505 4.635 7.085 ;
        RECT 172.760 6.505 173.340 7.085 ;
        RECT 39.000 -0.140 39.260 0.120 ;
        RECT 39.370 -0.140 39.630 0.120 ;
        RECT 39.740 -0.140 40.000 0.120 ;
        RECT 70.000 -0.140 70.260 0.120 ;
        RECT 70.370 -0.140 70.630 0.120 ;
        RECT 70.740 -0.140 71.000 0.120 ;
        RECT 112.000 -0.140 112.260 0.120 ;
        RECT 112.370 -0.140 112.630 0.120 ;
        RECT 112.740 -0.140 113.000 0.120 ;
        RECT 143.000 -0.140 143.260 0.120 ;
        RECT 143.370 -0.140 143.630 0.120 ;
        RECT 143.740 -0.140 144.000 0.120 ;
        RECT 179.475 -0.130 179.735 0.130 ;
        RECT 179.795 -0.130 180.055 0.130 ;
        RECT 180.115 -0.130 180.375 0.130 ;
      LAYER met2 ;
        RECT 39.000 37.870 40.000 38.270 ;
        RECT 17.890 31.635 18.785 31.665 ;
        RECT 14.420 30.935 18.785 31.635 ;
        RECT 14.420 20.050 15.120 30.935 ;
        RECT 17.890 30.905 18.785 30.935 ;
        RECT 46.820 28.920 47.620 39.370 ;
        RECT 70.000 37.870 71.000 38.270 ;
        RECT 76.320 28.920 77.120 39.370 ;
        RECT 105.820 28.920 106.620 39.370 ;
        RECT 112.000 37.870 113.000 38.270 ;
        RECT 135.320 28.920 136.120 39.370 ;
        RECT 143.000 37.870 144.000 38.270 ;
        RECT 164.470 31.635 165.390 31.665 ;
        RECT 164.470 30.935 169.490 31.635 ;
        RECT 164.470 30.905 165.390 30.935 ;
        RECT 4.000 19.350 15.120 20.050 ;
        RECT 17.120 28.210 18.865 28.910 ;
        RECT 46.550 28.210 47.890 28.920 ;
        RECT 76.050 28.210 77.390 28.920 ;
        RECT 105.550 28.210 106.890 28.920 ;
        RECT 135.050 28.210 136.390 28.920 ;
        RECT 164.450 28.210 166.790 28.910 ;
        RECT 4.000 18.535 4.700 19.350 ;
        RECT 3.995 12.965 4.700 18.535 ;
        RECT 17.120 17.350 17.820 28.210 ;
        RECT 39.000 21.550 40.000 21.950 ;
        RECT 70.000 21.550 71.000 21.950 ;
        RECT 112.000 21.550 113.000 21.950 ;
        RECT 143.000 21.550 144.000 21.950 ;
        RECT 6.705 16.650 17.820 17.350 ;
        RECT 3.995 6.415 4.695 12.965 ;
        RECT 6.705 9.170 7.405 16.650 ;
        RECT 13.270 -1.290 14.070 16.650 ;
        RECT 39.000 16.110 40.000 16.510 ;
        RECT 70.000 16.110 71.000 16.510 ;
        RECT 112.000 16.110 113.000 16.510 ;
        RECT 143.000 16.110 144.000 16.510 ;
        RECT 166.090 9.870 166.790 28.210 ;
        RECT 168.790 17.635 169.490 30.935 ;
        RECT 172.440 22.240 173.440 38.370 ;
        RECT 175.570 25.390 181.500 26.190 ;
        RECT 172.440 21.240 180.440 22.240 ;
        RECT 179.440 20.700 180.435 21.240 ;
        RECT 168.790 16.935 173.400 17.635 ;
        RECT 31.000 9.190 32.340 9.870 ;
        RECT 60.500 9.190 61.840 9.870 ;
        RECT 90.000 9.190 91.340 9.870 ;
        RECT 119.500 9.190 120.840 9.870 ;
        RECT 149.000 9.190 150.340 9.870 ;
        RECT 31.270 -1.290 32.070 9.190 ;
        RECT 39.000 -0.210 40.000 0.190 ;
        RECT 60.770 -1.290 61.570 9.190 ;
        RECT 70.000 -0.210 71.000 0.190 ;
        RECT 90.270 -1.290 91.070 9.190 ;
        RECT 112.000 -0.210 113.000 0.190 ;
        RECT 119.770 -1.290 120.570 9.190 ;
        RECT 143.000 -0.210 144.000 0.190 ;
        RECT 149.270 -1.290 150.070 9.190 ;
        RECT 166.090 9.140 167.460 9.870 ;
        RECT 166.360 -1.290 167.160 9.140 ;
        RECT 172.700 6.445 173.400 16.935 ;
        RECT 179.440 -0.290 180.440 20.700 ;
      LAYER via2 ;
        RECT 39.100 37.920 39.400 38.220 ;
        RECT 39.600 37.920 39.900 38.220 ;
        RECT 70.100 37.920 70.400 38.220 ;
        RECT 70.600 37.920 70.900 38.220 ;
        RECT 112.100 37.920 112.400 38.220 ;
        RECT 112.600 37.920 112.900 38.220 ;
        RECT 143.100 37.920 143.400 38.220 ;
        RECT 143.600 37.920 143.900 38.220 ;
        RECT 39.100 21.600 39.400 21.900 ;
        RECT 39.600 21.600 39.900 21.900 ;
        RECT 70.100 21.600 70.400 21.900 ;
        RECT 70.600 21.600 70.900 21.900 ;
        RECT 112.100 21.600 112.400 21.900 ;
        RECT 112.600 21.600 112.900 21.900 ;
        RECT 143.100 21.600 143.400 21.900 ;
        RECT 143.600 21.600 143.900 21.900 ;
        RECT 39.100 16.160 39.400 16.460 ;
        RECT 39.600 16.160 39.900 16.460 ;
        RECT 70.100 16.160 70.400 16.460 ;
        RECT 70.600 16.160 70.900 16.460 ;
        RECT 112.100 16.160 112.400 16.460 ;
        RECT 112.600 16.160 112.900 16.460 ;
        RECT 143.100 16.160 143.400 16.460 ;
        RECT 143.600 16.160 143.900 16.460 ;
        RECT 179.750 19.100 180.150 19.500 ;
        RECT 179.750 18.570 180.150 18.970 ;
        RECT 39.100 -0.160 39.400 0.140 ;
        RECT 39.600 -0.160 39.900 0.140 ;
        RECT 70.100 -0.160 70.400 0.140 ;
        RECT 70.600 -0.160 70.900 0.140 ;
        RECT 112.100 -0.160 112.400 0.140 ;
        RECT 112.600 -0.160 112.900 0.140 ;
        RECT 143.100 -0.160 143.400 0.140 ;
        RECT 143.600 -0.160 143.900 0.140 ;
      LAYER met3 ;
        RECT 39.000 19.610 40.000 38.320 ;
        RECT 70.000 19.610 71.000 38.320 ;
        RECT 112.000 19.610 113.000 38.320 ;
        RECT 143.000 19.610 144.000 38.320 ;
        RECT 39.000 18.460 180.440 19.610 ;
        RECT 39.000 -0.240 40.000 18.460 ;
        RECT 70.000 -0.240 71.000 18.460 ;
        RECT 112.000 -0.240 113.000 18.460 ;
        RECT 143.000 -0.240 144.000 18.460 ;
  END
END ring_osc_r100
MACRO pwell_co_ring
  CLASS BLOCK ;
  FOREIGN pwell_co_ring ;
  ORIGIN -0.880 -30.000 ;
  SIZE 179.740 BY 42.500 ;
  OBS
      LAYER li1 ;
        RECT 15.920 72.000 166.580 72.500 ;
        RECT 16.000 52.500 16.500 72.000 ;
        RECT 166.000 52.500 166.500 72.000 ;
        RECT 15.920 52.000 166.580 52.500 ;
        RECT 0.920 50.000 180.580 50.500 ;
        RECT 1.000 30.500 1.500 50.000 ;
        RECT 180.000 30.500 180.500 50.000 ;
        RECT 0.920 30.000 180.580 30.500 ;
  END
END pwell_co_ring
MACRO power_ring_2_2
  CLASS BLOCK ;
  FOREIGN power_ring_2_2 ;
  ORIGIN -135.000 -16.000 ;
  SIZE 182.000 BY 105.000 ;
  OBS
      LAYER met3 ;
        RECT 140.000 119.000 312.000 121.000 ;
        RECT 135.000 115.000 317.000 117.000 ;
        RECT 135.000 20.000 317.000 22.000 ;
        RECT 140.000 16.000 312.000 18.000 ;
      LAYER via3 ;
        RECT 140.200 120.400 140.600 120.800 ;
        RECT 140.800 120.400 141.200 120.800 ;
        RECT 141.400 120.400 141.800 120.800 ;
        RECT 153.200 120.400 153.600 120.800 ;
        RECT 153.800 120.400 154.200 120.800 ;
        RECT 154.400 120.400 154.800 120.800 ;
        RECT 189.200 120.400 189.600 120.800 ;
        RECT 189.800 120.400 190.200 120.800 ;
        RECT 190.400 120.400 190.800 120.800 ;
        RECT 225.200 120.400 225.600 120.800 ;
        RECT 225.800 120.400 226.200 120.800 ;
        RECT 226.400 120.400 226.800 120.800 ;
        RECT 261.200 120.400 261.600 120.800 ;
        RECT 261.800 120.400 262.200 120.800 ;
        RECT 262.400 120.400 262.800 120.800 ;
        RECT 297.200 120.400 297.600 120.800 ;
        RECT 297.800 120.400 298.200 120.800 ;
        RECT 298.400 120.400 298.800 120.800 ;
        RECT 310.200 120.400 310.600 120.800 ;
        RECT 310.800 120.400 311.200 120.800 ;
        RECT 311.400 120.400 311.800 120.800 ;
        RECT 140.200 119.800 140.600 120.200 ;
        RECT 140.800 119.800 141.200 120.200 ;
        RECT 141.400 119.800 141.800 120.200 ;
        RECT 153.200 119.800 153.600 120.200 ;
        RECT 153.800 119.800 154.200 120.200 ;
        RECT 154.400 119.800 154.800 120.200 ;
        RECT 189.200 119.800 189.600 120.200 ;
        RECT 189.800 119.800 190.200 120.200 ;
        RECT 190.400 119.800 190.800 120.200 ;
        RECT 225.200 119.800 225.600 120.200 ;
        RECT 225.800 119.800 226.200 120.200 ;
        RECT 226.400 119.800 226.800 120.200 ;
        RECT 261.200 119.800 261.600 120.200 ;
        RECT 261.800 119.800 262.200 120.200 ;
        RECT 262.400 119.800 262.800 120.200 ;
        RECT 297.200 119.800 297.600 120.200 ;
        RECT 297.800 119.800 298.200 120.200 ;
        RECT 298.400 119.800 298.800 120.200 ;
        RECT 310.200 119.800 310.600 120.200 ;
        RECT 310.800 119.800 311.200 120.200 ;
        RECT 311.400 119.800 311.800 120.200 ;
        RECT 140.200 119.200 140.600 119.600 ;
        RECT 140.800 119.200 141.200 119.600 ;
        RECT 141.400 119.200 141.800 119.600 ;
        RECT 153.200 119.200 153.600 119.600 ;
        RECT 153.800 119.200 154.200 119.600 ;
        RECT 154.400 119.200 154.800 119.600 ;
        RECT 189.200 119.200 189.600 119.600 ;
        RECT 189.800 119.200 190.200 119.600 ;
        RECT 190.400 119.200 190.800 119.600 ;
        RECT 225.200 119.200 225.600 119.600 ;
        RECT 225.800 119.200 226.200 119.600 ;
        RECT 226.400 119.200 226.800 119.600 ;
        RECT 261.200 119.200 261.600 119.600 ;
        RECT 261.800 119.200 262.200 119.600 ;
        RECT 262.400 119.200 262.800 119.600 ;
        RECT 297.200 119.200 297.600 119.600 ;
        RECT 297.800 119.200 298.200 119.600 ;
        RECT 298.400 119.200 298.800 119.600 ;
        RECT 310.200 119.200 310.600 119.600 ;
        RECT 310.800 119.200 311.200 119.600 ;
        RECT 311.400 119.200 311.800 119.600 ;
        RECT 135.200 116.400 135.600 116.800 ;
        RECT 135.800 116.400 136.200 116.800 ;
        RECT 136.400 116.400 136.800 116.800 ;
        RECT 171.200 116.400 171.600 116.800 ;
        RECT 171.800 116.400 172.200 116.800 ;
        RECT 172.400 116.400 172.800 116.800 ;
        RECT 207.200 116.400 207.600 116.800 ;
        RECT 207.800 116.400 208.200 116.800 ;
        RECT 208.400 116.400 208.800 116.800 ;
        RECT 243.200 116.400 243.600 116.800 ;
        RECT 243.800 116.400 244.200 116.800 ;
        RECT 244.400 116.400 244.800 116.800 ;
        RECT 279.200 116.400 279.600 116.800 ;
        RECT 279.800 116.400 280.200 116.800 ;
        RECT 280.400 116.400 280.800 116.800 ;
        RECT 315.200 116.400 315.600 116.800 ;
        RECT 315.800 116.400 316.200 116.800 ;
        RECT 316.400 116.400 316.800 116.800 ;
        RECT 135.200 115.800 135.600 116.200 ;
        RECT 135.800 115.800 136.200 116.200 ;
        RECT 136.400 115.800 136.800 116.200 ;
        RECT 171.200 115.800 171.600 116.200 ;
        RECT 171.800 115.800 172.200 116.200 ;
        RECT 172.400 115.800 172.800 116.200 ;
        RECT 207.200 115.800 207.600 116.200 ;
        RECT 207.800 115.800 208.200 116.200 ;
        RECT 208.400 115.800 208.800 116.200 ;
        RECT 243.200 115.800 243.600 116.200 ;
        RECT 243.800 115.800 244.200 116.200 ;
        RECT 244.400 115.800 244.800 116.200 ;
        RECT 279.200 115.800 279.600 116.200 ;
        RECT 279.800 115.800 280.200 116.200 ;
        RECT 280.400 115.800 280.800 116.200 ;
        RECT 315.200 115.800 315.600 116.200 ;
        RECT 315.800 115.800 316.200 116.200 ;
        RECT 316.400 115.800 316.800 116.200 ;
        RECT 135.200 115.200 135.600 115.600 ;
        RECT 135.800 115.200 136.200 115.600 ;
        RECT 136.400 115.200 136.800 115.600 ;
        RECT 171.200 115.200 171.600 115.600 ;
        RECT 171.800 115.200 172.200 115.600 ;
        RECT 172.400 115.200 172.800 115.600 ;
        RECT 207.200 115.200 207.600 115.600 ;
        RECT 207.800 115.200 208.200 115.600 ;
        RECT 208.400 115.200 208.800 115.600 ;
        RECT 243.200 115.200 243.600 115.600 ;
        RECT 243.800 115.200 244.200 115.600 ;
        RECT 244.400 115.200 244.800 115.600 ;
        RECT 279.200 115.200 279.600 115.600 ;
        RECT 279.800 115.200 280.200 115.600 ;
        RECT 280.400 115.200 280.800 115.600 ;
        RECT 315.200 115.200 315.600 115.600 ;
        RECT 315.800 115.200 316.200 115.600 ;
        RECT 316.400 115.200 316.800 115.600 ;
        RECT 135.200 21.400 135.600 21.800 ;
        RECT 135.800 21.400 136.200 21.800 ;
        RECT 136.400 21.400 136.800 21.800 ;
        RECT 171.200 21.400 171.600 21.800 ;
        RECT 171.800 21.400 172.200 21.800 ;
        RECT 172.400 21.400 172.800 21.800 ;
        RECT 207.200 21.400 207.600 21.800 ;
        RECT 207.800 21.400 208.200 21.800 ;
        RECT 208.400 21.400 208.800 21.800 ;
        RECT 243.200 21.400 243.600 21.800 ;
        RECT 243.800 21.400 244.200 21.800 ;
        RECT 244.400 21.400 244.800 21.800 ;
        RECT 279.200 21.400 279.600 21.800 ;
        RECT 279.800 21.400 280.200 21.800 ;
        RECT 280.400 21.400 280.800 21.800 ;
        RECT 315.200 21.400 315.600 21.800 ;
        RECT 315.800 21.400 316.200 21.800 ;
        RECT 316.400 21.400 316.800 21.800 ;
        RECT 135.200 20.800 135.600 21.200 ;
        RECT 135.800 20.800 136.200 21.200 ;
        RECT 136.400 20.800 136.800 21.200 ;
        RECT 171.200 20.800 171.600 21.200 ;
        RECT 171.800 20.800 172.200 21.200 ;
        RECT 172.400 20.800 172.800 21.200 ;
        RECT 207.200 20.800 207.600 21.200 ;
        RECT 207.800 20.800 208.200 21.200 ;
        RECT 208.400 20.800 208.800 21.200 ;
        RECT 243.200 20.800 243.600 21.200 ;
        RECT 243.800 20.800 244.200 21.200 ;
        RECT 244.400 20.800 244.800 21.200 ;
        RECT 279.200 20.800 279.600 21.200 ;
        RECT 279.800 20.800 280.200 21.200 ;
        RECT 280.400 20.800 280.800 21.200 ;
        RECT 315.200 20.800 315.600 21.200 ;
        RECT 315.800 20.800 316.200 21.200 ;
        RECT 316.400 20.800 316.800 21.200 ;
        RECT 135.200 20.200 135.600 20.600 ;
        RECT 135.800 20.200 136.200 20.600 ;
        RECT 136.400 20.200 136.800 20.600 ;
        RECT 171.200 20.200 171.600 20.600 ;
        RECT 171.800 20.200 172.200 20.600 ;
        RECT 172.400 20.200 172.800 20.600 ;
        RECT 207.200 20.200 207.600 20.600 ;
        RECT 207.800 20.200 208.200 20.600 ;
        RECT 208.400 20.200 208.800 20.600 ;
        RECT 243.200 20.200 243.600 20.600 ;
        RECT 243.800 20.200 244.200 20.600 ;
        RECT 244.400 20.200 244.800 20.600 ;
        RECT 279.200 20.200 279.600 20.600 ;
        RECT 279.800 20.200 280.200 20.600 ;
        RECT 280.400 20.200 280.800 20.600 ;
        RECT 315.200 20.200 315.600 20.600 ;
        RECT 315.800 20.200 316.200 20.600 ;
        RECT 316.400 20.200 316.800 20.600 ;
        RECT 140.200 17.400 140.600 17.800 ;
        RECT 140.800 17.400 141.200 17.800 ;
        RECT 141.400 17.400 141.800 17.800 ;
        RECT 153.200 17.400 153.600 17.800 ;
        RECT 153.800 17.400 154.200 17.800 ;
        RECT 154.400 17.400 154.800 17.800 ;
        RECT 189.200 17.400 189.600 17.800 ;
        RECT 189.800 17.400 190.200 17.800 ;
        RECT 190.400 17.400 190.800 17.800 ;
        RECT 225.200 17.400 225.600 17.800 ;
        RECT 225.800 17.400 226.200 17.800 ;
        RECT 226.400 17.400 226.800 17.800 ;
        RECT 261.200 17.400 261.600 17.800 ;
        RECT 261.800 17.400 262.200 17.800 ;
        RECT 262.400 17.400 262.800 17.800 ;
        RECT 297.200 17.400 297.600 17.800 ;
        RECT 297.800 17.400 298.200 17.800 ;
        RECT 298.400 17.400 298.800 17.800 ;
        RECT 310.200 17.400 310.600 17.800 ;
        RECT 310.800 17.400 311.200 17.800 ;
        RECT 311.400 17.400 311.800 17.800 ;
        RECT 140.200 16.800 140.600 17.200 ;
        RECT 140.800 16.800 141.200 17.200 ;
        RECT 141.400 16.800 141.800 17.200 ;
        RECT 153.200 16.800 153.600 17.200 ;
        RECT 153.800 16.800 154.200 17.200 ;
        RECT 154.400 16.800 154.800 17.200 ;
        RECT 189.200 16.800 189.600 17.200 ;
        RECT 189.800 16.800 190.200 17.200 ;
        RECT 190.400 16.800 190.800 17.200 ;
        RECT 225.200 16.800 225.600 17.200 ;
        RECT 225.800 16.800 226.200 17.200 ;
        RECT 226.400 16.800 226.800 17.200 ;
        RECT 261.200 16.800 261.600 17.200 ;
        RECT 261.800 16.800 262.200 17.200 ;
        RECT 262.400 16.800 262.800 17.200 ;
        RECT 297.200 16.800 297.600 17.200 ;
        RECT 297.800 16.800 298.200 17.200 ;
        RECT 298.400 16.800 298.800 17.200 ;
        RECT 310.200 16.800 310.600 17.200 ;
        RECT 310.800 16.800 311.200 17.200 ;
        RECT 311.400 16.800 311.800 17.200 ;
        RECT 140.200 16.200 140.600 16.600 ;
        RECT 140.800 16.200 141.200 16.600 ;
        RECT 141.400 16.200 141.800 16.600 ;
        RECT 153.200 16.200 153.600 16.600 ;
        RECT 153.800 16.200 154.200 16.600 ;
        RECT 154.400 16.200 154.800 16.600 ;
        RECT 189.200 16.200 189.600 16.600 ;
        RECT 189.800 16.200 190.200 16.600 ;
        RECT 190.400 16.200 190.800 16.600 ;
        RECT 225.200 16.200 225.600 16.600 ;
        RECT 225.800 16.200 226.200 16.600 ;
        RECT 226.400 16.200 226.800 16.600 ;
        RECT 261.200 16.200 261.600 16.600 ;
        RECT 261.800 16.200 262.200 16.600 ;
        RECT 262.400 16.200 262.800 16.600 ;
        RECT 297.200 16.200 297.600 16.600 ;
        RECT 297.800 16.200 298.200 16.600 ;
        RECT 298.400 16.200 298.800 16.600 ;
        RECT 310.200 16.200 310.600 16.600 ;
        RECT 310.800 16.200 311.200 16.600 ;
        RECT 311.400 16.200 311.800 16.600 ;
      LAYER met4 ;
        RECT 135.000 20.000 137.000 117.000 ;
        RECT 140.000 16.000 142.000 121.000 ;
        RECT 153.000 16.000 155.000 121.000 ;
        RECT 171.000 20.000 173.000 117.000 ;
        RECT 189.000 16.000 191.000 121.000 ;
        RECT 207.000 20.000 209.000 117.000 ;
        RECT 225.000 16.000 227.000 121.000 ;
        RECT 243.000 20.000 245.000 117.000 ;
        RECT 261.000 16.000 263.000 121.000 ;
        RECT 279.000 20.000 281.000 117.000 ;
        RECT 297.000 16.000 299.000 121.000 ;
        RECT 310.000 16.000 312.000 121.000 ;
        RECT 315.000 20.000 317.000 117.000 ;
  END
END power_ring_2_2
MACRO vco_r100
  CLASS BLOCK ;
  FOREIGN vco_r100 ;
  ORIGIN 0.000 1.000 ;
  SIZE 184.000 BY 105.000 ;
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 133.300 42.180 134.500 42.760 ;
        RECT 132.500 42.060 134.500 42.180 ;
        RECT 151.270 42.120 152.450 42.400 ;
        RECT 132.500 41.460 136.500 42.060 ;
        RECT 150.770 41.520 152.450 42.120 ;
        RECT 151.270 41.320 152.450 41.520 ;
        RECT 154.935 41.030 155.435 42.180 ;
        RECT 157.450 41.030 157.745 45.295 ;
        RECT 164.600 42.760 164.890 48.090 ;
        RECT 168.780 42.760 169.070 48.090 ;
        RECT 164.600 42.470 169.070 42.760 ;
        RECT 167.030 41.030 167.530 42.470 ;
        RECT 154.935 40.530 167.530 41.030 ;
        RECT 157.455 32.850 157.750 40.530 ;
        RECT 164.600 35.530 164.890 40.530 ;
      LAYER mcon ;
        RECT 132.560 41.520 133.200 42.150 ;
        RECT 133.400 41.460 134.100 42.150 ;
        RECT 134.300 41.460 134.900 42.060 ;
        RECT 135.100 41.460 135.700 42.060 ;
        RECT 135.900 41.460 136.500 42.060 ;
        RECT 150.820 41.570 151.220 42.070 ;
        RECT 151.420 41.570 152.370 42.070 ;
        RECT 154.935 41.520 155.435 42.120 ;
      LAYER met1 ;
        RECT 132.500 42.120 136.600 42.180 ;
        RECT 154.905 42.120 155.465 42.180 ;
        RECT 132.500 41.520 155.465 42.120 ;
        RECT 132.500 41.460 136.600 41.520 ;
        RECT 154.905 41.460 155.465 41.520 ;
        RECT 133.300 41.430 136.600 41.460 ;
      LAYER via ;
        RECT 149.010 41.530 149.590 42.110 ;
        RECT 149.750 41.530 150.330 42.110 ;
      LAYER met2 ;
        RECT 149.000 41.490 150.340 42.170 ;
        RECT 149.270 31.010 150.070 41.490 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 103.800 42.180 105.000 42.760 ;
        RECT 103.000 42.060 105.000 42.180 ;
        RECT 121.770 42.120 122.950 42.400 ;
        RECT 103.000 41.460 107.000 42.060 ;
        RECT 121.270 41.520 122.950 42.120 ;
        RECT 121.770 41.320 122.950 41.520 ;
        RECT 125.435 41.030 125.935 42.180 ;
        RECT 127.950 41.030 128.245 45.295 ;
        RECT 135.100 42.760 135.390 48.090 ;
        RECT 139.280 42.760 139.570 48.090 ;
        RECT 135.100 42.470 139.570 42.760 ;
        RECT 137.530 41.030 138.030 42.470 ;
        RECT 125.435 40.530 138.030 41.030 ;
        RECT 127.955 32.850 128.250 40.530 ;
        RECT 135.100 35.530 135.390 40.530 ;
      LAYER mcon ;
        RECT 103.060 41.520 103.700 42.150 ;
        RECT 103.900 41.460 104.600 42.150 ;
        RECT 104.800 41.460 105.400 42.060 ;
        RECT 105.600 41.460 106.200 42.060 ;
        RECT 106.400 41.460 107.000 42.060 ;
        RECT 121.320 41.570 121.720 42.070 ;
        RECT 121.920 41.570 122.870 42.070 ;
        RECT 125.435 41.520 125.935 42.120 ;
      LAYER met1 ;
        RECT 103.000 42.120 107.100 42.180 ;
        RECT 125.405 42.120 125.965 42.180 ;
        RECT 103.000 41.520 125.965 42.120 ;
        RECT 103.000 41.460 107.100 41.520 ;
        RECT 125.405 41.460 125.965 41.520 ;
        RECT 103.800 41.430 107.100 41.460 ;
      LAYER via ;
        RECT 119.510 41.530 120.090 42.110 ;
        RECT 120.250 41.530 120.830 42.110 ;
      LAYER met2 ;
        RECT 119.500 41.490 120.840 42.170 ;
        RECT 119.770 31.010 120.570 41.490 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 74.300 42.180 75.500 42.760 ;
        RECT 73.500 42.060 75.500 42.180 ;
        RECT 92.270 42.120 93.450 42.400 ;
        RECT 73.500 41.460 77.500 42.060 ;
        RECT 91.770 41.520 93.450 42.120 ;
        RECT 92.270 41.320 93.450 41.520 ;
        RECT 95.935 41.030 96.435 42.180 ;
        RECT 98.450 41.030 98.745 45.295 ;
        RECT 105.600 42.760 105.890 48.090 ;
        RECT 109.780 42.760 110.070 48.090 ;
        RECT 105.600 42.470 110.070 42.760 ;
        RECT 108.030 41.030 108.530 42.470 ;
        RECT 95.935 40.530 108.530 41.030 ;
        RECT 98.455 32.850 98.750 40.530 ;
        RECT 105.600 35.530 105.890 40.530 ;
      LAYER mcon ;
        RECT 73.560 41.520 74.200 42.150 ;
        RECT 74.400 41.460 75.100 42.150 ;
        RECT 75.300 41.460 75.900 42.060 ;
        RECT 76.100 41.460 76.700 42.060 ;
        RECT 76.900 41.460 77.500 42.060 ;
        RECT 91.820 41.570 92.220 42.070 ;
        RECT 92.420 41.570 93.370 42.070 ;
        RECT 95.935 41.520 96.435 42.120 ;
      LAYER met1 ;
        RECT 73.500 42.120 77.600 42.180 ;
        RECT 95.905 42.120 96.465 42.180 ;
        RECT 73.500 41.520 96.465 42.120 ;
        RECT 73.500 41.460 77.600 41.520 ;
        RECT 95.905 41.460 96.465 41.520 ;
        RECT 74.300 41.430 77.600 41.460 ;
      LAYER via ;
        RECT 90.010 41.530 90.590 42.110 ;
        RECT 90.750 41.530 91.330 42.110 ;
      LAYER met2 ;
        RECT 90.000 41.490 91.340 42.170 ;
        RECT 90.270 31.010 91.070 41.490 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 44.800 42.180 46.000 42.760 ;
        RECT 44.000 42.060 46.000 42.180 ;
        RECT 62.770 42.120 63.950 42.400 ;
        RECT 44.000 41.460 48.000 42.060 ;
        RECT 62.270 41.520 63.950 42.120 ;
        RECT 62.770 41.320 63.950 41.520 ;
        RECT 66.435 41.030 66.935 42.180 ;
        RECT 68.950 41.030 69.245 45.295 ;
        RECT 76.100 42.760 76.390 48.090 ;
        RECT 80.280 42.760 80.570 48.090 ;
        RECT 76.100 42.470 80.570 42.760 ;
        RECT 78.530 41.030 79.030 42.470 ;
        RECT 66.435 40.530 79.030 41.030 ;
        RECT 68.955 32.850 69.250 40.530 ;
        RECT 76.100 35.530 76.390 40.530 ;
      LAYER mcon ;
        RECT 44.060 41.520 44.700 42.150 ;
        RECT 44.900 41.460 45.600 42.150 ;
        RECT 45.800 41.460 46.400 42.060 ;
        RECT 46.600 41.460 47.200 42.060 ;
        RECT 47.400 41.460 48.000 42.060 ;
        RECT 62.320 41.570 62.720 42.070 ;
        RECT 62.920 41.570 63.870 42.070 ;
        RECT 66.435 41.520 66.935 42.120 ;
      LAYER met1 ;
        RECT 44.000 42.120 48.100 42.180 ;
        RECT 66.405 42.120 66.965 42.180 ;
        RECT 44.000 41.520 66.965 42.120 ;
        RECT 44.000 41.460 48.100 41.520 ;
        RECT 66.405 41.460 66.965 41.520 ;
        RECT 44.800 41.430 48.100 41.460 ;
      LAYER via ;
        RECT 60.510 41.530 61.090 42.110 ;
        RECT 61.250 41.530 61.830 42.110 ;
      LAYER met2 ;
        RECT 60.500 41.490 61.840 42.170 ;
        RECT 60.770 31.010 61.570 41.490 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 15.300 42.180 16.500 42.760 ;
        RECT 14.500 42.060 16.500 42.180 ;
        RECT 33.270 42.120 34.450 42.400 ;
        RECT 14.500 41.460 18.500 42.060 ;
        RECT 32.770 41.520 34.450 42.120 ;
        RECT 33.270 41.320 34.450 41.520 ;
        RECT 36.935 41.030 37.435 42.180 ;
        RECT 39.450 41.030 39.745 45.295 ;
        RECT 46.600 42.760 46.890 48.090 ;
        RECT 50.780 42.760 51.070 48.090 ;
        RECT 46.600 42.470 51.070 42.760 ;
        RECT 49.030 41.030 49.530 42.470 ;
        RECT 36.935 40.530 49.530 41.030 ;
        RECT 39.455 32.850 39.750 40.530 ;
        RECT 46.600 35.530 46.890 40.530 ;
      LAYER mcon ;
        RECT 14.560 41.520 15.200 42.150 ;
        RECT 15.400 41.460 16.100 42.150 ;
        RECT 16.300 41.460 16.900 42.060 ;
        RECT 17.100 41.460 17.700 42.060 ;
        RECT 17.900 41.460 18.500 42.060 ;
        RECT 32.820 41.570 33.220 42.070 ;
        RECT 33.420 41.570 34.370 42.070 ;
        RECT 36.935 41.520 37.435 42.120 ;
      LAYER met1 ;
        RECT 14.500 42.120 18.600 42.180 ;
        RECT 36.905 42.120 37.465 42.180 ;
        RECT 14.500 41.520 37.465 42.120 ;
        RECT 14.500 41.460 18.600 41.520 ;
        RECT 36.905 41.460 37.465 41.520 ;
        RECT 15.300 41.430 18.600 41.460 ;
      LAYER via ;
        RECT 31.010 41.530 31.590 42.110 ;
        RECT 31.750 41.530 32.330 42.110 ;
      LAYER met2 ;
        RECT 31.000 41.490 32.340 42.170 ;
        RECT 31.270 31.010 32.070 41.490 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.680500 ;
    PORT
      LAYER li1 ;
        RECT 5.440 61.625 6.035 61.965 ;
        RECT 5.440 60.305 5.615 61.625 ;
        RECT 5.440 60.175 6.035 60.305 ;
        RECT 6.860 60.175 7.160 61.010 ;
        RECT 30.890 60.620 34.890 61.220 ;
        RECT 5.440 59.875 7.160 60.175 ;
        RECT 32.890 60.500 34.890 60.620 ;
        RECT 32.890 59.920 34.090 60.500 ;
        RECT 5.440 59.755 6.035 59.875 ;
        RECT 3.770 42.120 4.950 42.400 ;
        RECT 3.270 41.520 4.950 42.120 ;
        RECT 3.770 41.320 4.950 41.520 ;
        RECT 7.435 41.030 7.935 42.180 ;
        RECT 9.950 41.030 10.245 45.295 ;
        RECT 17.100 42.760 17.390 48.090 ;
        RECT 21.280 42.760 21.570 48.090 ;
        RECT 17.100 42.470 21.570 42.760 ;
        RECT 19.530 41.030 20.030 42.470 ;
        RECT 7.435 40.530 20.030 41.030 ;
        RECT 9.955 32.850 10.250 40.530 ;
        RECT 17.100 35.530 17.390 40.530 ;
      LAYER mcon ;
        RECT 6.925 60.775 7.095 60.945 ;
        RECT 30.890 60.620 31.490 61.220 ;
        RECT 31.690 60.620 32.290 61.220 ;
        RECT 32.490 60.620 33.090 61.220 ;
        RECT 33.290 60.530 33.990 61.220 ;
        RECT 34.190 60.530 34.830 61.160 ;
        RECT 3.320 41.570 3.720 42.070 ;
        RECT 3.920 41.570 4.870 42.070 ;
        RECT 7.435 41.520 7.935 42.120 ;
      LAYER met1 ;
        RECT 30.790 61.220 34.090 61.250 ;
        RECT 30.790 61.160 34.890 61.220 ;
        RECT 6.800 61.010 7.220 61.040 ;
        RECT 17.000 61.010 34.890 61.160 ;
        RECT 6.800 60.710 34.890 61.010 ;
        RECT 6.800 60.680 7.220 60.710 ;
        RECT 17.000 60.560 34.890 60.710 ;
        RECT 30.790 60.500 34.890 60.560 ;
        RECT 7.405 42.120 7.965 42.180 ;
        RECT 2.000 41.520 7.965 42.120 ;
        RECT 7.405 41.460 7.965 41.520 ;
      LAYER via ;
        RECT 17.925 60.570 18.825 61.150 ;
        RECT 6.765 41.530 7.345 42.110 ;
      LAYER met2 ;
        RECT 17.120 60.510 18.865 61.210 ;
        RECT 17.120 49.650 17.820 60.510 ;
        RECT 6.705 48.950 17.820 49.650 ;
        RECT 6.705 41.470 7.405 48.950 ;
        RECT 13.270 31.010 14.070 48.950 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 32.000 62.150 32.290 67.150 ;
        RECT 39.140 62.150 39.435 69.830 ;
        RECT 29.360 61.650 41.955 62.150 ;
        RECT 29.360 60.210 29.860 61.650 ;
        RECT 27.820 59.920 32.290 60.210 ;
        RECT 27.820 54.590 28.110 59.920 ;
        RECT 32.000 54.590 32.290 59.920 ;
        RECT 39.145 57.385 39.440 61.650 ;
        RECT 41.455 60.500 41.955 61.650 ;
        RECT 44.440 61.160 45.620 61.360 ;
        RECT 44.440 60.560 46.120 61.160 ;
        RECT 60.390 60.620 64.390 61.220 ;
        RECT 44.440 60.280 45.620 60.560 ;
        RECT 62.390 60.500 64.390 60.620 ;
        RECT 62.390 59.920 63.590 60.500 ;
      LAYER mcon ;
        RECT 41.455 60.560 41.955 61.160 ;
        RECT 44.520 60.610 45.470 61.110 ;
        RECT 45.670 60.610 46.070 61.110 ;
        RECT 60.390 60.620 60.990 61.220 ;
        RECT 61.190 60.620 61.790 61.220 ;
        RECT 61.990 60.620 62.590 61.220 ;
        RECT 62.790 60.530 63.490 61.220 ;
        RECT 63.690 60.530 64.330 61.160 ;
      LAYER met1 ;
        RECT 60.290 61.220 63.590 61.250 ;
        RECT 41.425 61.160 41.985 61.220 ;
        RECT 60.290 61.160 64.390 61.220 ;
        RECT 41.425 60.560 64.390 61.160 ;
        RECT 41.425 60.500 41.985 60.560 ;
        RECT 60.290 60.500 64.390 60.560 ;
      LAYER via ;
        RECT 46.560 60.570 47.140 61.150 ;
        RECT 47.300 60.570 47.880 61.150 ;
      LAYER met2 ;
        RECT 46.820 61.220 47.620 71.670 ;
        RECT 46.550 60.510 47.890 61.220 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 61.500 62.150 61.790 67.150 ;
        RECT 68.640 62.150 68.935 69.830 ;
        RECT 58.860 61.650 71.455 62.150 ;
        RECT 58.860 60.210 59.360 61.650 ;
        RECT 57.320 59.920 61.790 60.210 ;
        RECT 57.320 54.590 57.610 59.920 ;
        RECT 61.500 54.590 61.790 59.920 ;
        RECT 68.645 57.385 68.940 61.650 ;
        RECT 70.955 60.500 71.455 61.650 ;
        RECT 73.940 61.160 75.120 61.360 ;
        RECT 73.940 60.560 75.620 61.160 ;
        RECT 89.890 60.620 93.890 61.220 ;
        RECT 73.940 60.280 75.120 60.560 ;
        RECT 91.890 60.500 93.890 60.620 ;
        RECT 91.890 59.920 93.090 60.500 ;
      LAYER mcon ;
        RECT 70.955 60.560 71.455 61.160 ;
        RECT 74.020 60.610 74.970 61.110 ;
        RECT 75.170 60.610 75.570 61.110 ;
        RECT 89.890 60.620 90.490 61.220 ;
        RECT 90.690 60.620 91.290 61.220 ;
        RECT 91.490 60.620 92.090 61.220 ;
        RECT 92.290 60.530 92.990 61.220 ;
        RECT 93.190 60.530 93.830 61.160 ;
      LAYER met1 ;
        RECT 89.790 61.220 93.090 61.250 ;
        RECT 70.925 61.160 71.485 61.220 ;
        RECT 89.790 61.160 93.890 61.220 ;
        RECT 70.925 60.560 93.890 61.160 ;
        RECT 70.925 60.500 71.485 60.560 ;
        RECT 89.790 60.500 93.890 60.560 ;
      LAYER via ;
        RECT 76.060 60.570 76.640 61.150 ;
        RECT 76.800 60.570 77.380 61.150 ;
      LAYER met2 ;
        RECT 76.320 61.220 77.120 71.670 ;
        RECT 76.050 60.510 77.390 61.220 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 91.000 62.150 91.290 67.150 ;
        RECT 98.140 62.150 98.435 69.830 ;
        RECT 88.360 61.650 100.955 62.150 ;
        RECT 88.360 60.210 88.860 61.650 ;
        RECT 86.820 59.920 91.290 60.210 ;
        RECT 86.820 54.590 87.110 59.920 ;
        RECT 91.000 54.590 91.290 59.920 ;
        RECT 98.145 57.385 98.440 61.650 ;
        RECT 100.455 60.500 100.955 61.650 ;
        RECT 103.440 61.160 104.620 61.360 ;
        RECT 103.440 60.560 105.120 61.160 ;
        RECT 119.390 60.620 123.390 61.220 ;
        RECT 103.440 60.280 104.620 60.560 ;
        RECT 121.390 60.500 123.390 60.620 ;
        RECT 121.390 59.920 122.590 60.500 ;
      LAYER mcon ;
        RECT 100.455 60.560 100.955 61.160 ;
        RECT 103.520 60.610 104.470 61.110 ;
        RECT 104.670 60.610 105.070 61.110 ;
        RECT 119.390 60.620 119.990 61.220 ;
        RECT 120.190 60.620 120.790 61.220 ;
        RECT 120.990 60.620 121.590 61.220 ;
        RECT 121.790 60.530 122.490 61.220 ;
        RECT 122.690 60.530 123.330 61.160 ;
      LAYER met1 ;
        RECT 119.290 61.220 122.590 61.250 ;
        RECT 100.425 61.160 100.985 61.220 ;
        RECT 119.290 61.160 123.390 61.220 ;
        RECT 100.425 60.560 123.390 61.160 ;
        RECT 100.425 60.500 100.985 60.560 ;
        RECT 119.290 60.500 123.390 60.560 ;
      LAYER via ;
        RECT 105.560 60.570 106.140 61.150 ;
        RECT 106.300 60.570 106.880 61.150 ;
      LAYER met2 ;
        RECT 105.820 61.220 106.620 71.670 ;
        RECT 105.550 60.510 106.890 61.220 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 120.500 62.150 120.790 67.150 ;
        RECT 127.640 62.150 127.935 69.830 ;
        RECT 117.860 61.650 130.455 62.150 ;
        RECT 117.860 60.210 118.360 61.650 ;
        RECT 116.320 59.920 120.790 60.210 ;
        RECT 116.320 54.590 116.610 59.920 ;
        RECT 120.500 54.590 120.790 59.920 ;
        RECT 127.645 57.385 127.940 61.650 ;
        RECT 129.955 60.500 130.455 61.650 ;
        RECT 132.940 61.160 134.120 61.360 ;
        RECT 132.940 60.560 134.620 61.160 ;
        RECT 148.890 60.620 152.890 61.220 ;
        RECT 132.940 60.280 134.120 60.560 ;
        RECT 150.890 60.500 152.890 60.620 ;
        RECT 150.890 59.920 152.090 60.500 ;
      LAYER mcon ;
        RECT 129.955 60.560 130.455 61.160 ;
        RECT 133.020 60.610 133.970 61.110 ;
        RECT 134.170 60.610 134.570 61.110 ;
        RECT 148.890 60.620 149.490 61.220 ;
        RECT 149.690 60.620 150.290 61.220 ;
        RECT 150.490 60.620 151.090 61.220 ;
        RECT 151.290 60.530 151.990 61.220 ;
        RECT 152.190 60.530 152.830 61.160 ;
      LAYER met1 ;
        RECT 148.790 61.220 152.090 61.250 ;
        RECT 129.925 61.160 130.485 61.220 ;
        RECT 148.790 61.160 152.890 61.220 ;
        RECT 129.925 60.560 152.890 61.160 ;
        RECT 129.925 60.500 130.485 60.560 ;
        RECT 148.790 60.500 152.890 60.560 ;
      LAYER via ;
        RECT 135.060 60.570 135.640 61.150 ;
        RECT 135.800 60.570 136.380 61.150 ;
      LAYER met2 ;
        RECT 135.320 61.220 136.120 71.670 ;
        RECT 135.050 60.510 136.390 61.220 ;
    END
  END p[9]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 150.000 62.150 150.290 67.150 ;
        RECT 157.140 62.150 157.435 69.830 ;
        RECT 147.360 61.650 159.955 62.150 ;
        RECT 147.360 60.210 147.860 61.650 ;
        RECT 145.820 59.920 150.290 60.210 ;
        RECT 145.820 54.590 146.110 59.920 ;
        RECT 150.000 54.590 150.290 59.920 ;
        RECT 157.145 57.385 157.440 61.650 ;
        RECT 159.455 60.500 159.955 61.650 ;
        RECT 162.440 61.160 163.620 61.360 ;
        RECT 162.440 60.560 164.120 61.160 ;
        RECT 162.440 60.280 163.620 60.560 ;
        RECT 162.800 42.180 164.000 42.760 ;
        RECT 162.000 42.060 164.000 42.180 ;
        RECT 162.000 41.460 166.000 42.060 ;
      LAYER mcon ;
        RECT 159.455 60.560 159.955 61.160 ;
        RECT 162.520 60.610 163.470 61.110 ;
        RECT 163.670 60.610 164.070 61.110 ;
        RECT 162.060 41.520 162.700 42.150 ;
        RECT 162.900 41.460 163.600 42.150 ;
        RECT 163.800 41.460 164.400 42.060 ;
        RECT 164.600 41.460 165.200 42.060 ;
        RECT 165.400 41.460 166.000 42.060 ;
      LAYER met1 ;
        RECT 159.425 61.160 159.985 61.220 ;
        RECT 159.425 60.560 165.440 61.160 ;
        RECT 159.425 60.500 159.985 60.560 ;
        RECT 162.000 42.120 166.100 42.180 ;
        RECT 162.000 41.520 179.000 42.120 ;
        RECT 162.000 41.460 166.100 41.520 ;
        RECT 162.800 41.430 166.100 41.460 ;
      LAYER via ;
        RECT 164.470 60.570 165.370 61.150 ;
        RECT 166.150 41.530 166.730 42.110 ;
        RECT 166.870 41.530 167.450 42.110 ;
      LAYER met2 ;
        RECT 164.450 60.510 166.790 61.210 ;
        RECT 166.090 42.170 166.790 60.510 ;
        RECT 166.090 41.440 167.460 42.170 ;
        RECT 166.360 31.010 167.160 41.440 ;
    END
  END p[10]
  PIN input_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 175.550 58.040 177.550 58.210 ;
        RECT 175.630 58.010 177.470 58.040 ;
      LAYER mcon ;
        RECT 175.745 58.025 175.915 58.195 ;
        RECT 176.105 58.025 176.275 58.195 ;
        RECT 176.465 58.025 176.635 58.195 ;
        RECT 176.825 58.025 176.995 58.195 ;
        RECT 177.185 58.025 177.355 58.195 ;
      LAYER met1 ;
        RECT 175.520 57.980 177.580 58.240 ;
      LAYER via ;
        RECT 175.620 57.980 175.880 58.240 ;
        RECT 175.940 57.980 176.200 58.240 ;
        RECT 176.260 57.980 176.520 58.240 ;
        RECT 176.580 57.980 176.840 58.240 ;
        RECT 176.900 57.980 177.160 58.240 ;
        RECT 177.220 57.980 177.480 58.240 ;
      LAYER met2 ;
        RECT 175.570 57.690 184.000 58.490 ;
      LAYER via2 ;
        RECT 183.000 57.890 183.400 58.290 ;
        RECT 183.530 57.890 183.930 58.290 ;
      LAYER met3 ;
        RECT 182.970 57.690 184.000 58.490 ;
    END
  END input_analog
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 3.630 60.805 6.310 62.640 ;
        RECT 7.800 60.805 9.560 62.640 ;
        RECT 18.390 56.545 24.240 62.420 ;
        RECT 29.220 62.080 35.070 67.935 ;
        RECT 42.840 62.610 46.600 67.885 ;
        RECT 36.365 56.550 40.125 61.860 ;
        RECT 47.890 56.545 53.740 62.420 ;
        RECT 58.720 62.080 64.570 67.935 ;
        RECT 72.340 62.610 76.100 67.885 ;
        RECT 65.865 56.550 69.625 61.860 ;
        RECT 77.390 56.545 83.240 62.420 ;
        RECT 88.220 62.080 94.070 67.935 ;
        RECT 101.840 62.610 105.600 67.885 ;
        RECT 95.365 56.550 99.125 61.860 ;
        RECT 106.890 56.545 112.740 62.420 ;
        RECT 117.720 62.080 123.570 67.935 ;
        RECT 131.340 62.610 135.100 67.885 ;
        RECT 124.865 56.550 128.625 61.860 ;
        RECT 136.390 56.545 142.240 62.420 ;
        RECT 147.220 62.080 153.070 67.935 ;
        RECT 160.840 62.610 164.600 67.885 ;
        RECT 154.365 56.550 158.125 61.860 ;
        RECT 9.265 40.820 13.025 46.130 ;
        RECT 2.790 34.795 6.550 40.070 ;
        RECT 14.320 34.745 20.170 40.600 ;
        RECT 25.150 40.260 31.000 46.135 ;
        RECT 38.765 40.820 42.525 46.130 ;
        RECT 32.290 34.795 36.050 40.070 ;
        RECT 43.820 34.745 49.670 40.600 ;
        RECT 54.650 40.260 60.500 46.135 ;
        RECT 68.265 40.820 72.025 46.130 ;
        RECT 61.790 34.795 65.550 40.070 ;
        RECT 73.320 34.745 79.170 40.600 ;
        RECT 84.150 40.260 90.000 46.135 ;
        RECT 97.765 40.820 101.525 46.130 ;
        RECT 91.290 34.795 95.050 40.070 ;
        RECT 102.820 34.745 108.670 40.600 ;
        RECT 113.650 40.260 119.500 46.135 ;
        RECT 127.265 40.820 131.025 46.130 ;
        RECT 120.790 34.795 124.550 40.070 ;
        RECT 132.320 34.745 138.170 40.600 ;
        RECT 143.150 40.260 149.000 46.135 ;
        RECT 156.765 40.820 160.525 46.130 ;
        RECT 150.290 34.795 154.050 40.070 ;
        RECT 161.820 34.745 167.670 40.600 ;
        RECT 172.650 40.260 178.500 46.135 ;
      LAYER li1 ;
        RECT 29.400 67.755 31.745 67.900 ;
        RECT 32.545 67.755 34.890 67.900 ;
        RECT 44.325 67.870 46.420 67.900 ;
        RECT 29.400 67.585 34.890 67.755 ;
        RECT 44.170 67.705 46.420 67.870 ;
        RECT 29.400 67.420 31.745 67.585 ;
        RECT 32.545 67.420 34.890 67.585 ;
        RECT 29.400 62.760 29.570 67.420 ;
        RECT 29.910 62.590 30.200 67.420 ;
        RECT 34.090 62.590 34.380 67.420 ;
        RECT 34.720 62.820 34.890 67.420 ;
        RECT 43.020 67.535 46.420 67.705 ;
        RECT 43.020 64.560 43.190 67.535 ;
        RECT 44.170 67.450 46.420 67.535 ;
        RECT 44.325 67.420 46.420 67.450 ;
        RECT 45.620 63.010 45.910 67.420 ;
        RECT 46.250 63.005 46.420 67.420 ;
        RECT 58.900 67.755 61.245 67.900 ;
        RECT 62.045 67.755 64.390 67.900 ;
        RECT 73.825 67.870 75.920 67.900 ;
        RECT 58.900 67.585 64.390 67.755 ;
        RECT 73.670 67.705 75.920 67.870 ;
        RECT 58.900 67.420 61.245 67.585 ;
        RECT 62.045 67.420 64.390 67.585 ;
        RECT 58.900 62.760 59.070 67.420 ;
        RECT 59.410 62.590 59.700 67.420 ;
        RECT 63.590 62.590 63.880 67.420 ;
        RECT 64.220 62.820 64.390 67.420 ;
        RECT 72.520 67.535 75.920 67.705 ;
        RECT 72.520 64.560 72.690 67.535 ;
        RECT 73.670 67.450 75.920 67.535 ;
        RECT 73.825 67.420 75.920 67.450 ;
        RECT 75.120 63.010 75.410 67.420 ;
        RECT 75.750 63.005 75.920 67.420 ;
        RECT 88.400 67.755 90.745 67.900 ;
        RECT 91.545 67.755 93.890 67.900 ;
        RECT 103.325 67.870 105.420 67.900 ;
        RECT 88.400 67.585 93.890 67.755 ;
        RECT 103.170 67.705 105.420 67.870 ;
        RECT 88.400 67.420 90.745 67.585 ;
        RECT 91.545 67.420 93.890 67.585 ;
        RECT 88.400 62.760 88.570 67.420 ;
        RECT 88.910 62.590 89.200 67.420 ;
        RECT 93.090 62.590 93.380 67.420 ;
        RECT 93.720 62.820 93.890 67.420 ;
        RECT 102.020 67.535 105.420 67.705 ;
        RECT 102.020 64.560 102.190 67.535 ;
        RECT 103.170 67.450 105.420 67.535 ;
        RECT 103.325 67.420 105.420 67.450 ;
        RECT 104.620 63.010 104.910 67.420 ;
        RECT 105.250 63.005 105.420 67.420 ;
        RECT 117.900 67.755 120.245 67.900 ;
        RECT 121.045 67.755 123.390 67.900 ;
        RECT 132.825 67.870 134.920 67.900 ;
        RECT 117.900 67.585 123.390 67.755 ;
        RECT 132.670 67.705 134.920 67.870 ;
        RECT 117.900 67.420 120.245 67.585 ;
        RECT 121.045 67.420 123.390 67.585 ;
        RECT 117.900 62.760 118.070 67.420 ;
        RECT 118.410 62.590 118.700 67.420 ;
        RECT 122.590 62.590 122.880 67.420 ;
        RECT 123.220 62.820 123.390 67.420 ;
        RECT 131.520 67.535 134.920 67.705 ;
        RECT 131.520 64.560 131.690 67.535 ;
        RECT 132.670 67.450 134.920 67.535 ;
        RECT 132.825 67.420 134.920 67.450 ;
        RECT 134.120 63.010 134.410 67.420 ;
        RECT 134.750 63.005 134.920 67.420 ;
        RECT 147.400 67.755 149.745 67.900 ;
        RECT 150.545 67.755 152.890 67.900 ;
        RECT 162.325 67.870 164.420 67.900 ;
        RECT 147.400 67.585 152.890 67.755 ;
        RECT 162.170 67.705 164.420 67.870 ;
        RECT 147.400 67.420 149.745 67.585 ;
        RECT 150.545 67.420 152.890 67.585 ;
        RECT 147.400 62.760 147.570 67.420 ;
        RECT 147.910 62.590 148.200 67.420 ;
        RECT 152.090 62.590 152.380 67.420 ;
        RECT 152.720 62.820 152.890 67.420 ;
        RECT 161.020 67.535 164.420 67.705 ;
        RECT 161.020 64.560 161.190 67.535 ;
        RECT 162.170 67.450 164.420 67.535 ;
        RECT 162.325 67.420 164.420 67.450 ;
        RECT 163.620 63.010 163.910 67.420 ;
        RECT 164.250 63.005 164.420 67.420 ;
        RECT 4.340 62.305 5.310 62.460 ;
        RECT 8.340 62.305 9.310 62.460 ;
        RECT 3.820 62.135 6.120 62.305 ;
        RECT 7.990 62.135 9.370 62.305 ;
        RECT 4.335 61.735 5.270 62.135 ;
        RECT 8.265 61.410 8.595 62.135 ;
        RECT 18.570 57.020 18.740 61.875 ;
        RECT 19.080 57.020 19.370 61.870 ;
        RECT 23.260 57.020 23.550 61.870 ;
        RECT 23.890 57.020 24.060 61.875 ;
        RECT 18.570 56.895 20.915 57.020 ;
        RECT 21.715 56.990 24.060 57.020 ;
        RECT 36.545 57.020 36.715 60.945 ;
        RECT 37.055 57.020 37.345 61.090 ;
        RECT 36.545 56.990 38.640 57.020 ;
        RECT 21.715 56.895 24.240 56.990 ;
        RECT 18.570 56.725 24.240 56.895 ;
        RECT 18.570 56.540 20.915 56.725 ;
        RECT 21.715 56.570 24.240 56.725 ;
        RECT 36.545 56.900 38.795 56.990 ;
        RECT 39.775 56.900 39.945 60.935 ;
        RECT 36.545 56.730 39.945 56.900 ;
        RECT 48.070 57.020 48.240 61.875 ;
        RECT 48.580 57.020 48.870 61.870 ;
        RECT 52.760 57.020 53.050 61.870 ;
        RECT 53.390 57.020 53.560 61.875 ;
        RECT 48.070 56.895 50.415 57.020 ;
        RECT 51.215 56.990 53.560 57.020 ;
        RECT 66.045 57.020 66.215 60.945 ;
        RECT 66.555 57.020 66.845 61.090 ;
        RECT 66.045 56.990 68.140 57.020 ;
        RECT 51.215 56.895 53.740 56.990 ;
        RECT 36.545 56.570 38.795 56.730 ;
        RECT 48.070 56.725 53.740 56.895 ;
        RECT 21.715 56.540 24.060 56.570 ;
        RECT 36.545 56.540 38.640 56.570 ;
        RECT 48.070 56.540 50.415 56.725 ;
        RECT 51.215 56.570 53.740 56.725 ;
        RECT 66.045 56.900 68.295 56.990 ;
        RECT 69.275 56.900 69.445 60.935 ;
        RECT 66.045 56.730 69.445 56.900 ;
        RECT 77.570 57.020 77.740 61.875 ;
        RECT 78.080 57.020 78.370 61.870 ;
        RECT 82.260 57.020 82.550 61.870 ;
        RECT 82.890 57.020 83.060 61.875 ;
        RECT 77.570 56.895 79.915 57.020 ;
        RECT 80.715 56.990 83.060 57.020 ;
        RECT 95.545 57.020 95.715 60.945 ;
        RECT 96.055 57.020 96.345 61.090 ;
        RECT 95.545 56.990 97.640 57.020 ;
        RECT 80.715 56.895 83.240 56.990 ;
        RECT 66.045 56.570 68.295 56.730 ;
        RECT 77.570 56.725 83.240 56.895 ;
        RECT 51.215 56.540 53.560 56.570 ;
        RECT 66.045 56.540 68.140 56.570 ;
        RECT 77.570 56.540 79.915 56.725 ;
        RECT 80.715 56.570 83.240 56.725 ;
        RECT 95.545 56.900 97.795 56.990 ;
        RECT 98.775 56.900 98.945 60.935 ;
        RECT 95.545 56.730 98.945 56.900 ;
        RECT 107.070 57.020 107.240 61.875 ;
        RECT 107.580 57.020 107.870 61.870 ;
        RECT 111.760 57.020 112.050 61.870 ;
        RECT 112.390 57.020 112.560 61.875 ;
        RECT 107.070 56.895 109.415 57.020 ;
        RECT 110.215 56.990 112.560 57.020 ;
        RECT 125.045 57.020 125.215 60.945 ;
        RECT 125.555 57.020 125.845 61.090 ;
        RECT 125.045 56.990 127.140 57.020 ;
        RECT 110.215 56.895 112.740 56.990 ;
        RECT 95.545 56.570 97.795 56.730 ;
        RECT 107.070 56.725 112.740 56.895 ;
        RECT 80.715 56.540 83.060 56.570 ;
        RECT 95.545 56.540 97.640 56.570 ;
        RECT 107.070 56.540 109.415 56.725 ;
        RECT 110.215 56.570 112.740 56.725 ;
        RECT 125.045 56.900 127.295 56.990 ;
        RECT 128.275 56.900 128.445 60.935 ;
        RECT 125.045 56.730 128.445 56.900 ;
        RECT 136.570 57.020 136.740 61.875 ;
        RECT 137.080 57.020 137.370 61.870 ;
        RECT 141.260 57.020 141.550 61.870 ;
        RECT 141.890 57.020 142.060 61.875 ;
        RECT 136.570 56.895 138.915 57.020 ;
        RECT 139.715 56.990 142.060 57.020 ;
        RECT 154.545 57.020 154.715 60.945 ;
        RECT 155.055 57.020 155.345 61.090 ;
        RECT 154.545 56.990 156.640 57.020 ;
        RECT 139.715 56.895 142.240 56.990 ;
        RECT 125.045 56.570 127.295 56.730 ;
        RECT 136.570 56.725 142.240 56.895 ;
        RECT 110.215 56.540 112.560 56.570 ;
        RECT 125.045 56.540 127.140 56.570 ;
        RECT 136.570 56.540 138.915 56.725 ;
        RECT 139.715 56.570 142.240 56.725 ;
        RECT 154.545 56.900 156.795 56.990 ;
        RECT 157.775 56.900 157.945 60.935 ;
        RECT 154.545 56.730 157.945 56.900 ;
        RECT 154.545 56.570 156.795 56.730 ;
        RECT 139.715 56.540 142.060 56.570 ;
        RECT 154.545 56.540 156.640 56.570 ;
        RECT 10.750 46.110 12.845 46.140 ;
        RECT 25.330 46.110 27.675 46.140 ;
        RECT 10.595 45.950 12.845 46.110 ;
        RECT 9.445 45.780 12.845 45.950 ;
        RECT 9.445 41.745 9.615 45.780 ;
        RECT 10.595 45.690 12.845 45.780 ;
        RECT 25.150 45.955 27.675 46.110 ;
        RECT 28.475 45.955 30.820 46.140 ;
        RECT 40.250 46.110 42.345 46.140 ;
        RECT 54.830 46.110 57.175 46.140 ;
        RECT 25.150 45.785 30.820 45.955 ;
        RECT 40.095 45.950 42.345 46.110 ;
        RECT 25.150 45.690 27.675 45.785 ;
        RECT 10.750 45.660 12.845 45.690 ;
        RECT 12.045 41.590 12.335 45.660 ;
        RECT 12.675 41.735 12.845 45.660 ;
        RECT 25.330 45.660 27.675 45.690 ;
        RECT 28.475 45.660 30.820 45.785 ;
        RECT 25.330 40.805 25.500 45.660 ;
        RECT 25.840 40.810 26.130 45.660 ;
        RECT 30.020 40.810 30.310 45.660 ;
        RECT 30.650 40.805 30.820 45.660 ;
        RECT 38.945 45.780 42.345 45.950 ;
        RECT 38.945 41.745 39.115 45.780 ;
        RECT 40.095 45.690 42.345 45.780 ;
        RECT 54.650 45.955 57.175 46.110 ;
        RECT 57.975 45.955 60.320 46.140 ;
        RECT 69.750 46.110 71.845 46.140 ;
        RECT 84.330 46.110 86.675 46.140 ;
        RECT 54.650 45.785 60.320 45.955 ;
        RECT 69.595 45.950 71.845 46.110 ;
        RECT 54.650 45.690 57.175 45.785 ;
        RECT 40.250 45.660 42.345 45.690 ;
        RECT 41.545 41.590 41.835 45.660 ;
        RECT 42.175 41.735 42.345 45.660 ;
        RECT 54.830 45.660 57.175 45.690 ;
        RECT 57.975 45.660 60.320 45.785 ;
        RECT 54.830 40.805 55.000 45.660 ;
        RECT 55.340 40.810 55.630 45.660 ;
        RECT 59.520 40.810 59.810 45.660 ;
        RECT 60.150 40.805 60.320 45.660 ;
        RECT 68.445 45.780 71.845 45.950 ;
        RECT 68.445 41.745 68.615 45.780 ;
        RECT 69.595 45.690 71.845 45.780 ;
        RECT 84.150 45.955 86.675 46.110 ;
        RECT 87.475 45.955 89.820 46.140 ;
        RECT 99.250 46.110 101.345 46.140 ;
        RECT 113.830 46.110 116.175 46.140 ;
        RECT 84.150 45.785 89.820 45.955 ;
        RECT 99.095 45.950 101.345 46.110 ;
        RECT 84.150 45.690 86.675 45.785 ;
        RECT 69.750 45.660 71.845 45.690 ;
        RECT 71.045 41.590 71.335 45.660 ;
        RECT 71.675 41.735 71.845 45.660 ;
        RECT 84.330 45.660 86.675 45.690 ;
        RECT 87.475 45.660 89.820 45.785 ;
        RECT 84.330 40.805 84.500 45.660 ;
        RECT 84.840 40.810 85.130 45.660 ;
        RECT 89.020 40.810 89.310 45.660 ;
        RECT 89.650 40.805 89.820 45.660 ;
        RECT 97.945 45.780 101.345 45.950 ;
        RECT 97.945 41.745 98.115 45.780 ;
        RECT 99.095 45.690 101.345 45.780 ;
        RECT 113.650 45.955 116.175 46.110 ;
        RECT 116.975 45.955 119.320 46.140 ;
        RECT 128.750 46.110 130.845 46.140 ;
        RECT 143.330 46.110 145.675 46.140 ;
        RECT 113.650 45.785 119.320 45.955 ;
        RECT 128.595 45.950 130.845 46.110 ;
        RECT 113.650 45.690 116.175 45.785 ;
        RECT 99.250 45.660 101.345 45.690 ;
        RECT 100.545 41.590 100.835 45.660 ;
        RECT 101.175 41.735 101.345 45.660 ;
        RECT 113.830 45.660 116.175 45.690 ;
        RECT 116.975 45.660 119.320 45.785 ;
        RECT 113.830 40.805 114.000 45.660 ;
        RECT 114.340 40.810 114.630 45.660 ;
        RECT 118.520 40.810 118.810 45.660 ;
        RECT 119.150 40.805 119.320 45.660 ;
        RECT 127.445 45.780 130.845 45.950 ;
        RECT 127.445 41.745 127.615 45.780 ;
        RECT 128.595 45.690 130.845 45.780 ;
        RECT 143.150 45.955 145.675 46.110 ;
        RECT 146.475 45.955 148.820 46.140 ;
        RECT 158.250 46.110 160.345 46.140 ;
        RECT 172.830 46.110 175.175 46.140 ;
        RECT 143.150 45.785 148.820 45.955 ;
        RECT 158.095 45.950 160.345 46.110 ;
        RECT 143.150 45.690 145.675 45.785 ;
        RECT 128.750 45.660 130.845 45.690 ;
        RECT 130.045 41.590 130.335 45.660 ;
        RECT 130.675 41.735 130.845 45.660 ;
        RECT 143.330 45.660 145.675 45.690 ;
        RECT 146.475 45.660 148.820 45.785 ;
        RECT 143.330 40.805 143.500 45.660 ;
        RECT 143.840 40.810 144.130 45.660 ;
        RECT 148.020 40.810 148.310 45.660 ;
        RECT 148.650 40.805 148.820 45.660 ;
        RECT 156.945 45.780 160.345 45.950 ;
        RECT 156.945 41.745 157.115 45.780 ;
        RECT 158.095 45.690 160.345 45.780 ;
        RECT 172.650 45.955 175.175 46.110 ;
        RECT 175.975 45.955 178.320 46.140 ;
        RECT 172.650 45.785 178.320 45.955 ;
        RECT 172.650 45.690 175.175 45.785 ;
        RECT 158.250 45.660 160.345 45.690 ;
        RECT 159.545 41.590 159.835 45.660 ;
        RECT 160.175 41.735 160.345 45.660 ;
        RECT 172.830 45.660 175.175 45.690 ;
        RECT 175.975 45.660 178.320 45.785 ;
        RECT 172.830 40.805 173.000 45.660 ;
        RECT 173.340 40.810 173.630 45.660 ;
        RECT 177.520 40.810 177.810 45.660 ;
        RECT 178.150 40.805 178.320 45.660 ;
        RECT 2.970 35.260 3.140 39.675 ;
        RECT 3.480 35.260 3.770 39.670 ;
        RECT 2.970 35.230 5.065 35.260 ;
        RECT 2.970 35.145 5.220 35.230 ;
        RECT 6.200 35.145 6.370 38.120 ;
        RECT 2.970 34.975 6.370 35.145 ;
        RECT 14.500 35.260 14.670 39.860 ;
        RECT 15.010 35.260 15.300 40.090 ;
        RECT 19.190 35.260 19.480 40.090 ;
        RECT 19.820 35.260 19.990 39.920 ;
        RECT 14.500 35.095 16.845 35.260 ;
        RECT 17.645 35.095 19.990 35.260 ;
        RECT 2.970 34.810 5.220 34.975 ;
        RECT 14.500 34.925 19.990 35.095 ;
        RECT 2.970 34.780 5.065 34.810 ;
        RECT 14.500 34.780 16.845 34.925 ;
        RECT 17.645 34.780 19.990 34.925 ;
        RECT 32.470 35.260 32.640 39.675 ;
        RECT 32.980 35.260 33.270 39.670 ;
        RECT 32.470 35.230 34.565 35.260 ;
        RECT 32.470 35.145 34.720 35.230 ;
        RECT 35.700 35.145 35.870 38.120 ;
        RECT 32.470 34.975 35.870 35.145 ;
        RECT 44.000 35.260 44.170 39.860 ;
        RECT 44.510 35.260 44.800 40.090 ;
        RECT 48.690 35.260 48.980 40.090 ;
        RECT 49.320 35.260 49.490 39.920 ;
        RECT 44.000 35.095 46.345 35.260 ;
        RECT 47.145 35.095 49.490 35.260 ;
        RECT 32.470 34.810 34.720 34.975 ;
        RECT 44.000 34.925 49.490 35.095 ;
        RECT 32.470 34.780 34.565 34.810 ;
        RECT 44.000 34.780 46.345 34.925 ;
        RECT 47.145 34.780 49.490 34.925 ;
        RECT 61.970 35.260 62.140 39.675 ;
        RECT 62.480 35.260 62.770 39.670 ;
        RECT 61.970 35.230 64.065 35.260 ;
        RECT 61.970 35.145 64.220 35.230 ;
        RECT 65.200 35.145 65.370 38.120 ;
        RECT 61.970 34.975 65.370 35.145 ;
        RECT 73.500 35.260 73.670 39.860 ;
        RECT 74.010 35.260 74.300 40.090 ;
        RECT 78.190 35.260 78.480 40.090 ;
        RECT 78.820 35.260 78.990 39.920 ;
        RECT 73.500 35.095 75.845 35.260 ;
        RECT 76.645 35.095 78.990 35.260 ;
        RECT 61.970 34.810 64.220 34.975 ;
        RECT 73.500 34.925 78.990 35.095 ;
        RECT 61.970 34.780 64.065 34.810 ;
        RECT 73.500 34.780 75.845 34.925 ;
        RECT 76.645 34.780 78.990 34.925 ;
        RECT 91.470 35.260 91.640 39.675 ;
        RECT 91.980 35.260 92.270 39.670 ;
        RECT 91.470 35.230 93.565 35.260 ;
        RECT 91.470 35.145 93.720 35.230 ;
        RECT 94.700 35.145 94.870 38.120 ;
        RECT 91.470 34.975 94.870 35.145 ;
        RECT 103.000 35.260 103.170 39.860 ;
        RECT 103.510 35.260 103.800 40.090 ;
        RECT 107.690 35.260 107.980 40.090 ;
        RECT 108.320 35.260 108.490 39.920 ;
        RECT 103.000 35.095 105.345 35.260 ;
        RECT 106.145 35.095 108.490 35.260 ;
        RECT 91.470 34.810 93.720 34.975 ;
        RECT 103.000 34.925 108.490 35.095 ;
        RECT 91.470 34.780 93.565 34.810 ;
        RECT 103.000 34.780 105.345 34.925 ;
        RECT 106.145 34.780 108.490 34.925 ;
        RECT 120.970 35.260 121.140 39.675 ;
        RECT 121.480 35.260 121.770 39.670 ;
        RECT 120.970 35.230 123.065 35.260 ;
        RECT 120.970 35.145 123.220 35.230 ;
        RECT 124.200 35.145 124.370 38.120 ;
        RECT 120.970 34.975 124.370 35.145 ;
        RECT 132.500 35.260 132.670 39.860 ;
        RECT 133.010 35.260 133.300 40.090 ;
        RECT 137.190 35.260 137.480 40.090 ;
        RECT 137.820 35.260 137.990 39.920 ;
        RECT 132.500 35.095 134.845 35.260 ;
        RECT 135.645 35.095 137.990 35.260 ;
        RECT 120.970 34.810 123.220 34.975 ;
        RECT 132.500 34.925 137.990 35.095 ;
        RECT 120.970 34.780 123.065 34.810 ;
        RECT 132.500 34.780 134.845 34.925 ;
        RECT 135.645 34.780 137.990 34.925 ;
        RECT 150.470 35.260 150.640 39.675 ;
        RECT 150.980 35.260 151.270 39.670 ;
        RECT 150.470 35.230 152.565 35.260 ;
        RECT 150.470 35.145 152.720 35.230 ;
        RECT 153.700 35.145 153.870 38.120 ;
        RECT 150.470 34.975 153.870 35.145 ;
        RECT 162.000 35.260 162.170 39.860 ;
        RECT 162.510 35.260 162.800 40.090 ;
        RECT 166.690 35.260 166.980 40.090 ;
        RECT 167.320 35.260 167.490 39.920 ;
        RECT 162.000 35.095 164.345 35.260 ;
        RECT 165.145 35.095 167.490 35.260 ;
        RECT 150.470 34.810 152.720 34.975 ;
        RECT 162.000 34.925 167.490 35.095 ;
        RECT 150.470 34.780 152.565 34.810 ;
        RECT 162.000 34.780 164.345 34.925 ;
        RECT 165.145 34.780 167.490 34.925 ;
      LAYER mcon ;
        RECT 29.400 67.450 29.915 67.870 ;
        RECT 30.105 67.450 30.525 67.870 ;
        RECT 30.715 67.450 31.135 67.870 ;
        RECT 31.325 67.450 31.745 67.870 ;
        RECT 32.545 67.450 32.965 67.870 ;
        RECT 33.155 67.450 33.575 67.870 ;
        RECT 33.765 67.450 34.185 67.870 ;
        RECT 34.375 67.450 34.890 67.870 ;
        RECT 44.780 67.450 45.200 67.870 ;
        RECT 45.390 67.450 45.810 67.870 ;
        RECT 46.000 67.450 46.420 67.870 ;
        RECT 58.900 67.450 59.415 67.870 ;
        RECT 59.605 67.450 60.025 67.870 ;
        RECT 60.215 67.450 60.635 67.870 ;
        RECT 60.825 67.450 61.245 67.870 ;
        RECT 62.045 67.450 62.465 67.870 ;
        RECT 62.655 67.450 63.075 67.870 ;
        RECT 63.265 67.450 63.685 67.870 ;
        RECT 63.875 67.450 64.390 67.870 ;
        RECT 74.280 67.450 74.700 67.870 ;
        RECT 74.890 67.450 75.310 67.870 ;
        RECT 75.500 67.450 75.920 67.870 ;
        RECT 88.400 67.450 88.915 67.870 ;
        RECT 89.105 67.450 89.525 67.870 ;
        RECT 89.715 67.450 90.135 67.870 ;
        RECT 90.325 67.450 90.745 67.870 ;
        RECT 91.545 67.450 91.965 67.870 ;
        RECT 92.155 67.450 92.575 67.870 ;
        RECT 92.765 67.450 93.185 67.870 ;
        RECT 93.375 67.450 93.890 67.870 ;
        RECT 103.780 67.450 104.200 67.870 ;
        RECT 104.390 67.450 104.810 67.870 ;
        RECT 105.000 67.450 105.420 67.870 ;
        RECT 117.900 67.450 118.415 67.870 ;
        RECT 118.605 67.450 119.025 67.870 ;
        RECT 119.215 67.450 119.635 67.870 ;
        RECT 119.825 67.450 120.245 67.870 ;
        RECT 121.045 67.450 121.465 67.870 ;
        RECT 121.655 67.450 122.075 67.870 ;
        RECT 122.265 67.450 122.685 67.870 ;
        RECT 122.875 67.450 123.390 67.870 ;
        RECT 133.280 67.450 133.700 67.870 ;
        RECT 133.890 67.450 134.310 67.870 ;
        RECT 134.500 67.450 134.920 67.870 ;
        RECT 147.400 67.450 147.915 67.870 ;
        RECT 148.105 67.450 148.525 67.870 ;
        RECT 148.715 67.450 149.135 67.870 ;
        RECT 149.325 67.450 149.745 67.870 ;
        RECT 150.545 67.450 150.965 67.870 ;
        RECT 151.155 67.450 151.575 67.870 ;
        RECT 151.765 67.450 152.185 67.870 ;
        RECT 152.375 67.450 152.890 67.870 ;
        RECT 162.780 67.450 163.200 67.870 ;
        RECT 163.390 67.450 163.810 67.870 ;
        RECT 164.000 67.450 164.420 67.870 ;
        RECT 3.965 62.135 4.135 62.305 ;
        RECT 4.425 62.135 4.595 62.305 ;
        RECT 4.885 62.135 5.055 62.305 ;
        RECT 5.345 62.135 5.515 62.305 ;
        RECT 5.805 62.135 5.975 62.305 ;
        RECT 8.135 62.135 8.305 62.305 ;
        RECT 8.595 62.135 8.765 62.305 ;
        RECT 9.055 62.135 9.225 62.305 ;
        RECT 18.570 56.570 19.085 56.990 ;
        RECT 19.275 56.570 19.695 56.990 ;
        RECT 19.885 56.570 20.305 56.990 ;
        RECT 20.495 56.570 20.915 56.990 ;
        RECT 21.895 56.570 22.315 56.990 ;
        RECT 22.505 56.570 22.925 56.990 ;
        RECT 23.115 56.570 23.535 56.990 ;
        RECT 23.725 56.570 24.240 56.990 ;
        RECT 37.155 56.570 37.575 56.990 ;
        RECT 37.765 56.570 38.185 56.990 ;
        RECT 38.375 56.570 38.795 56.990 ;
        RECT 48.070 56.570 48.585 56.990 ;
        RECT 48.775 56.570 49.195 56.990 ;
        RECT 49.385 56.570 49.805 56.990 ;
        RECT 49.995 56.570 50.415 56.990 ;
        RECT 51.395 56.570 51.815 56.990 ;
        RECT 52.005 56.570 52.425 56.990 ;
        RECT 52.615 56.570 53.035 56.990 ;
        RECT 53.225 56.570 53.740 56.990 ;
        RECT 66.655 56.570 67.075 56.990 ;
        RECT 67.265 56.570 67.685 56.990 ;
        RECT 67.875 56.570 68.295 56.990 ;
        RECT 77.570 56.570 78.085 56.990 ;
        RECT 78.275 56.570 78.695 56.990 ;
        RECT 78.885 56.570 79.305 56.990 ;
        RECT 79.495 56.570 79.915 56.990 ;
        RECT 80.895 56.570 81.315 56.990 ;
        RECT 81.505 56.570 81.925 56.990 ;
        RECT 82.115 56.570 82.535 56.990 ;
        RECT 82.725 56.570 83.240 56.990 ;
        RECT 96.155 56.570 96.575 56.990 ;
        RECT 96.765 56.570 97.185 56.990 ;
        RECT 97.375 56.570 97.795 56.990 ;
        RECT 107.070 56.570 107.585 56.990 ;
        RECT 107.775 56.570 108.195 56.990 ;
        RECT 108.385 56.570 108.805 56.990 ;
        RECT 108.995 56.570 109.415 56.990 ;
        RECT 110.395 56.570 110.815 56.990 ;
        RECT 111.005 56.570 111.425 56.990 ;
        RECT 111.615 56.570 112.035 56.990 ;
        RECT 112.225 56.570 112.740 56.990 ;
        RECT 125.655 56.570 126.075 56.990 ;
        RECT 126.265 56.570 126.685 56.990 ;
        RECT 126.875 56.570 127.295 56.990 ;
        RECT 136.570 56.570 137.085 56.990 ;
        RECT 137.275 56.570 137.695 56.990 ;
        RECT 137.885 56.570 138.305 56.990 ;
        RECT 138.495 56.570 138.915 56.990 ;
        RECT 139.895 56.570 140.315 56.990 ;
        RECT 140.505 56.570 140.925 56.990 ;
        RECT 141.115 56.570 141.535 56.990 ;
        RECT 141.725 56.570 142.240 56.990 ;
        RECT 155.155 56.570 155.575 56.990 ;
        RECT 155.765 56.570 156.185 56.990 ;
        RECT 156.375 56.570 156.795 56.990 ;
        RECT 11.205 45.690 11.625 46.110 ;
        RECT 11.815 45.690 12.235 46.110 ;
        RECT 12.425 45.690 12.845 46.110 ;
        RECT 25.855 45.690 26.275 46.110 ;
        RECT 26.465 45.690 26.885 46.110 ;
        RECT 27.075 45.690 27.495 46.110 ;
        RECT 28.475 45.690 28.895 46.110 ;
        RECT 29.085 45.690 29.505 46.110 ;
        RECT 29.695 45.690 30.115 46.110 ;
        RECT 30.305 45.690 30.820 46.110 ;
        RECT 40.705 45.690 41.125 46.110 ;
        RECT 41.315 45.690 41.735 46.110 ;
        RECT 41.925 45.690 42.345 46.110 ;
        RECT 55.355 45.690 55.775 46.110 ;
        RECT 55.965 45.690 56.385 46.110 ;
        RECT 56.575 45.690 56.995 46.110 ;
        RECT 57.975 45.690 58.395 46.110 ;
        RECT 58.585 45.690 59.005 46.110 ;
        RECT 59.195 45.690 59.615 46.110 ;
        RECT 59.805 45.690 60.320 46.110 ;
        RECT 70.205 45.690 70.625 46.110 ;
        RECT 70.815 45.690 71.235 46.110 ;
        RECT 71.425 45.690 71.845 46.110 ;
        RECT 84.855 45.690 85.275 46.110 ;
        RECT 85.465 45.690 85.885 46.110 ;
        RECT 86.075 45.690 86.495 46.110 ;
        RECT 87.475 45.690 87.895 46.110 ;
        RECT 88.085 45.690 88.505 46.110 ;
        RECT 88.695 45.690 89.115 46.110 ;
        RECT 89.305 45.690 89.820 46.110 ;
        RECT 99.705 45.690 100.125 46.110 ;
        RECT 100.315 45.690 100.735 46.110 ;
        RECT 100.925 45.690 101.345 46.110 ;
        RECT 114.355 45.690 114.775 46.110 ;
        RECT 114.965 45.690 115.385 46.110 ;
        RECT 115.575 45.690 115.995 46.110 ;
        RECT 116.975 45.690 117.395 46.110 ;
        RECT 117.585 45.690 118.005 46.110 ;
        RECT 118.195 45.690 118.615 46.110 ;
        RECT 118.805 45.690 119.320 46.110 ;
        RECT 129.205 45.690 129.625 46.110 ;
        RECT 129.815 45.690 130.235 46.110 ;
        RECT 130.425 45.690 130.845 46.110 ;
        RECT 143.855 45.690 144.275 46.110 ;
        RECT 144.465 45.690 144.885 46.110 ;
        RECT 145.075 45.690 145.495 46.110 ;
        RECT 146.475 45.690 146.895 46.110 ;
        RECT 147.085 45.690 147.505 46.110 ;
        RECT 147.695 45.690 148.115 46.110 ;
        RECT 148.305 45.690 148.820 46.110 ;
        RECT 158.705 45.690 159.125 46.110 ;
        RECT 159.315 45.690 159.735 46.110 ;
        RECT 159.925 45.690 160.345 46.110 ;
        RECT 173.355 45.690 173.775 46.110 ;
        RECT 173.965 45.690 174.385 46.110 ;
        RECT 174.575 45.690 174.995 46.110 ;
        RECT 175.975 45.690 176.395 46.110 ;
        RECT 176.585 45.690 177.005 46.110 ;
        RECT 177.195 45.690 177.615 46.110 ;
        RECT 177.805 45.690 178.320 46.110 ;
        RECT 3.580 34.810 4.000 35.230 ;
        RECT 4.190 34.810 4.610 35.230 ;
        RECT 4.800 34.810 5.220 35.230 ;
        RECT 14.500 34.810 15.015 35.230 ;
        RECT 15.205 34.810 15.625 35.230 ;
        RECT 15.815 34.810 16.235 35.230 ;
        RECT 16.425 34.810 16.845 35.230 ;
        RECT 17.645 34.810 18.065 35.230 ;
        RECT 18.255 34.810 18.675 35.230 ;
        RECT 18.865 34.810 19.285 35.230 ;
        RECT 19.475 34.810 19.990 35.230 ;
        RECT 33.080 34.810 33.500 35.230 ;
        RECT 33.690 34.810 34.110 35.230 ;
        RECT 34.300 34.810 34.720 35.230 ;
        RECT 44.000 34.810 44.515 35.230 ;
        RECT 44.705 34.810 45.125 35.230 ;
        RECT 45.315 34.810 45.735 35.230 ;
        RECT 45.925 34.810 46.345 35.230 ;
        RECT 47.145 34.810 47.565 35.230 ;
        RECT 47.755 34.810 48.175 35.230 ;
        RECT 48.365 34.810 48.785 35.230 ;
        RECT 48.975 34.810 49.490 35.230 ;
        RECT 62.580 34.810 63.000 35.230 ;
        RECT 63.190 34.810 63.610 35.230 ;
        RECT 63.800 34.810 64.220 35.230 ;
        RECT 73.500 34.810 74.015 35.230 ;
        RECT 74.205 34.810 74.625 35.230 ;
        RECT 74.815 34.810 75.235 35.230 ;
        RECT 75.425 34.810 75.845 35.230 ;
        RECT 76.645 34.810 77.065 35.230 ;
        RECT 77.255 34.810 77.675 35.230 ;
        RECT 77.865 34.810 78.285 35.230 ;
        RECT 78.475 34.810 78.990 35.230 ;
        RECT 92.080 34.810 92.500 35.230 ;
        RECT 92.690 34.810 93.110 35.230 ;
        RECT 93.300 34.810 93.720 35.230 ;
        RECT 103.000 34.810 103.515 35.230 ;
        RECT 103.705 34.810 104.125 35.230 ;
        RECT 104.315 34.810 104.735 35.230 ;
        RECT 104.925 34.810 105.345 35.230 ;
        RECT 106.145 34.810 106.565 35.230 ;
        RECT 106.755 34.810 107.175 35.230 ;
        RECT 107.365 34.810 107.785 35.230 ;
        RECT 107.975 34.810 108.490 35.230 ;
        RECT 121.580 34.810 122.000 35.230 ;
        RECT 122.190 34.810 122.610 35.230 ;
        RECT 122.800 34.810 123.220 35.230 ;
        RECT 132.500 34.810 133.015 35.230 ;
        RECT 133.205 34.810 133.625 35.230 ;
        RECT 133.815 34.810 134.235 35.230 ;
        RECT 134.425 34.810 134.845 35.230 ;
        RECT 135.645 34.810 136.065 35.230 ;
        RECT 136.255 34.810 136.675 35.230 ;
        RECT 136.865 34.810 137.285 35.230 ;
        RECT 137.475 34.810 137.990 35.230 ;
        RECT 151.080 34.810 151.500 35.230 ;
        RECT 151.690 34.810 152.110 35.230 ;
        RECT 152.300 34.810 152.720 35.230 ;
        RECT 162.000 34.810 162.515 35.230 ;
        RECT 162.705 34.810 163.125 35.230 ;
        RECT 163.315 34.810 163.735 35.230 ;
        RECT 163.925 34.810 164.345 35.230 ;
        RECT 165.145 34.810 165.565 35.230 ;
        RECT 165.755 34.810 166.175 35.230 ;
        RECT 166.365 34.810 166.785 35.230 ;
        RECT 166.975 34.810 167.490 35.230 ;
      LAYER met1 ;
        RECT 16.000 67.420 165.390 67.900 ;
        RECT 3.820 61.980 20.490 62.460 ;
        RECT 15.005 56.540 172.440 57.020 ;
        RECT 162.490 56.535 164.490 56.540 ;
        RECT 0.000 45.660 179.445 46.140 ;
        RECT 0.000 34.780 179.440 35.260 ;
      LAYER via ;
        RECT 18.620 67.510 18.920 67.810 ;
        RECT 18.980 67.510 19.280 67.810 ;
        RECT 19.340 67.510 19.640 67.810 ;
        RECT 19.700 67.510 20.000 67.810 ;
        RECT 20.060 67.510 20.360 67.810 ;
        RECT 54.620 67.510 54.920 67.810 ;
        RECT 54.980 67.510 55.280 67.810 ;
        RECT 55.340 67.510 55.640 67.810 ;
        RECT 55.700 67.510 56.000 67.810 ;
        RECT 56.060 67.510 56.360 67.810 ;
        RECT 90.620 67.510 90.920 67.810 ;
        RECT 90.980 67.510 91.280 67.810 ;
        RECT 91.340 67.510 91.640 67.810 ;
        RECT 91.700 67.510 92.000 67.810 ;
        RECT 92.060 67.510 92.360 67.810 ;
        RECT 126.620 67.510 126.920 67.810 ;
        RECT 126.980 67.510 127.280 67.810 ;
        RECT 127.340 67.510 127.640 67.810 ;
        RECT 127.700 67.510 128.000 67.810 ;
        RECT 128.060 67.510 128.360 67.810 ;
        RECT 162.620 67.510 162.920 67.810 ;
        RECT 162.980 67.510 163.280 67.810 ;
        RECT 163.340 67.510 163.640 67.810 ;
        RECT 163.700 67.510 164.000 67.810 ;
        RECT 164.060 67.510 164.360 67.810 ;
        RECT 18.620 62.070 18.920 62.370 ;
        RECT 18.980 62.070 19.280 62.370 ;
        RECT 19.340 62.070 19.640 62.370 ;
        RECT 19.700 62.070 20.000 62.370 ;
        RECT 20.060 62.070 20.360 62.370 ;
        RECT 18.620 56.630 18.920 56.930 ;
        RECT 18.980 56.630 19.280 56.930 ;
        RECT 19.340 56.630 19.640 56.930 ;
        RECT 19.700 56.630 20.000 56.930 ;
        RECT 20.060 56.630 20.360 56.930 ;
        RECT 54.620 56.630 54.920 56.930 ;
        RECT 54.980 56.630 55.280 56.930 ;
        RECT 55.340 56.630 55.640 56.930 ;
        RECT 55.700 56.630 56.000 56.930 ;
        RECT 56.060 56.630 56.360 56.930 ;
        RECT 90.620 56.630 90.920 56.930 ;
        RECT 90.980 56.630 91.280 56.930 ;
        RECT 91.340 56.630 91.640 56.930 ;
        RECT 91.700 56.630 92.000 56.930 ;
        RECT 92.060 56.630 92.360 56.930 ;
        RECT 126.620 56.630 126.920 56.930 ;
        RECT 126.980 56.630 127.280 56.930 ;
        RECT 127.340 56.630 127.640 56.930 ;
        RECT 127.700 56.630 128.000 56.930 ;
        RECT 128.060 56.630 128.360 56.930 ;
        RECT 162.620 56.625 162.920 56.925 ;
        RECT 162.980 56.625 163.280 56.925 ;
        RECT 163.340 56.625 163.640 56.925 ;
        RECT 163.700 56.625 164.000 56.925 ;
        RECT 164.060 56.625 164.360 56.925 ;
        RECT 18.620 45.750 18.920 46.050 ;
        RECT 18.980 45.750 19.280 46.050 ;
        RECT 19.340 45.750 19.640 46.050 ;
        RECT 19.700 45.750 20.000 46.050 ;
        RECT 20.060 45.750 20.360 46.050 ;
        RECT 54.620 45.750 54.920 46.050 ;
        RECT 54.980 45.750 55.280 46.050 ;
        RECT 55.340 45.750 55.640 46.050 ;
        RECT 55.700 45.750 56.000 46.050 ;
        RECT 56.060 45.750 56.360 46.050 ;
        RECT 90.620 45.750 90.920 46.050 ;
        RECT 90.980 45.750 91.280 46.050 ;
        RECT 91.340 45.750 91.640 46.050 ;
        RECT 91.700 45.750 92.000 46.050 ;
        RECT 92.060 45.750 92.360 46.050 ;
        RECT 126.620 45.750 126.920 46.050 ;
        RECT 126.980 45.750 127.280 46.050 ;
        RECT 127.340 45.750 127.640 46.050 ;
        RECT 127.700 45.750 128.000 46.050 ;
        RECT 128.060 45.750 128.360 46.050 ;
        RECT 162.620 45.750 162.920 46.050 ;
        RECT 162.980 45.750 163.280 46.050 ;
        RECT 163.340 45.750 163.640 46.050 ;
        RECT 163.700 45.750 164.000 46.050 ;
        RECT 164.060 45.750 164.360 46.050 ;
        RECT 18.620 34.870 18.920 35.170 ;
        RECT 18.980 34.870 19.280 35.170 ;
        RECT 19.340 34.870 19.640 35.170 ;
        RECT 19.700 34.870 20.000 35.170 ;
        RECT 20.060 34.870 20.360 35.170 ;
        RECT 54.620 34.870 54.920 35.170 ;
        RECT 54.980 34.870 55.280 35.170 ;
        RECT 55.340 34.870 55.640 35.170 ;
        RECT 55.700 34.870 56.000 35.170 ;
        RECT 56.060 34.870 56.360 35.170 ;
        RECT 126.620 34.870 126.920 35.170 ;
        RECT 126.980 34.870 127.280 35.170 ;
        RECT 127.340 34.870 127.640 35.170 ;
        RECT 127.700 34.870 128.000 35.170 ;
        RECT 128.060 34.870 128.360 35.170 ;
        RECT 162.620 34.870 162.920 35.170 ;
        RECT 162.980 34.870 163.280 35.170 ;
        RECT 163.340 34.870 163.640 35.170 ;
        RECT 163.700 34.870 164.000 35.170 ;
        RECT 164.060 34.870 164.360 35.170 ;
      LAYER met2 ;
        RECT 18.490 67.420 20.490 67.900 ;
        RECT 54.490 67.420 56.490 67.900 ;
        RECT 90.490 67.420 92.490 67.900 ;
        RECT 126.490 67.420 128.490 67.900 ;
        RECT 162.490 67.420 164.490 67.900 ;
        RECT 18.490 61.980 20.490 62.460 ;
        RECT 18.490 56.540 20.490 57.020 ;
        RECT 54.490 56.540 56.490 57.020 ;
        RECT 90.490 56.540 92.490 57.020 ;
        RECT 126.490 56.540 128.490 57.020 ;
        RECT 162.490 56.535 164.490 57.020 ;
        RECT 18.490 45.660 20.490 46.140 ;
        RECT 54.490 45.660 56.490 46.140 ;
        RECT 90.490 45.660 92.490 46.140 ;
        RECT 126.490 45.660 128.490 46.140 ;
        RECT 162.490 45.660 164.490 46.140 ;
        RECT 18.490 34.780 20.490 35.260 ;
        RECT 54.490 34.780 56.490 35.260 ;
        RECT 126.490 34.780 128.490 35.260 ;
        RECT 162.490 34.780 164.490 35.260 ;
      LAYER via2 ;
        RECT 18.670 67.500 18.990 67.820 ;
        RECT 19.110 67.500 19.430 67.820 ;
        RECT 19.550 67.500 19.870 67.820 ;
        RECT 19.990 67.500 20.310 67.820 ;
        RECT 54.670 67.500 54.990 67.820 ;
        RECT 55.110 67.500 55.430 67.820 ;
        RECT 55.550 67.500 55.870 67.820 ;
        RECT 55.990 67.500 56.310 67.820 ;
        RECT 90.670 67.500 90.990 67.820 ;
        RECT 91.110 67.500 91.430 67.820 ;
        RECT 91.550 67.500 91.870 67.820 ;
        RECT 91.990 67.500 92.310 67.820 ;
        RECT 126.670 67.500 126.990 67.820 ;
        RECT 127.110 67.500 127.430 67.820 ;
        RECT 127.550 67.500 127.870 67.820 ;
        RECT 127.990 67.500 128.310 67.820 ;
        RECT 162.670 67.500 162.990 67.820 ;
        RECT 163.110 67.500 163.430 67.820 ;
        RECT 163.550 67.500 163.870 67.820 ;
        RECT 163.990 67.500 164.310 67.820 ;
        RECT 18.670 62.060 18.990 62.380 ;
        RECT 19.110 62.060 19.430 62.380 ;
        RECT 19.550 62.060 19.870 62.380 ;
        RECT 19.990 62.060 20.310 62.380 ;
        RECT 18.670 56.620 18.990 56.940 ;
        RECT 19.110 56.620 19.430 56.940 ;
        RECT 19.550 56.620 19.870 56.940 ;
        RECT 19.990 56.620 20.310 56.940 ;
        RECT 54.670 56.620 54.990 56.940 ;
        RECT 55.110 56.620 55.430 56.940 ;
        RECT 55.550 56.620 55.870 56.940 ;
        RECT 55.990 56.620 56.310 56.940 ;
        RECT 90.670 56.620 90.990 56.940 ;
        RECT 91.110 56.620 91.430 56.940 ;
        RECT 91.550 56.620 91.870 56.940 ;
        RECT 91.990 56.620 92.310 56.940 ;
        RECT 126.670 56.620 126.990 56.940 ;
        RECT 127.110 56.620 127.430 56.940 ;
        RECT 127.550 56.620 127.870 56.940 ;
        RECT 127.990 56.620 128.310 56.940 ;
        RECT 162.670 56.615 162.990 56.935 ;
        RECT 163.110 56.615 163.430 56.935 ;
        RECT 163.550 56.615 163.870 56.935 ;
        RECT 163.990 56.615 164.310 56.935 ;
        RECT 18.670 45.740 18.990 46.060 ;
        RECT 19.110 45.740 19.430 46.060 ;
        RECT 19.550 45.740 19.870 46.060 ;
        RECT 19.990 45.740 20.310 46.060 ;
        RECT 54.670 45.740 54.990 46.060 ;
        RECT 55.110 45.740 55.430 46.060 ;
        RECT 55.550 45.740 55.870 46.060 ;
        RECT 55.990 45.740 56.310 46.060 ;
        RECT 90.670 45.740 90.990 46.060 ;
        RECT 91.110 45.740 91.430 46.060 ;
        RECT 91.550 45.740 91.870 46.060 ;
        RECT 91.990 45.740 92.310 46.060 ;
        RECT 126.670 45.740 126.990 46.060 ;
        RECT 127.110 45.740 127.430 46.060 ;
        RECT 127.550 45.740 127.870 46.060 ;
        RECT 127.990 45.740 128.310 46.060 ;
        RECT 162.670 45.740 162.990 46.060 ;
        RECT 163.110 45.740 163.430 46.060 ;
        RECT 163.550 45.740 163.870 46.060 ;
        RECT 163.990 45.740 164.310 46.060 ;
        RECT 18.670 34.860 18.990 35.180 ;
        RECT 19.110 34.860 19.430 35.180 ;
        RECT 19.550 34.860 19.870 35.180 ;
        RECT 19.990 34.860 20.310 35.180 ;
        RECT 54.670 34.860 54.990 35.180 ;
        RECT 55.110 34.860 55.430 35.180 ;
        RECT 55.550 34.860 55.870 35.180 ;
        RECT 55.990 34.860 56.310 35.180 ;
        RECT 126.670 34.860 126.990 35.180 ;
        RECT 127.110 34.860 127.430 35.180 ;
        RECT 127.550 34.860 127.870 35.180 ;
        RECT 127.990 34.860 128.310 35.180 ;
        RECT 162.670 34.860 162.990 35.180 ;
        RECT 163.110 34.860 163.430 35.180 ;
        RECT 163.550 34.860 163.870 35.180 ;
        RECT 163.990 34.860 164.310 35.180 ;
      LAYER met3 ;
        RECT 5.490 102.000 177.490 104.000 ;
        RECT 18.490 67.420 20.490 67.900 ;
        RECT 54.490 67.420 56.490 67.900 ;
        RECT 90.490 67.420 92.490 67.900 ;
        RECT 126.490 67.420 128.490 67.900 ;
        RECT 162.490 67.420 164.490 67.900 ;
        RECT 18.490 61.980 20.490 62.460 ;
        RECT 18.490 56.540 20.490 57.020 ;
        RECT 54.490 56.540 56.490 57.020 ;
        RECT 90.490 56.540 92.490 57.020 ;
        RECT 126.490 56.540 128.490 57.020 ;
        RECT 162.490 56.535 164.490 57.020 ;
        RECT 18.490 45.660 20.490 46.140 ;
        RECT 54.490 45.660 56.490 46.140 ;
        RECT 90.490 45.660 92.490 46.140 ;
        RECT 126.490 45.660 128.490 46.140 ;
        RECT 162.490 45.660 164.490 46.140 ;
        RECT 18.490 34.780 20.490 35.260 ;
        RECT 54.490 34.780 56.490 35.260 ;
        RECT 126.490 34.780 128.490 35.260 ;
        RECT 162.490 34.780 164.490 35.260 ;
        RECT 5.490 -1.000 177.490 1.000 ;
      LAYER via3 ;
        RECT 5.690 103.400 6.090 103.800 ;
        RECT 6.290 103.400 6.690 103.800 ;
        RECT 6.890 103.400 7.290 103.800 ;
        RECT 18.690 103.400 19.090 103.800 ;
        RECT 19.290 103.400 19.690 103.800 ;
        RECT 19.890 103.400 20.290 103.800 ;
        RECT 54.690 103.400 55.090 103.800 ;
        RECT 55.290 103.400 55.690 103.800 ;
        RECT 55.890 103.400 56.290 103.800 ;
        RECT 90.690 103.400 91.090 103.800 ;
        RECT 91.290 103.400 91.690 103.800 ;
        RECT 91.890 103.400 92.290 103.800 ;
        RECT 126.690 103.400 127.090 103.800 ;
        RECT 127.290 103.400 127.690 103.800 ;
        RECT 127.890 103.400 128.290 103.800 ;
        RECT 162.690 103.400 163.090 103.800 ;
        RECT 163.290 103.400 163.690 103.800 ;
        RECT 163.890 103.400 164.290 103.800 ;
        RECT 175.690 103.400 176.090 103.800 ;
        RECT 176.290 103.400 176.690 103.800 ;
        RECT 176.890 103.400 177.290 103.800 ;
        RECT 5.690 102.800 6.090 103.200 ;
        RECT 6.290 102.800 6.690 103.200 ;
        RECT 6.890 102.800 7.290 103.200 ;
        RECT 18.690 102.800 19.090 103.200 ;
        RECT 19.290 102.800 19.690 103.200 ;
        RECT 19.890 102.800 20.290 103.200 ;
        RECT 54.690 102.800 55.090 103.200 ;
        RECT 55.290 102.800 55.690 103.200 ;
        RECT 55.890 102.800 56.290 103.200 ;
        RECT 90.690 102.800 91.090 103.200 ;
        RECT 91.290 102.800 91.690 103.200 ;
        RECT 91.890 102.800 92.290 103.200 ;
        RECT 126.690 102.800 127.090 103.200 ;
        RECT 127.290 102.800 127.690 103.200 ;
        RECT 127.890 102.800 128.290 103.200 ;
        RECT 162.690 102.800 163.090 103.200 ;
        RECT 163.290 102.800 163.690 103.200 ;
        RECT 163.890 102.800 164.290 103.200 ;
        RECT 175.690 102.800 176.090 103.200 ;
        RECT 176.290 102.800 176.690 103.200 ;
        RECT 176.890 102.800 177.290 103.200 ;
        RECT 5.690 102.200 6.090 102.600 ;
        RECT 6.290 102.200 6.690 102.600 ;
        RECT 6.890 102.200 7.290 102.600 ;
        RECT 18.690 102.200 19.090 102.600 ;
        RECT 19.290 102.200 19.690 102.600 ;
        RECT 19.890 102.200 20.290 102.600 ;
        RECT 54.690 102.200 55.090 102.600 ;
        RECT 55.290 102.200 55.690 102.600 ;
        RECT 55.890 102.200 56.290 102.600 ;
        RECT 90.690 102.200 91.090 102.600 ;
        RECT 91.290 102.200 91.690 102.600 ;
        RECT 91.890 102.200 92.290 102.600 ;
        RECT 126.690 102.200 127.090 102.600 ;
        RECT 127.290 102.200 127.690 102.600 ;
        RECT 127.890 102.200 128.290 102.600 ;
        RECT 162.690 102.200 163.090 102.600 ;
        RECT 163.290 102.200 163.690 102.600 ;
        RECT 163.890 102.200 164.290 102.600 ;
        RECT 175.690 102.200 176.090 102.600 ;
        RECT 176.290 102.200 176.690 102.600 ;
        RECT 176.890 102.200 177.290 102.600 ;
        RECT 18.650 67.480 19.010 67.840 ;
        RECT 19.090 67.480 19.450 67.840 ;
        RECT 19.530 67.480 19.890 67.840 ;
        RECT 19.970 67.480 20.330 67.840 ;
        RECT 54.650 67.480 55.010 67.840 ;
        RECT 55.090 67.480 55.450 67.840 ;
        RECT 55.530 67.480 55.890 67.840 ;
        RECT 55.970 67.480 56.330 67.840 ;
        RECT 90.650 67.480 91.010 67.840 ;
        RECT 91.090 67.480 91.450 67.840 ;
        RECT 91.530 67.480 91.890 67.840 ;
        RECT 91.970 67.480 92.330 67.840 ;
        RECT 126.650 67.480 127.010 67.840 ;
        RECT 127.090 67.480 127.450 67.840 ;
        RECT 127.530 67.480 127.890 67.840 ;
        RECT 127.970 67.480 128.330 67.840 ;
        RECT 162.650 67.480 163.010 67.840 ;
        RECT 163.090 67.480 163.450 67.840 ;
        RECT 163.530 67.480 163.890 67.840 ;
        RECT 163.970 67.480 164.330 67.840 ;
        RECT 18.650 62.040 19.010 62.400 ;
        RECT 19.090 62.040 19.450 62.400 ;
        RECT 19.530 62.040 19.890 62.400 ;
        RECT 19.970 62.040 20.330 62.400 ;
        RECT 18.650 56.600 19.010 56.960 ;
        RECT 19.090 56.600 19.450 56.960 ;
        RECT 19.530 56.600 19.890 56.960 ;
        RECT 19.970 56.600 20.330 56.960 ;
        RECT 54.650 56.600 55.010 56.960 ;
        RECT 55.090 56.600 55.450 56.960 ;
        RECT 55.530 56.600 55.890 56.960 ;
        RECT 55.970 56.600 56.330 56.960 ;
        RECT 90.650 56.600 91.010 56.960 ;
        RECT 91.090 56.600 91.450 56.960 ;
        RECT 91.530 56.600 91.890 56.960 ;
        RECT 91.970 56.600 92.330 56.960 ;
        RECT 126.650 56.600 127.010 56.960 ;
        RECT 127.090 56.600 127.450 56.960 ;
        RECT 127.530 56.600 127.890 56.960 ;
        RECT 127.970 56.600 128.330 56.960 ;
        RECT 162.650 56.595 163.010 56.960 ;
        RECT 163.090 56.595 163.450 56.960 ;
        RECT 163.530 56.595 163.890 56.960 ;
        RECT 163.970 56.595 164.330 56.960 ;
        RECT 18.650 45.720 19.010 46.085 ;
        RECT 19.090 45.720 19.450 46.085 ;
        RECT 19.530 45.720 19.890 46.085 ;
        RECT 19.970 45.720 20.330 46.085 ;
        RECT 54.650 45.720 55.010 46.085 ;
        RECT 55.090 45.720 55.450 46.085 ;
        RECT 55.530 45.720 55.890 46.085 ;
        RECT 55.970 45.720 56.330 46.085 ;
        RECT 90.650 45.720 91.010 46.085 ;
        RECT 91.090 45.720 91.450 46.085 ;
        RECT 91.530 45.720 91.890 46.085 ;
        RECT 91.970 45.720 92.330 46.085 ;
        RECT 126.650 45.720 127.010 46.085 ;
        RECT 127.090 45.720 127.450 46.085 ;
        RECT 127.530 45.720 127.890 46.085 ;
        RECT 127.970 45.720 128.330 46.085 ;
        RECT 162.650 45.720 163.010 46.085 ;
        RECT 163.090 45.720 163.450 46.085 ;
        RECT 163.530 45.720 163.890 46.085 ;
        RECT 163.970 45.720 164.330 46.085 ;
        RECT 18.650 34.840 19.010 35.205 ;
        RECT 19.090 34.840 19.450 35.205 ;
        RECT 19.530 34.840 19.890 35.205 ;
        RECT 19.970 34.840 20.330 35.205 ;
        RECT 54.650 34.840 55.010 35.205 ;
        RECT 55.090 34.840 55.450 35.205 ;
        RECT 55.530 34.840 55.890 35.205 ;
        RECT 55.970 34.840 56.330 35.205 ;
        RECT 126.650 34.840 127.010 35.205 ;
        RECT 127.090 34.840 127.450 35.205 ;
        RECT 127.530 34.840 127.890 35.205 ;
        RECT 127.970 34.840 128.330 35.205 ;
        RECT 162.650 34.840 163.010 35.205 ;
        RECT 163.090 34.840 163.450 35.205 ;
        RECT 163.530 34.840 163.890 35.205 ;
        RECT 163.970 34.840 164.330 35.205 ;
        RECT 5.690 0.400 6.090 0.800 ;
        RECT 6.290 0.400 6.690 0.800 ;
        RECT 6.890 0.400 7.290 0.800 ;
        RECT 18.690 0.400 19.090 0.800 ;
        RECT 19.290 0.400 19.690 0.800 ;
        RECT 19.890 0.400 20.290 0.800 ;
        RECT 54.690 0.400 55.090 0.800 ;
        RECT 55.290 0.400 55.690 0.800 ;
        RECT 55.890 0.400 56.290 0.800 ;
        RECT 90.690 0.400 91.090 0.800 ;
        RECT 91.290 0.400 91.690 0.800 ;
        RECT 91.890 0.400 92.290 0.800 ;
        RECT 126.690 0.400 127.090 0.800 ;
        RECT 127.290 0.400 127.690 0.800 ;
        RECT 127.890 0.400 128.290 0.800 ;
        RECT 162.690 0.400 163.090 0.800 ;
        RECT 163.290 0.400 163.690 0.800 ;
        RECT 163.890 0.400 164.290 0.800 ;
        RECT 175.690 0.400 176.090 0.800 ;
        RECT 176.290 0.400 176.690 0.800 ;
        RECT 176.890 0.400 177.290 0.800 ;
        RECT 5.690 -0.200 6.090 0.200 ;
        RECT 6.290 -0.200 6.690 0.200 ;
        RECT 6.890 -0.200 7.290 0.200 ;
        RECT 18.690 -0.200 19.090 0.200 ;
        RECT 19.290 -0.200 19.690 0.200 ;
        RECT 19.890 -0.200 20.290 0.200 ;
        RECT 54.690 -0.200 55.090 0.200 ;
        RECT 55.290 -0.200 55.690 0.200 ;
        RECT 55.890 -0.200 56.290 0.200 ;
        RECT 90.690 -0.200 91.090 0.200 ;
        RECT 91.290 -0.200 91.690 0.200 ;
        RECT 91.890 -0.200 92.290 0.200 ;
        RECT 126.690 -0.200 127.090 0.200 ;
        RECT 127.290 -0.200 127.690 0.200 ;
        RECT 127.890 -0.200 128.290 0.200 ;
        RECT 162.690 -0.200 163.090 0.200 ;
        RECT 163.290 -0.200 163.690 0.200 ;
        RECT 163.890 -0.200 164.290 0.200 ;
        RECT 175.690 -0.200 176.090 0.200 ;
        RECT 176.290 -0.200 176.690 0.200 ;
        RECT 176.890 -0.200 177.290 0.200 ;
        RECT 5.690 -0.800 6.090 -0.400 ;
        RECT 6.290 -0.800 6.690 -0.400 ;
        RECT 6.890 -0.800 7.290 -0.400 ;
        RECT 18.690 -0.800 19.090 -0.400 ;
        RECT 19.290 -0.800 19.690 -0.400 ;
        RECT 19.890 -0.800 20.290 -0.400 ;
        RECT 54.690 -0.800 55.090 -0.400 ;
        RECT 55.290 -0.800 55.690 -0.400 ;
        RECT 55.890 -0.800 56.290 -0.400 ;
        RECT 90.690 -0.800 91.090 -0.400 ;
        RECT 91.290 -0.800 91.690 -0.400 ;
        RECT 91.890 -0.800 92.290 -0.400 ;
        RECT 126.690 -0.800 127.090 -0.400 ;
        RECT 127.290 -0.800 127.690 -0.400 ;
        RECT 127.890 -0.800 128.290 -0.400 ;
        RECT 162.690 -0.800 163.090 -0.400 ;
        RECT 163.290 -0.800 163.690 -0.400 ;
        RECT 163.890 -0.800 164.290 -0.400 ;
        RECT 175.690 -0.800 176.090 -0.400 ;
        RECT 176.290 -0.800 176.690 -0.400 ;
        RECT 176.890 -0.800 177.290 -0.400 ;
      LAYER met4 ;
        RECT 5.490 -1.000 7.490 104.000 ;
        RECT 18.490 -1.000 20.490 104.000 ;
        RECT 54.490 -1.000 56.490 104.000 ;
        RECT 90.490 -1.000 92.490 104.000 ;
        RECT 126.490 -1.000 128.490 104.000 ;
        RECT 162.490 -1.000 164.490 104.000 ;
        RECT 175.490 -1.000 177.490 104.000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 15.920 72.000 166.580 72.500 ;
        RECT 4.335 59.585 5.270 59.985 ;
        RECT 8.765 59.585 9.105 60.245 ;
        RECT 3.820 59.415 6.120 59.585 ;
        RECT 7.990 59.415 9.370 59.585 ;
        RECT 16.000 52.500 16.500 72.000 ;
        RECT 166.000 52.500 166.500 72.000 ;
        RECT 172.420 58.500 174.420 58.670 ;
        RECT 172.500 58.470 174.340 58.500 ;
        RECT 15.920 52.000 166.580 52.500 ;
        RECT 0.920 50.000 180.580 50.500 ;
        RECT 1.000 30.500 1.500 50.000 ;
        RECT 180.000 30.500 180.500 50.000 ;
        RECT 0.920 30.000 180.580 30.500 ;
      LAYER mcon ;
        RECT 36.590 72.100 36.890 72.400 ;
        RECT 37.090 72.100 37.390 72.400 ;
        RECT 37.590 72.100 37.890 72.400 ;
        RECT 38.090 72.100 38.390 72.400 ;
        RECT 72.590 72.100 72.890 72.400 ;
        RECT 73.090 72.100 73.390 72.400 ;
        RECT 73.590 72.100 73.890 72.400 ;
        RECT 74.090 72.100 74.390 72.400 ;
        RECT 108.590 72.100 108.890 72.400 ;
        RECT 109.090 72.100 109.390 72.400 ;
        RECT 109.590 72.100 109.890 72.400 ;
        RECT 110.090 72.100 110.390 72.400 ;
        RECT 144.590 72.100 144.890 72.400 ;
        RECT 145.090 72.100 145.390 72.400 ;
        RECT 145.590 72.100 145.890 72.400 ;
        RECT 146.090 72.100 146.390 72.400 ;
        RECT 3.965 59.415 4.135 59.585 ;
        RECT 4.425 59.415 4.595 59.585 ;
        RECT 4.885 59.415 5.055 59.585 ;
        RECT 5.345 59.415 5.515 59.585 ;
        RECT 5.805 59.415 5.975 59.585 ;
        RECT 8.135 59.415 8.305 59.585 ;
        RECT 8.595 59.415 8.765 59.585 ;
        RECT 9.055 59.415 9.225 59.585 ;
        RECT 172.615 58.485 172.785 58.655 ;
        RECT 172.975 58.485 173.145 58.655 ;
        RECT 173.335 58.485 173.505 58.655 ;
        RECT 173.695 58.485 173.865 58.655 ;
        RECT 174.055 58.485 174.225 58.655 ;
        RECT 36.590 30.100 36.890 30.400 ;
        RECT 37.090 30.100 37.390 30.400 ;
        RECT 37.590 30.100 37.890 30.400 ;
        RECT 38.090 30.100 38.390 30.400 ;
        RECT 72.590 30.100 72.890 30.400 ;
        RECT 73.090 30.100 73.390 30.400 ;
        RECT 73.590 30.100 73.890 30.400 ;
        RECT 74.090 30.100 74.390 30.400 ;
        RECT 108.590 30.100 108.890 30.400 ;
        RECT 109.090 30.100 109.390 30.400 ;
        RECT 109.590 30.100 109.890 30.400 ;
        RECT 110.090 30.100 110.390 30.400 ;
        RECT 144.590 30.100 144.890 30.400 ;
        RECT 145.090 30.100 145.390 30.400 ;
        RECT 145.590 30.100 145.890 30.400 ;
        RECT 146.090 30.100 146.390 30.400 ;
      LAYER met1 ;
        RECT 36.490 72.000 38.490 72.500 ;
        RECT 72.490 72.000 74.490 72.500 ;
        RECT 108.490 72.000 110.490 72.500 ;
        RECT 144.490 72.000 146.490 72.500 ;
        RECT 0.000 59.260 9.965 59.740 ;
        RECT 171.590 59.260 182.490 59.740 ;
        RECT 172.440 58.440 174.400 59.260 ;
        RECT 36.490 30.000 38.490 30.500 ;
        RECT 72.490 30.000 74.490 30.500 ;
        RECT 108.490 30.000 110.490 30.500 ;
        RECT 144.490 30.000 146.490 30.500 ;
      LAYER via ;
        RECT 36.620 72.100 36.920 72.400 ;
        RECT 36.980 72.100 37.280 72.400 ;
        RECT 37.340 72.100 37.640 72.400 ;
        RECT 37.700 72.100 38.000 72.400 ;
        RECT 38.060 72.100 38.360 72.400 ;
        RECT 72.620 72.100 72.920 72.400 ;
        RECT 72.980 72.100 73.280 72.400 ;
        RECT 73.340 72.100 73.640 72.400 ;
        RECT 73.700 72.100 74.000 72.400 ;
        RECT 74.060 72.100 74.360 72.400 ;
        RECT 108.620 72.100 108.920 72.400 ;
        RECT 108.980 72.100 109.280 72.400 ;
        RECT 109.340 72.100 109.640 72.400 ;
        RECT 109.700 72.100 110.000 72.400 ;
        RECT 110.060 72.100 110.360 72.400 ;
        RECT 144.620 72.100 144.920 72.400 ;
        RECT 144.980 72.100 145.280 72.400 ;
        RECT 145.340 72.100 145.640 72.400 ;
        RECT 145.700 72.100 146.000 72.400 ;
        RECT 146.060 72.100 146.360 72.400 ;
        RECT 0.620 59.350 0.920 59.650 ;
        RECT 0.980 59.350 1.280 59.650 ;
        RECT 1.340 59.350 1.640 59.650 ;
        RECT 1.700 59.350 2.000 59.650 ;
        RECT 2.060 59.350 2.360 59.650 ;
        RECT 180.620 59.350 180.920 59.650 ;
        RECT 180.980 59.350 181.280 59.650 ;
        RECT 181.340 59.350 181.640 59.650 ;
        RECT 181.700 59.350 182.000 59.650 ;
        RECT 182.060 59.350 182.360 59.650 ;
        RECT 36.620 30.100 36.920 30.400 ;
        RECT 36.980 30.100 37.280 30.400 ;
        RECT 37.340 30.100 37.640 30.400 ;
        RECT 37.700 30.100 38.000 30.400 ;
        RECT 38.060 30.100 38.360 30.400 ;
        RECT 72.620 30.100 72.920 30.400 ;
        RECT 72.980 30.100 73.280 30.400 ;
        RECT 73.340 30.100 73.640 30.400 ;
        RECT 73.700 30.100 74.000 30.400 ;
        RECT 74.060 30.100 74.360 30.400 ;
        RECT 108.620 30.100 108.920 30.400 ;
        RECT 108.980 30.100 109.280 30.400 ;
        RECT 109.340 30.100 109.640 30.400 ;
        RECT 109.700 30.100 110.000 30.400 ;
        RECT 110.060 30.100 110.360 30.400 ;
        RECT 144.620 30.100 144.920 30.400 ;
        RECT 144.980 30.100 145.280 30.400 ;
        RECT 145.340 30.100 145.640 30.400 ;
        RECT 145.700 30.100 146.000 30.400 ;
        RECT 146.060 30.100 146.360 30.400 ;
      LAYER met2 ;
        RECT 36.490 72.000 38.490 72.500 ;
        RECT 72.490 72.000 74.490 72.500 ;
        RECT 108.490 72.000 110.490 72.500 ;
        RECT 144.490 72.000 146.490 72.500 ;
        RECT 0.490 59.260 2.490 59.740 ;
        RECT 180.490 59.260 182.490 59.740 ;
        RECT 36.490 30.000 38.490 30.500 ;
        RECT 72.490 30.000 74.490 30.500 ;
        RECT 108.490 30.000 110.490 30.500 ;
        RECT 144.490 30.000 146.490 30.500 ;
      LAYER via2 ;
        RECT 36.670 72.090 36.990 72.410 ;
        RECT 37.110 72.090 37.430 72.410 ;
        RECT 37.550 72.090 37.870 72.410 ;
        RECT 37.990 72.090 38.310 72.410 ;
        RECT 72.670 72.090 72.990 72.410 ;
        RECT 73.110 72.090 73.430 72.410 ;
        RECT 73.550 72.090 73.870 72.410 ;
        RECT 73.990 72.090 74.310 72.410 ;
        RECT 108.670 72.090 108.990 72.410 ;
        RECT 109.110 72.090 109.430 72.410 ;
        RECT 109.550 72.090 109.870 72.410 ;
        RECT 109.990 72.090 110.310 72.410 ;
        RECT 144.670 72.090 144.990 72.410 ;
        RECT 145.110 72.090 145.430 72.410 ;
        RECT 145.550 72.090 145.870 72.410 ;
        RECT 145.990 72.090 146.310 72.410 ;
        RECT 0.670 59.340 0.990 59.660 ;
        RECT 1.110 59.340 1.430 59.660 ;
        RECT 1.550 59.340 1.870 59.660 ;
        RECT 1.990 59.340 2.310 59.660 ;
        RECT 180.670 59.340 180.990 59.660 ;
        RECT 181.110 59.340 181.430 59.660 ;
        RECT 181.550 59.340 181.870 59.660 ;
        RECT 181.990 59.340 182.310 59.660 ;
        RECT 36.670 30.090 36.990 30.410 ;
        RECT 37.110 30.090 37.430 30.410 ;
        RECT 37.550 30.090 37.870 30.410 ;
        RECT 37.990 30.090 38.310 30.410 ;
        RECT 72.670 30.090 72.990 30.410 ;
        RECT 73.110 30.090 73.430 30.410 ;
        RECT 73.550 30.090 73.870 30.410 ;
        RECT 73.990 30.090 74.310 30.410 ;
        RECT 108.670 30.090 108.990 30.410 ;
        RECT 109.110 30.090 109.430 30.410 ;
        RECT 109.550 30.090 109.870 30.410 ;
        RECT 109.990 30.090 110.310 30.410 ;
        RECT 144.670 30.090 144.990 30.410 ;
        RECT 145.110 30.090 145.430 30.410 ;
        RECT 145.550 30.090 145.870 30.410 ;
        RECT 145.990 30.090 146.310 30.410 ;
      LAYER met3 ;
        RECT 0.490 98.000 182.490 100.000 ;
        RECT 36.490 72.000 38.490 72.500 ;
        RECT 72.490 72.000 74.490 72.500 ;
        RECT 108.490 72.000 110.490 72.500 ;
        RECT 144.490 72.000 146.490 72.500 ;
        RECT 0.490 59.260 2.490 59.740 ;
        RECT 180.490 59.260 182.490 59.740 ;
        RECT 36.490 30.000 38.490 30.500 ;
        RECT 72.490 30.000 74.490 30.500 ;
        RECT 108.490 30.000 110.490 30.500 ;
        RECT 144.490 30.000 146.490 30.500 ;
        RECT 0.490 3.000 182.490 5.000 ;
      LAYER via3 ;
        RECT 0.690 99.400 1.090 99.800 ;
        RECT 1.290 99.400 1.690 99.800 ;
        RECT 1.890 99.400 2.290 99.800 ;
        RECT 36.690 99.400 37.090 99.800 ;
        RECT 37.290 99.400 37.690 99.800 ;
        RECT 37.890 99.400 38.290 99.800 ;
        RECT 72.690 99.400 73.090 99.800 ;
        RECT 73.290 99.400 73.690 99.800 ;
        RECT 73.890 99.400 74.290 99.800 ;
        RECT 108.690 99.400 109.090 99.800 ;
        RECT 109.290 99.400 109.690 99.800 ;
        RECT 109.890 99.400 110.290 99.800 ;
        RECT 144.690 99.400 145.090 99.800 ;
        RECT 145.290 99.400 145.690 99.800 ;
        RECT 145.890 99.400 146.290 99.800 ;
        RECT 180.690 99.400 181.090 99.800 ;
        RECT 181.290 99.400 181.690 99.800 ;
        RECT 181.890 99.400 182.290 99.800 ;
        RECT 0.690 98.800 1.090 99.200 ;
        RECT 1.290 98.800 1.690 99.200 ;
        RECT 1.890 98.800 2.290 99.200 ;
        RECT 36.690 98.800 37.090 99.200 ;
        RECT 37.290 98.800 37.690 99.200 ;
        RECT 37.890 98.800 38.290 99.200 ;
        RECT 72.690 98.800 73.090 99.200 ;
        RECT 73.290 98.800 73.690 99.200 ;
        RECT 73.890 98.800 74.290 99.200 ;
        RECT 108.690 98.800 109.090 99.200 ;
        RECT 109.290 98.800 109.690 99.200 ;
        RECT 109.890 98.800 110.290 99.200 ;
        RECT 144.690 98.800 145.090 99.200 ;
        RECT 145.290 98.800 145.690 99.200 ;
        RECT 145.890 98.800 146.290 99.200 ;
        RECT 180.690 98.800 181.090 99.200 ;
        RECT 181.290 98.800 181.690 99.200 ;
        RECT 181.890 98.800 182.290 99.200 ;
        RECT 0.690 98.200 1.090 98.600 ;
        RECT 1.290 98.200 1.690 98.600 ;
        RECT 1.890 98.200 2.290 98.600 ;
        RECT 36.690 98.200 37.090 98.600 ;
        RECT 37.290 98.200 37.690 98.600 ;
        RECT 37.890 98.200 38.290 98.600 ;
        RECT 72.690 98.200 73.090 98.600 ;
        RECT 73.290 98.200 73.690 98.600 ;
        RECT 73.890 98.200 74.290 98.600 ;
        RECT 108.690 98.200 109.090 98.600 ;
        RECT 109.290 98.200 109.690 98.600 ;
        RECT 109.890 98.200 110.290 98.600 ;
        RECT 144.690 98.200 145.090 98.600 ;
        RECT 145.290 98.200 145.690 98.600 ;
        RECT 145.890 98.200 146.290 98.600 ;
        RECT 180.690 98.200 181.090 98.600 ;
        RECT 181.290 98.200 181.690 98.600 ;
        RECT 181.890 98.200 182.290 98.600 ;
        RECT 36.650 72.070 37.010 72.435 ;
        RECT 37.090 72.070 37.450 72.435 ;
        RECT 37.530 72.070 37.890 72.435 ;
        RECT 37.970 72.070 38.330 72.435 ;
        RECT 72.650 72.070 73.010 72.435 ;
        RECT 73.090 72.070 73.450 72.435 ;
        RECT 73.530 72.070 73.890 72.435 ;
        RECT 73.970 72.070 74.330 72.435 ;
        RECT 108.650 72.070 109.010 72.435 ;
        RECT 109.090 72.070 109.450 72.435 ;
        RECT 109.530 72.070 109.890 72.435 ;
        RECT 109.970 72.070 110.330 72.435 ;
        RECT 144.650 72.070 145.010 72.435 ;
        RECT 145.090 72.070 145.450 72.435 ;
        RECT 145.530 72.070 145.890 72.435 ;
        RECT 145.970 72.070 146.330 72.435 ;
        RECT 0.650 59.320 1.010 59.685 ;
        RECT 1.090 59.320 1.450 59.685 ;
        RECT 1.530 59.320 1.890 59.685 ;
        RECT 1.970 59.320 2.330 59.685 ;
        RECT 180.650 59.320 181.010 59.685 ;
        RECT 181.090 59.320 181.450 59.685 ;
        RECT 181.530 59.320 181.890 59.685 ;
        RECT 181.970 59.320 182.330 59.685 ;
        RECT 36.650 30.070 37.010 30.435 ;
        RECT 37.090 30.070 37.450 30.435 ;
        RECT 37.530 30.070 37.890 30.435 ;
        RECT 37.970 30.070 38.330 30.435 ;
        RECT 72.650 30.070 73.010 30.435 ;
        RECT 73.090 30.070 73.450 30.435 ;
        RECT 73.530 30.070 73.890 30.435 ;
        RECT 73.970 30.070 74.330 30.435 ;
        RECT 108.650 30.070 109.010 30.435 ;
        RECT 109.090 30.070 109.450 30.435 ;
        RECT 109.530 30.070 109.890 30.435 ;
        RECT 109.970 30.070 110.330 30.435 ;
        RECT 144.650 30.070 145.010 30.435 ;
        RECT 145.090 30.070 145.450 30.435 ;
        RECT 145.530 30.070 145.890 30.435 ;
        RECT 145.970 30.070 146.330 30.435 ;
        RECT 0.690 4.400 1.090 4.800 ;
        RECT 1.290 4.400 1.690 4.800 ;
        RECT 1.890 4.400 2.290 4.800 ;
        RECT 36.690 4.400 37.090 4.800 ;
        RECT 37.290 4.400 37.690 4.800 ;
        RECT 37.890 4.400 38.290 4.800 ;
        RECT 72.690 4.400 73.090 4.800 ;
        RECT 73.290 4.400 73.690 4.800 ;
        RECT 73.890 4.400 74.290 4.800 ;
        RECT 108.690 4.400 109.090 4.800 ;
        RECT 109.290 4.400 109.690 4.800 ;
        RECT 109.890 4.400 110.290 4.800 ;
        RECT 144.690 4.400 145.090 4.800 ;
        RECT 145.290 4.400 145.690 4.800 ;
        RECT 145.890 4.400 146.290 4.800 ;
        RECT 180.690 4.400 181.090 4.800 ;
        RECT 181.290 4.400 181.690 4.800 ;
        RECT 181.890 4.400 182.290 4.800 ;
        RECT 0.690 3.800 1.090 4.200 ;
        RECT 1.290 3.800 1.690 4.200 ;
        RECT 1.890 3.800 2.290 4.200 ;
        RECT 36.690 3.800 37.090 4.200 ;
        RECT 37.290 3.800 37.690 4.200 ;
        RECT 37.890 3.800 38.290 4.200 ;
        RECT 72.690 3.800 73.090 4.200 ;
        RECT 73.290 3.800 73.690 4.200 ;
        RECT 73.890 3.800 74.290 4.200 ;
        RECT 108.690 3.800 109.090 4.200 ;
        RECT 109.290 3.800 109.690 4.200 ;
        RECT 109.890 3.800 110.290 4.200 ;
        RECT 144.690 3.800 145.090 4.200 ;
        RECT 145.290 3.800 145.690 4.200 ;
        RECT 145.890 3.800 146.290 4.200 ;
        RECT 180.690 3.800 181.090 4.200 ;
        RECT 181.290 3.800 181.690 4.200 ;
        RECT 181.890 3.800 182.290 4.200 ;
        RECT 0.690 3.200 1.090 3.600 ;
        RECT 1.290 3.200 1.690 3.600 ;
        RECT 1.890 3.200 2.290 3.600 ;
        RECT 36.690 3.200 37.090 3.600 ;
        RECT 37.290 3.200 37.690 3.600 ;
        RECT 37.890 3.200 38.290 3.600 ;
        RECT 72.690 3.200 73.090 3.600 ;
        RECT 73.290 3.200 73.690 3.600 ;
        RECT 73.890 3.200 74.290 3.600 ;
        RECT 108.690 3.200 109.090 3.600 ;
        RECT 109.290 3.200 109.690 3.600 ;
        RECT 109.890 3.200 110.290 3.600 ;
        RECT 144.690 3.200 145.090 3.600 ;
        RECT 145.290 3.200 145.690 3.600 ;
        RECT 145.890 3.200 146.290 3.600 ;
        RECT 180.690 3.200 181.090 3.600 ;
        RECT 181.290 3.200 181.690 3.600 ;
        RECT 181.890 3.200 182.290 3.600 ;
      LAYER met4 ;
        RECT 0.490 3.000 2.490 100.000 ;
        RECT 36.490 3.000 38.490 100.000 ;
        RECT 72.490 3.000 74.490 100.000 ;
        RECT 108.490 3.000 110.490 100.000 ;
        RECT 144.490 3.000 146.490 100.000 ;
        RECT 180.490 3.000 182.490 100.000 ;
    END
  END vssd2
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER li1 ;
        RECT 3.905 60.495 4.365 61.225 ;
    END
  END enb
  OBS
      LAYER pwell ;
        RECT 18.390 64.610 28.420 70.670 ;
        RECT 36.365 64.570 42.215 70.670 ;
        RECT 47.890 64.610 57.920 70.670 ;
        RECT 65.865 64.570 71.715 70.670 ;
        RECT 77.390 64.610 87.420 70.670 ;
        RECT 95.365 64.570 101.215 70.670 ;
        RECT 106.890 64.610 116.920 70.670 ;
        RECT 124.865 64.570 130.715 70.670 ;
        RECT 136.390 64.610 146.420 70.670 ;
        RECT 154.365 64.570 160.215 70.670 ;
        RECT 4.310 60.285 6.115 60.515 ;
        RECT 3.825 59.605 6.115 60.285 ;
        RECT 3.970 59.415 4.140 59.605 ;
        RECT 8.135 59.415 8.305 59.585 ;
        RECT 25.040 53.760 35.070 60.160 ;
        RECT 40.745 58.925 46.595 59.865 ;
        RECT 40.745 58.875 46.600 58.925 ;
        RECT 40.750 53.765 46.600 58.875 ;
        RECT 54.540 53.760 64.570 60.160 ;
        RECT 70.245 58.925 76.095 59.865 ;
        RECT 70.245 58.875 76.100 58.925 ;
        RECT 70.250 53.765 76.100 58.875 ;
        RECT 84.040 53.760 94.070 60.160 ;
        RECT 99.745 58.925 105.595 59.865 ;
        RECT 99.745 58.875 105.600 58.925 ;
        RECT 99.750 53.765 105.600 58.875 ;
        RECT 113.540 53.760 123.570 60.160 ;
        RECT 129.245 58.925 135.095 59.865 ;
        RECT 129.245 58.875 135.100 58.925 ;
        RECT 129.250 53.765 135.100 58.875 ;
        RECT 143.040 53.760 153.070 60.160 ;
        RECT 158.745 58.925 164.595 59.865 ;
        RECT 158.745 58.875 164.600 58.925 ;
        RECT 158.750 53.765 164.600 58.875 ;
        RECT 171.590 52.580 178.380 59.580 ;
        RECT 2.790 43.805 8.640 48.915 ;
        RECT 2.790 43.755 8.645 43.805 ;
        RECT 2.795 42.815 8.645 43.755 ;
        RECT 14.320 42.520 24.350 48.920 ;
        RECT 32.290 43.805 38.140 48.915 ;
        RECT 32.290 43.755 38.145 43.805 ;
        RECT 32.295 42.815 38.145 43.755 ;
        RECT 43.820 42.520 53.850 48.920 ;
        RECT 61.790 43.805 67.640 48.915 ;
        RECT 61.790 43.755 67.645 43.805 ;
        RECT 61.795 42.815 67.645 43.755 ;
        RECT 73.320 42.520 83.350 48.920 ;
        RECT 91.290 43.805 97.140 48.915 ;
        RECT 91.290 43.755 97.145 43.805 ;
        RECT 91.295 42.815 97.145 43.755 ;
        RECT 102.820 42.520 112.850 48.920 ;
        RECT 120.790 43.805 126.640 48.915 ;
        RECT 120.790 43.755 126.645 43.805 ;
        RECT 120.795 42.815 126.645 43.755 ;
        RECT 132.320 42.520 142.350 48.920 ;
        RECT 150.290 43.805 156.140 48.915 ;
        RECT 150.290 43.755 156.145 43.805 ;
        RECT 150.295 42.815 156.145 43.755 ;
        RECT 161.820 42.520 171.850 48.920 ;
        RECT 7.175 32.010 13.025 38.110 ;
        RECT 20.970 32.010 31.000 38.070 ;
        RECT 36.675 32.010 42.525 38.110 ;
        RECT 50.470 32.010 60.500 38.070 ;
        RECT 66.175 32.010 72.025 38.110 ;
        RECT 79.970 32.010 90.000 38.070 ;
        RECT 95.675 32.010 101.525 38.110 ;
        RECT 109.470 32.010 119.500 38.070 ;
        RECT 125.175 32.010 131.025 38.110 ;
        RECT 138.970 32.010 149.000 38.070 ;
        RECT 154.675 32.010 160.525 38.110 ;
        RECT 168.470 32.010 178.500 38.070 ;
      LAYER li1 ;
        RECT 18.570 70.140 20.915 70.620 ;
        RECT 21.980 70.140 24.840 70.620 ;
        RECT 25.895 70.140 28.240 70.620 ;
        RECT 36.545 70.140 38.890 70.620 ;
        RECT 39.690 70.140 42.035 70.620 ;
        RECT 48.070 70.140 50.415 70.620 ;
        RECT 51.480 70.140 54.340 70.620 ;
        RECT 55.395 70.140 57.740 70.620 ;
        RECT 66.045 70.140 68.390 70.620 ;
        RECT 69.190 70.140 71.535 70.620 ;
        RECT 77.570 70.140 79.915 70.620 ;
        RECT 80.980 70.140 83.840 70.620 ;
        RECT 84.895 70.140 87.240 70.620 ;
        RECT 95.545 70.140 97.890 70.620 ;
        RECT 98.690 70.140 101.035 70.620 ;
        RECT 107.070 70.140 109.415 70.620 ;
        RECT 110.480 70.140 113.340 70.620 ;
        RECT 114.395 70.140 116.740 70.620 ;
        RECT 125.045 70.140 127.390 70.620 ;
        RECT 128.190 70.140 130.535 70.620 ;
        RECT 136.570 70.140 138.915 70.620 ;
        RECT 139.980 70.140 142.840 70.620 ;
        RECT 143.895 70.140 146.240 70.620 ;
        RECT 154.545 70.140 156.890 70.620 ;
        RECT 157.690 70.140 160.035 70.620 ;
        RECT 19.080 65.545 19.370 70.140 ;
        RECT 19.140 65.300 19.310 65.545 ;
        RECT 19.290 63.090 20.420 64.090 ;
        RECT 21.170 63.780 21.460 69.840 ;
        RECT 23.260 65.545 23.550 70.140 ;
        RECT 23.320 65.300 23.490 65.545 ;
        RECT 25.350 63.880 25.640 69.840 ;
        RECT 27.440 65.545 27.730 70.140 ;
        RECT 37.055 65.790 37.345 70.140 ;
        RECT 41.235 65.790 41.525 70.140 ;
        RECT 27.500 65.535 27.695 65.545 ;
        RECT 27.500 65.300 27.670 65.535 ;
        RECT 37.290 63.880 38.490 64.190 ;
        RECT 43.525 63.975 43.820 67.050 ;
        RECT 48.580 65.545 48.870 70.140 ;
        RECT 48.640 65.300 48.810 65.545 ;
        RECT 25.350 63.780 26.170 63.880 ;
        RECT 21.170 63.280 26.170 63.780 ;
        RECT 3.905 61.565 4.165 61.965 ;
        RECT 3.905 61.395 5.270 61.565 ;
        RECT 6.330 61.455 7.780 61.675 ;
        RECT 4.535 60.325 5.270 61.395 ;
        RECT 5.795 61.375 7.780 61.455 ;
        RECT 5.795 61.155 6.630 61.375 ;
        RECT 7.480 61.240 7.780 61.375 ;
        RECT 5.795 60.475 6.035 61.155 ;
        RECT 7.480 60.940 8.595 61.240 ;
        RECT 3.905 60.155 5.270 60.325 ;
        RECT 3.905 59.755 4.165 60.155 ;
        RECT 8.075 59.755 8.595 60.940 ;
        RECT 8.765 60.415 9.285 61.965 ;
        RECT 21.170 57.330 21.460 63.280 ;
        RECT 36.790 63.260 38.490 63.880 ;
        RECT 37.290 63.060 38.490 63.260 ;
        RECT 43.295 63.195 44.035 63.975 ;
        RECT 25.790 58.895 25.960 59.130 ;
        RECT 25.765 58.885 25.960 58.895 ;
        RECT 29.970 58.885 30.140 59.110 ;
        RECT 34.150 58.885 34.320 59.110 ;
        RECT 25.730 54.300 26.020 58.885 ;
        RECT 29.910 54.300 30.200 58.885 ;
        RECT 34.090 54.300 34.380 58.885 ;
        RECT 41.440 54.300 41.730 58.645 ;
        RECT 43.525 54.605 43.820 63.195 ;
        RECT 48.790 63.090 49.920 64.090 ;
        RECT 50.670 63.780 50.960 69.840 ;
        RECT 52.760 65.545 53.050 70.140 ;
        RECT 52.820 65.300 52.990 65.545 ;
        RECT 54.850 63.880 55.140 69.840 ;
        RECT 56.940 65.545 57.230 70.140 ;
        RECT 66.555 65.790 66.845 70.140 ;
        RECT 70.735 65.790 71.025 70.140 ;
        RECT 57.000 65.535 57.195 65.545 ;
        RECT 57.000 65.300 57.170 65.535 ;
        RECT 66.790 63.880 67.990 64.190 ;
        RECT 73.025 63.975 73.320 67.050 ;
        RECT 78.080 65.545 78.370 70.140 ;
        RECT 78.140 65.300 78.310 65.545 ;
        RECT 54.850 63.780 55.670 63.880 ;
        RECT 50.670 63.280 55.670 63.780 ;
        RECT 45.620 54.300 45.910 58.645 ;
        RECT 50.670 57.330 50.960 63.280 ;
        RECT 66.290 63.260 67.990 63.880 ;
        RECT 66.790 63.060 67.990 63.260 ;
        RECT 72.795 63.195 73.535 63.975 ;
        RECT 55.290 58.895 55.460 59.130 ;
        RECT 55.265 58.885 55.460 58.895 ;
        RECT 59.470 58.885 59.640 59.110 ;
        RECT 63.650 58.885 63.820 59.110 ;
        RECT 55.230 54.300 55.520 58.885 ;
        RECT 59.410 54.300 59.700 58.885 ;
        RECT 63.590 54.300 63.880 58.885 ;
        RECT 70.940 54.300 71.230 58.645 ;
        RECT 73.025 54.605 73.320 63.195 ;
        RECT 78.290 63.090 79.420 64.090 ;
        RECT 80.170 63.780 80.460 69.840 ;
        RECT 82.260 65.545 82.550 70.140 ;
        RECT 82.320 65.300 82.490 65.545 ;
        RECT 84.350 63.880 84.640 69.840 ;
        RECT 86.440 65.545 86.730 70.140 ;
        RECT 96.055 65.790 96.345 70.140 ;
        RECT 100.235 65.790 100.525 70.140 ;
        RECT 86.500 65.535 86.695 65.545 ;
        RECT 86.500 65.300 86.670 65.535 ;
        RECT 96.290 63.880 97.490 64.190 ;
        RECT 102.525 63.975 102.820 67.050 ;
        RECT 107.580 65.545 107.870 70.140 ;
        RECT 107.640 65.300 107.810 65.545 ;
        RECT 84.350 63.780 85.170 63.880 ;
        RECT 80.170 63.280 85.170 63.780 ;
        RECT 75.120 54.300 75.410 58.645 ;
        RECT 80.170 57.330 80.460 63.280 ;
        RECT 95.790 63.260 97.490 63.880 ;
        RECT 96.290 63.060 97.490 63.260 ;
        RECT 102.295 63.195 103.035 63.975 ;
        RECT 84.790 58.895 84.960 59.130 ;
        RECT 84.765 58.885 84.960 58.895 ;
        RECT 88.970 58.885 89.140 59.110 ;
        RECT 93.150 58.885 93.320 59.110 ;
        RECT 84.730 54.300 85.020 58.885 ;
        RECT 88.910 54.300 89.200 58.885 ;
        RECT 93.090 54.300 93.380 58.885 ;
        RECT 100.440 54.300 100.730 58.645 ;
        RECT 102.525 54.605 102.820 63.195 ;
        RECT 107.790 63.090 108.920 64.090 ;
        RECT 109.670 63.780 109.960 69.840 ;
        RECT 111.760 65.545 112.050 70.140 ;
        RECT 111.820 65.300 111.990 65.545 ;
        RECT 113.850 63.880 114.140 69.840 ;
        RECT 115.940 65.545 116.230 70.140 ;
        RECT 125.555 65.790 125.845 70.140 ;
        RECT 129.735 65.790 130.025 70.140 ;
        RECT 116.000 65.535 116.195 65.545 ;
        RECT 116.000 65.300 116.170 65.535 ;
        RECT 125.790 63.880 126.990 64.190 ;
        RECT 132.025 63.975 132.320 67.050 ;
        RECT 137.080 65.545 137.370 70.140 ;
        RECT 137.140 65.300 137.310 65.545 ;
        RECT 113.850 63.780 114.670 63.880 ;
        RECT 109.670 63.280 114.670 63.780 ;
        RECT 104.620 54.300 104.910 58.645 ;
        RECT 109.670 57.330 109.960 63.280 ;
        RECT 125.290 63.260 126.990 63.880 ;
        RECT 125.790 63.060 126.990 63.260 ;
        RECT 131.795 63.195 132.535 63.975 ;
        RECT 114.290 58.895 114.460 59.130 ;
        RECT 114.265 58.885 114.460 58.895 ;
        RECT 118.470 58.885 118.640 59.110 ;
        RECT 122.650 58.885 122.820 59.110 ;
        RECT 114.230 54.300 114.520 58.885 ;
        RECT 118.410 54.300 118.700 58.885 ;
        RECT 122.590 54.300 122.880 58.885 ;
        RECT 129.940 54.300 130.230 58.645 ;
        RECT 132.025 54.605 132.320 63.195 ;
        RECT 137.290 63.090 138.420 64.090 ;
        RECT 139.170 63.780 139.460 69.840 ;
        RECT 141.260 65.545 141.550 70.140 ;
        RECT 141.320 65.300 141.490 65.545 ;
        RECT 143.350 63.880 143.640 69.840 ;
        RECT 145.440 65.545 145.730 70.140 ;
        RECT 155.055 65.790 155.345 70.140 ;
        RECT 159.235 65.790 159.525 70.140 ;
        RECT 145.500 65.535 145.695 65.545 ;
        RECT 145.500 65.300 145.670 65.535 ;
        RECT 155.290 63.880 156.490 64.190 ;
        RECT 161.525 63.975 161.820 67.050 ;
        RECT 143.350 63.780 144.170 63.880 ;
        RECT 139.170 63.280 144.170 63.780 ;
        RECT 134.120 54.300 134.410 58.645 ;
        RECT 139.170 57.330 139.460 63.280 ;
        RECT 154.790 63.260 156.490 63.880 ;
        RECT 155.290 63.060 156.490 63.260 ;
        RECT 161.295 63.195 162.035 63.975 ;
        RECT 143.790 58.895 143.960 59.130 ;
        RECT 143.765 58.885 143.960 58.895 ;
        RECT 147.970 58.885 148.140 59.110 ;
        RECT 152.150 58.885 152.320 59.110 ;
        RECT 143.730 54.300 144.020 58.885 ;
        RECT 147.910 54.300 148.200 58.885 ;
        RECT 152.090 54.300 152.380 58.885 ;
        RECT 159.440 54.300 159.730 58.645 ;
        RECT 161.525 54.605 161.820 63.195 ;
        RECT 163.620 54.300 163.910 58.645 ;
        RECT 25.220 53.820 27.570 54.300 ;
        RECT 28.620 53.820 31.480 54.300 ;
        RECT 32.545 53.820 34.890 54.300 ;
        RECT 40.930 54.270 43.270 54.300 ;
        RECT 44.080 54.270 46.420 54.300 ;
        RECT 40.930 53.850 43.275 54.270 ;
        RECT 44.075 53.850 46.420 54.270 ;
        RECT 40.930 53.820 43.270 53.850 ;
        RECT 44.080 53.820 46.420 53.850 ;
        RECT 54.720 53.820 57.070 54.300 ;
        RECT 58.120 53.820 60.980 54.300 ;
        RECT 62.045 53.820 64.390 54.300 ;
        RECT 70.430 54.270 72.770 54.300 ;
        RECT 73.580 54.270 75.920 54.300 ;
        RECT 70.430 53.850 72.775 54.270 ;
        RECT 73.575 53.850 75.920 54.270 ;
        RECT 70.430 53.820 72.770 53.850 ;
        RECT 73.580 53.820 75.920 53.850 ;
        RECT 84.220 53.820 86.570 54.300 ;
        RECT 87.620 53.820 90.480 54.300 ;
        RECT 91.545 53.820 93.890 54.300 ;
        RECT 99.930 54.270 102.270 54.300 ;
        RECT 103.080 54.270 105.420 54.300 ;
        RECT 99.930 53.850 102.275 54.270 ;
        RECT 103.075 53.850 105.420 54.270 ;
        RECT 99.930 53.820 102.270 53.850 ;
        RECT 103.080 53.820 105.420 53.850 ;
        RECT 113.720 53.820 116.070 54.300 ;
        RECT 117.120 53.820 119.980 54.300 ;
        RECT 121.045 53.820 123.390 54.300 ;
        RECT 129.430 54.270 131.770 54.300 ;
        RECT 132.580 54.270 134.920 54.300 ;
        RECT 129.430 53.850 131.775 54.270 ;
        RECT 132.575 53.850 134.920 54.270 ;
        RECT 129.430 53.820 131.770 53.850 ;
        RECT 132.580 53.820 134.920 53.850 ;
        RECT 143.220 53.820 145.570 54.300 ;
        RECT 146.620 53.820 149.480 54.300 ;
        RECT 150.545 53.820 152.890 54.300 ;
        RECT 158.930 54.270 161.270 54.300 ;
        RECT 162.080 54.270 164.420 54.300 ;
        RECT 158.930 53.850 161.275 54.270 ;
        RECT 162.075 53.850 164.420 54.270 ;
        RECT 172.500 54.120 174.340 54.150 ;
        RECT 172.420 53.950 174.420 54.120 ;
        RECT 158.930 53.820 161.270 53.850 ;
        RECT 162.080 53.820 164.420 53.850 ;
        RECT 175.630 53.660 177.470 53.690 ;
        RECT 175.550 53.490 177.550 53.660 ;
        RECT 2.970 48.830 5.310 48.860 ;
        RECT 6.120 48.830 8.460 48.860 ;
        RECT 2.970 48.410 5.315 48.830 ;
        RECT 6.115 48.410 8.460 48.830 ;
        RECT 2.970 48.380 5.310 48.410 ;
        RECT 6.120 48.380 8.460 48.410 ;
        RECT 14.500 48.380 16.845 48.860 ;
        RECT 17.910 48.380 20.770 48.860 ;
        RECT 21.820 48.380 24.170 48.860 ;
        RECT 32.470 48.830 34.810 48.860 ;
        RECT 35.620 48.830 37.960 48.860 ;
        RECT 32.470 48.410 34.815 48.830 ;
        RECT 35.615 48.410 37.960 48.830 ;
        RECT 32.470 48.380 34.810 48.410 ;
        RECT 35.620 48.380 37.960 48.410 ;
        RECT 44.000 48.380 46.345 48.860 ;
        RECT 47.410 48.380 50.270 48.860 ;
        RECT 51.320 48.380 53.670 48.860 ;
        RECT 61.970 48.830 64.310 48.860 ;
        RECT 65.120 48.830 67.460 48.860 ;
        RECT 61.970 48.410 64.315 48.830 ;
        RECT 65.115 48.410 67.460 48.830 ;
        RECT 61.970 48.380 64.310 48.410 ;
        RECT 65.120 48.380 67.460 48.410 ;
        RECT 73.500 48.380 75.845 48.860 ;
        RECT 76.910 48.380 79.770 48.860 ;
        RECT 80.820 48.380 83.170 48.860 ;
        RECT 91.470 48.830 93.810 48.860 ;
        RECT 94.620 48.830 96.960 48.860 ;
        RECT 91.470 48.410 93.815 48.830 ;
        RECT 94.615 48.410 96.960 48.830 ;
        RECT 91.470 48.380 93.810 48.410 ;
        RECT 94.620 48.380 96.960 48.410 ;
        RECT 103.000 48.380 105.345 48.860 ;
        RECT 106.410 48.380 109.270 48.860 ;
        RECT 110.320 48.380 112.670 48.860 ;
        RECT 120.970 48.830 123.310 48.860 ;
        RECT 124.120 48.830 126.460 48.860 ;
        RECT 120.970 48.410 123.315 48.830 ;
        RECT 124.115 48.410 126.460 48.830 ;
        RECT 120.970 48.380 123.310 48.410 ;
        RECT 124.120 48.380 126.460 48.410 ;
        RECT 132.500 48.380 134.845 48.860 ;
        RECT 135.910 48.380 138.770 48.860 ;
        RECT 139.820 48.380 142.170 48.860 ;
        RECT 150.470 48.830 152.810 48.860 ;
        RECT 153.620 48.830 155.960 48.860 ;
        RECT 150.470 48.410 152.815 48.830 ;
        RECT 153.615 48.410 155.960 48.830 ;
        RECT 150.470 48.380 152.810 48.410 ;
        RECT 153.620 48.380 155.960 48.410 ;
        RECT 162.000 48.380 164.345 48.860 ;
        RECT 165.410 48.380 168.270 48.860 ;
        RECT 169.320 48.380 171.670 48.860 ;
        RECT 3.480 44.035 3.770 48.380 ;
        RECT 5.570 39.485 5.865 48.075 ;
        RECT 7.660 44.035 7.950 48.380 ;
        RECT 15.010 43.795 15.300 48.380 ;
        RECT 19.190 43.795 19.480 48.380 ;
        RECT 23.370 43.795 23.660 48.380 ;
        RECT 15.070 43.570 15.240 43.795 ;
        RECT 19.250 43.570 19.420 43.795 ;
        RECT 23.430 43.785 23.625 43.795 ;
        RECT 23.430 43.550 23.600 43.785 ;
        RECT 5.355 38.705 6.095 39.485 ;
        RECT 10.900 39.420 12.100 39.620 ;
        RECT 10.900 38.800 12.600 39.420 ;
        RECT 27.930 39.400 28.220 45.350 ;
        RECT 32.980 44.035 33.270 48.380 ;
        RECT 23.220 38.900 28.220 39.400 ;
        RECT 23.220 38.800 24.040 38.900 ;
        RECT 5.570 35.630 5.865 38.705 ;
        RECT 10.900 38.490 12.100 38.800 ;
        RECT 21.720 37.145 21.890 37.380 ;
        RECT 21.695 37.135 21.890 37.145 ;
        RECT 7.865 32.540 8.155 36.890 ;
        RECT 12.045 32.540 12.335 36.890 ;
        RECT 21.660 32.540 21.950 37.135 ;
        RECT 23.750 32.840 24.040 38.800 ;
        RECT 25.900 37.135 26.070 37.380 ;
        RECT 25.840 32.540 26.130 37.135 ;
        RECT 27.930 32.840 28.220 38.900 ;
        RECT 28.970 38.590 30.100 39.590 ;
        RECT 35.070 39.485 35.365 48.075 ;
        RECT 37.160 44.035 37.450 48.380 ;
        RECT 44.510 43.795 44.800 48.380 ;
        RECT 48.690 43.795 48.980 48.380 ;
        RECT 52.870 43.795 53.160 48.380 ;
        RECT 44.570 43.570 44.740 43.795 ;
        RECT 48.750 43.570 48.920 43.795 ;
        RECT 52.930 43.785 53.125 43.795 ;
        RECT 52.930 43.550 53.100 43.785 ;
        RECT 34.855 38.705 35.595 39.485 ;
        RECT 40.400 39.420 41.600 39.620 ;
        RECT 40.400 38.800 42.100 39.420 ;
        RECT 57.430 39.400 57.720 45.350 ;
        RECT 62.480 44.035 62.770 48.380 ;
        RECT 52.720 38.900 57.720 39.400 ;
        RECT 52.720 38.800 53.540 38.900 ;
        RECT 30.080 37.135 30.250 37.380 ;
        RECT 30.020 32.540 30.310 37.135 ;
        RECT 35.070 35.630 35.365 38.705 ;
        RECT 40.400 38.490 41.600 38.800 ;
        RECT 51.220 37.145 51.390 37.380 ;
        RECT 51.195 37.135 51.390 37.145 ;
        RECT 37.365 32.540 37.655 36.890 ;
        RECT 41.545 32.540 41.835 36.890 ;
        RECT 51.160 32.540 51.450 37.135 ;
        RECT 53.250 32.840 53.540 38.800 ;
        RECT 55.400 37.135 55.570 37.380 ;
        RECT 55.340 32.540 55.630 37.135 ;
        RECT 57.430 32.840 57.720 38.900 ;
        RECT 58.470 38.590 59.600 39.590 ;
        RECT 64.570 39.485 64.865 48.075 ;
        RECT 66.660 44.035 66.950 48.380 ;
        RECT 74.010 43.795 74.300 48.380 ;
        RECT 78.190 43.795 78.480 48.380 ;
        RECT 82.370 43.795 82.660 48.380 ;
        RECT 74.070 43.570 74.240 43.795 ;
        RECT 78.250 43.570 78.420 43.795 ;
        RECT 82.430 43.785 82.625 43.795 ;
        RECT 82.430 43.550 82.600 43.785 ;
        RECT 64.355 38.705 65.095 39.485 ;
        RECT 69.900 39.420 71.100 39.620 ;
        RECT 69.900 38.800 71.600 39.420 ;
        RECT 86.930 39.400 87.220 45.350 ;
        RECT 91.980 44.035 92.270 48.380 ;
        RECT 82.220 38.900 87.220 39.400 ;
        RECT 82.220 38.800 83.040 38.900 ;
        RECT 59.580 37.135 59.750 37.380 ;
        RECT 59.520 32.540 59.810 37.135 ;
        RECT 64.570 35.630 64.865 38.705 ;
        RECT 69.900 38.490 71.100 38.800 ;
        RECT 80.720 37.145 80.890 37.380 ;
        RECT 80.695 37.135 80.890 37.145 ;
        RECT 66.865 32.540 67.155 36.890 ;
        RECT 71.045 32.540 71.335 36.890 ;
        RECT 80.660 32.540 80.950 37.135 ;
        RECT 82.750 32.840 83.040 38.800 ;
        RECT 84.900 37.135 85.070 37.380 ;
        RECT 84.840 32.540 85.130 37.135 ;
        RECT 86.930 32.840 87.220 38.900 ;
        RECT 87.970 38.590 89.100 39.590 ;
        RECT 94.070 39.485 94.365 48.075 ;
        RECT 96.160 44.035 96.450 48.380 ;
        RECT 103.510 43.795 103.800 48.380 ;
        RECT 107.690 43.795 107.980 48.380 ;
        RECT 111.870 43.795 112.160 48.380 ;
        RECT 103.570 43.570 103.740 43.795 ;
        RECT 107.750 43.570 107.920 43.795 ;
        RECT 111.930 43.785 112.125 43.795 ;
        RECT 111.930 43.550 112.100 43.785 ;
        RECT 93.855 38.705 94.595 39.485 ;
        RECT 99.400 39.420 100.600 39.620 ;
        RECT 99.400 38.800 101.100 39.420 ;
        RECT 116.430 39.400 116.720 45.350 ;
        RECT 121.480 44.035 121.770 48.380 ;
        RECT 111.720 38.900 116.720 39.400 ;
        RECT 111.720 38.800 112.540 38.900 ;
        RECT 89.080 37.135 89.250 37.380 ;
        RECT 89.020 32.540 89.310 37.135 ;
        RECT 94.070 35.630 94.365 38.705 ;
        RECT 99.400 38.490 100.600 38.800 ;
        RECT 110.220 37.145 110.390 37.380 ;
        RECT 110.195 37.135 110.390 37.145 ;
        RECT 96.365 32.540 96.655 36.890 ;
        RECT 100.545 32.540 100.835 36.890 ;
        RECT 110.160 32.540 110.450 37.135 ;
        RECT 112.250 32.840 112.540 38.800 ;
        RECT 114.400 37.135 114.570 37.380 ;
        RECT 114.340 32.540 114.630 37.135 ;
        RECT 116.430 32.840 116.720 38.900 ;
        RECT 117.470 38.590 118.600 39.590 ;
        RECT 123.570 39.485 123.865 48.075 ;
        RECT 125.660 44.035 125.950 48.380 ;
        RECT 133.010 43.795 133.300 48.380 ;
        RECT 137.190 43.795 137.480 48.380 ;
        RECT 141.370 43.795 141.660 48.380 ;
        RECT 133.070 43.570 133.240 43.795 ;
        RECT 137.250 43.570 137.420 43.795 ;
        RECT 141.430 43.785 141.625 43.795 ;
        RECT 141.430 43.550 141.600 43.785 ;
        RECT 123.355 38.705 124.095 39.485 ;
        RECT 128.900 39.420 130.100 39.620 ;
        RECT 128.900 38.800 130.600 39.420 ;
        RECT 145.930 39.400 146.220 45.350 ;
        RECT 150.980 44.035 151.270 48.380 ;
        RECT 141.220 38.900 146.220 39.400 ;
        RECT 141.220 38.800 142.040 38.900 ;
        RECT 118.580 37.135 118.750 37.380 ;
        RECT 118.520 32.540 118.810 37.135 ;
        RECT 123.570 35.630 123.865 38.705 ;
        RECT 128.900 38.490 130.100 38.800 ;
        RECT 139.720 37.145 139.890 37.380 ;
        RECT 139.695 37.135 139.890 37.145 ;
        RECT 125.865 32.540 126.155 36.890 ;
        RECT 130.045 32.540 130.335 36.890 ;
        RECT 139.660 32.540 139.950 37.135 ;
        RECT 141.750 32.840 142.040 38.800 ;
        RECT 143.900 37.135 144.070 37.380 ;
        RECT 143.840 32.540 144.130 37.135 ;
        RECT 145.930 32.840 146.220 38.900 ;
        RECT 146.970 38.590 148.100 39.590 ;
        RECT 153.070 39.485 153.365 48.075 ;
        RECT 155.160 44.035 155.450 48.380 ;
        RECT 162.510 43.795 162.800 48.380 ;
        RECT 166.690 43.795 166.980 48.380 ;
        RECT 170.870 43.795 171.160 48.380 ;
        RECT 162.570 43.570 162.740 43.795 ;
        RECT 166.750 43.570 166.920 43.795 ;
        RECT 170.930 43.785 171.125 43.795 ;
        RECT 170.930 43.550 171.100 43.785 ;
        RECT 152.855 38.705 153.595 39.485 ;
        RECT 158.400 39.420 159.600 39.620 ;
        RECT 158.400 38.800 160.100 39.420 ;
        RECT 175.430 39.400 175.720 45.350 ;
        RECT 170.720 38.900 175.720 39.400 ;
        RECT 170.720 38.800 171.540 38.900 ;
        RECT 148.080 37.135 148.250 37.380 ;
        RECT 148.020 32.540 148.310 37.135 ;
        RECT 153.070 35.630 153.365 38.705 ;
        RECT 158.400 38.490 159.600 38.800 ;
        RECT 169.220 37.145 169.390 37.380 ;
        RECT 169.195 37.135 169.390 37.145 ;
        RECT 155.365 32.540 155.655 36.890 ;
        RECT 159.545 32.540 159.835 36.890 ;
        RECT 169.160 32.540 169.450 37.135 ;
        RECT 171.250 32.840 171.540 38.800 ;
        RECT 173.400 37.135 173.570 37.380 ;
        RECT 173.340 32.540 173.630 37.135 ;
        RECT 175.430 32.840 175.720 38.900 ;
        RECT 176.470 38.590 177.600 39.590 ;
        RECT 177.580 37.135 177.750 37.380 ;
        RECT 177.520 32.540 177.810 37.135 ;
        RECT 7.355 32.060 9.700 32.540 ;
        RECT 10.500 32.060 12.845 32.540 ;
        RECT 21.150 32.060 23.495 32.540 ;
        RECT 24.550 32.060 27.410 32.540 ;
        RECT 28.475 32.060 30.820 32.540 ;
        RECT 36.855 32.060 39.200 32.540 ;
        RECT 40.000 32.060 42.345 32.540 ;
        RECT 50.650 32.060 52.995 32.540 ;
        RECT 54.050 32.060 56.910 32.540 ;
        RECT 57.975 32.060 60.320 32.540 ;
        RECT 66.355 32.060 68.700 32.540 ;
        RECT 69.500 32.060 71.845 32.540 ;
        RECT 80.150 32.060 82.495 32.540 ;
        RECT 83.550 32.060 86.410 32.540 ;
        RECT 87.475 32.060 89.820 32.540 ;
        RECT 95.855 32.060 98.200 32.540 ;
        RECT 99.000 32.060 101.345 32.540 ;
        RECT 109.650 32.060 111.995 32.540 ;
        RECT 113.050 32.060 115.910 32.540 ;
        RECT 116.975 32.060 119.320 32.540 ;
        RECT 125.355 32.060 127.700 32.540 ;
        RECT 128.500 32.060 130.845 32.540 ;
        RECT 139.150 32.060 141.495 32.540 ;
        RECT 142.550 32.060 145.410 32.540 ;
        RECT 146.475 32.060 148.820 32.540 ;
        RECT 154.855 32.060 157.200 32.540 ;
        RECT 158.000 32.060 160.345 32.540 ;
        RECT 168.650 32.060 170.995 32.540 ;
        RECT 172.050 32.060 174.910 32.540 ;
        RECT 175.975 32.060 178.320 32.540 ;
      LAYER mcon ;
        RECT 18.570 70.170 19.085 70.590 ;
        RECT 19.275 70.170 19.695 70.590 ;
        RECT 19.885 70.170 20.305 70.590 ;
        RECT 20.495 70.170 20.915 70.590 ;
        RECT 21.980 70.170 22.400 70.590 ;
        RECT 22.590 70.170 23.010 70.590 ;
        RECT 23.200 70.170 23.620 70.590 ;
        RECT 23.810 70.170 24.230 70.590 ;
        RECT 24.420 70.170 24.840 70.590 ;
        RECT 25.895 70.170 26.315 70.590 ;
        RECT 26.505 70.170 26.925 70.590 ;
        RECT 27.115 70.170 27.535 70.590 ;
        RECT 27.725 70.170 28.240 70.590 ;
        RECT 36.545 70.170 36.965 70.590 ;
        RECT 37.155 70.170 37.575 70.590 ;
        RECT 37.765 70.170 38.185 70.590 ;
        RECT 38.375 70.170 38.890 70.590 ;
        RECT 39.690 70.170 40.205 70.590 ;
        RECT 40.395 70.170 40.815 70.590 ;
        RECT 41.005 70.170 41.425 70.590 ;
        RECT 41.615 70.170 42.035 70.590 ;
        RECT 48.070 70.170 48.585 70.590 ;
        RECT 48.775 70.170 49.195 70.590 ;
        RECT 49.385 70.170 49.805 70.590 ;
        RECT 49.995 70.170 50.415 70.590 ;
        RECT 51.480 70.170 51.900 70.590 ;
        RECT 52.090 70.170 52.510 70.590 ;
        RECT 52.700 70.170 53.120 70.590 ;
        RECT 53.310 70.170 53.730 70.590 ;
        RECT 53.920 70.170 54.340 70.590 ;
        RECT 55.395 70.170 55.815 70.590 ;
        RECT 56.005 70.170 56.425 70.590 ;
        RECT 56.615 70.170 57.035 70.590 ;
        RECT 57.225 70.170 57.740 70.590 ;
        RECT 66.045 70.170 66.465 70.590 ;
        RECT 66.655 70.170 67.075 70.590 ;
        RECT 67.265 70.170 67.685 70.590 ;
        RECT 67.875 70.170 68.390 70.590 ;
        RECT 69.190 70.170 69.705 70.590 ;
        RECT 69.895 70.170 70.315 70.590 ;
        RECT 70.505 70.170 70.925 70.590 ;
        RECT 71.115 70.170 71.535 70.590 ;
        RECT 77.570 70.170 78.085 70.590 ;
        RECT 78.275 70.170 78.695 70.590 ;
        RECT 78.885 70.170 79.305 70.590 ;
        RECT 79.495 70.170 79.915 70.590 ;
        RECT 80.980 70.170 81.400 70.590 ;
        RECT 81.590 70.170 82.010 70.590 ;
        RECT 82.200 70.170 82.620 70.590 ;
        RECT 82.810 70.170 83.230 70.590 ;
        RECT 83.420 70.170 83.840 70.590 ;
        RECT 84.895 70.170 85.315 70.590 ;
        RECT 85.505 70.170 85.925 70.590 ;
        RECT 86.115 70.170 86.535 70.590 ;
        RECT 86.725 70.170 87.240 70.590 ;
        RECT 95.545 70.170 95.965 70.590 ;
        RECT 96.155 70.170 96.575 70.590 ;
        RECT 96.765 70.170 97.185 70.590 ;
        RECT 97.375 70.170 97.890 70.590 ;
        RECT 98.690 70.170 99.205 70.590 ;
        RECT 99.395 70.170 99.815 70.590 ;
        RECT 100.005 70.170 100.425 70.590 ;
        RECT 100.615 70.170 101.035 70.590 ;
        RECT 107.070 70.170 107.585 70.590 ;
        RECT 107.775 70.170 108.195 70.590 ;
        RECT 108.385 70.170 108.805 70.590 ;
        RECT 108.995 70.170 109.415 70.590 ;
        RECT 110.480 70.170 110.900 70.590 ;
        RECT 111.090 70.170 111.510 70.590 ;
        RECT 111.700 70.170 112.120 70.590 ;
        RECT 112.310 70.170 112.730 70.590 ;
        RECT 112.920 70.170 113.340 70.590 ;
        RECT 114.395 70.170 114.815 70.590 ;
        RECT 115.005 70.170 115.425 70.590 ;
        RECT 115.615 70.170 116.035 70.590 ;
        RECT 116.225 70.170 116.740 70.590 ;
        RECT 125.045 70.170 125.465 70.590 ;
        RECT 125.655 70.170 126.075 70.590 ;
        RECT 126.265 70.170 126.685 70.590 ;
        RECT 126.875 70.170 127.390 70.590 ;
        RECT 128.190 70.170 128.705 70.590 ;
        RECT 128.895 70.170 129.315 70.590 ;
        RECT 129.505 70.170 129.925 70.590 ;
        RECT 130.115 70.170 130.535 70.590 ;
        RECT 136.570 70.170 137.085 70.590 ;
        RECT 137.275 70.170 137.695 70.590 ;
        RECT 137.885 70.170 138.305 70.590 ;
        RECT 138.495 70.170 138.915 70.590 ;
        RECT 139.980 70.170 140.400 70.590 ;
        RECT 140.590 70.170 141.010 70.590 ;
        RECT 141.200 70.170 141.620 70.590 ;
        RECT 141.810 70.170 142.230 70.590 ;
        RECT 142.420 70.170 142.840 70.590 ;
        RECT 143.895 70.170 144.315 70.590 ;
        RECT 144.505 70.170 144.925 70.590 ;
        RECT 145.115 70.170 145.535 70.590 ;
        RECT 145.725 70.170 146.240 70.590 ;
        RECT 154.545 70.170 154.965 70.590 ;
        RECT 155.155 70.170 155.575 70.590 ;
        RECT 155.765 70.170 156.185 70.590 ;
        RECT 156.375 70.170 156.890 70.590 ;
        RECT 157.690 70.170 158.205 70.590 ;
        RECT 158.395 70.170 158.815 70.590 ;
        RECT 159.005 70.170 159.425 70.590 ;
        RECT 159.615 70.170 160.035 70.590 ;
        RECT 19.320 63.120 20.330 64.060 ;
        RECT 25.350 63.280 26.170 63.880 ;
        RECT 36.820 63.290 37.270 63.880 ;
        RECT 37.460 63.290 38.490 63.880 ;
        RECT 43.355 63.225 43.975 63.945 ;
        RECT 48.820 63.120 49.830 64.060 ;
        RECT 54.850 63.280 55.670 63.880 ;
        RECT 66.320 63.290 66.770 63.880 ;
        RECT 66.960 63.290 67.990 63.880 ;
        RECT 72.855 63.225 73.475 63.945 ;
        RECT 78.320 63.120 79.330 64.060 ;
        RECT 84.350 63.280 85.170 63.880 ;
        RECT 95.820 63.290 96.270 63.880 ;
        RECT 96.460 63.290 97.490 63.880 ;
        RECT 102.355 63.225 102.975 63.945 ;
        RECT 107.820 63.120 108.830 64.060 ;
        RECT 113.850 63.280 114.670 63.880 ;
        RECT 125.320 63.290 125.770 63.880 ;
        RECT 125.960 63.290 126.990 63.880 ;
        RECT 131.855 63.225 132.475 63.945 ;
        RECT 137.320 63.120 138.330 64.060 ;
        RECT 143.350 63.280 144.170 63.880 ;
        RECT 154.820 63.290 155.270 63.880 ;
        RECT 155.460 63.290 156.490 63.880 ;
        RECT 161.355 63.225 161.975 63.945 ;
        RECT 25.220 53.850 25.735 54.270 ;
        RECT 25.925 53.850 26.345 54.270 ;
        RECT 26.535 53.850 26.955 54.270 ;
        RECT 27.145 53.850 27.565 54.270 ;
        RECT 28.620 53.850 29.040 54.270 ;
        RECT 29.230 53.850 29.650 54.270 ;
        RECT 29.840 53.850 30.260 54.270 ;
        RECT 30.450 53.850 30.870 54.270 ;
        RECT 31.060 53.850 31.480 54.270 ;
        RECT 32.545 53.850 32.965 54.270 ;
        RECT 33.155 53.850 33.575 54.270 ;
        RECT 33.765 53.850 34.185 54.270 ;
        RECT 34.375 53.850 34.890 54.270 ;
        RECT 41.640 53.850 42.050 54.270 ;
        RECT 42.250 53.850 42.660 54.270 ;
        RECT 42.860 53.850 43.275 54.270 ;
        RECT 44.685 53.850 45.105 54.270 ;
        RECT 45.295 53.850 45.715 54.270 ;
        RECT 45.905 53.850 46.420 54.270 ;
        RECT 54.720 53.850 55.235 54.270 ;
        RECT 55.425 53.850 55.845 54.270 ;
        RECT 56.035 53.850 56.455 54.270 ;
        RECT 56.645 53.850 57.065 54.270 ;
        RECT 58.120 53.850 58.540 54.270 ;
        RECT 58.730 53.850 59.150 54.270 ;
        RECT 59.340 53.850 59.760 54.270 ;
        RECT 59.950 53.850 60.370 54.270 ;
        RECT 60.560 53.850 60.980 54.270 ;
        RECT 62.045 53.850 62.465 54.270 ;
        RECT 62.655 53.850 63.075 54.270 ;
        RECT 63.265 53.850 63.685 54.270 ;
        RECT 63.875 53.850 64.390 54.270 ;
        RECT 71.140 53.850 71.550 54.270 ;
        RECT 71.750 53.850 72.160 54.270 ;
        RECT 72.360 53.850 72.775 54.270 ;
        RECT 74.185 53.850 74.605 54.270 ;
        RECT 74.795 53.850 75.215 54.270 ;
        RECT 75.405 53.850 75.920 54.270 ;
        RECT 84.220 53.850 84.735 54.270 ;
        RECT 84.925 53.850 85.345 54.270 ;
        RECT 85.535 53.850 85.955 54.270 ;
        RECT 86.145 53.850 86.565 54.270 ;
        RECT 87.620 53.850 88.040 54.270 ;
        RECT 88.230 53.850 88.650 54.270 ;
        RECT 88.840 53.850 89.260 54.270 ;
        RECT 89.450 53.850 89.870 54.270 ;
        RECT 90.060 53.850 90.480 54.270 ;
        RECT 91.545 53.850 91.965 54.270 ;
        RECT 92.155 53.850 92.575 54.270 ;
        RECT 92.765 53.850 93.185 54.270 ;
        RECT 93.375 53.850 93.890 54.270 ;
        RECT 100.640 53.850 101.050 54.270 ;
        RECT 101.250 53.850 101.660 54.270 ;
        RECT 101.860 53.850 102.275 54.270 ;
        RECT 103.685 53.850 104.105 54.270 ;
        RECT 104.295 53.850 104.715 54.270 ;
        RECT 104.905 53.850 105.420 54.270 ;
        RECT 113.720 53.850 114.235 54.270 ;
        RECT 114.425 53.850 114.845 54.270 ;
        RECT 115.035 53.850 115.455 54.270 ;
        RECT 115.645 53.850 116.065 54.270 ;
        RECT 117.120 53.850 117.540 54.270 ;
        RECT 117.730 53.850 118.150 54.270 ;
        RECT 118.340 53.850 118.760 54.270 ;
        RECT 118.950 53.850 119.370 54.270 ;
        RECT 119.560 53.850 119.980 54.270 ;
        RECT 121.045 53.850 121.465 54.270 ;
        RECT 121.655 53.850 122.075 54.270 ;
        RECT 122.265 53.850 122.685 54.270 ;
        RECT 122.875 53.850 123.390 54.270 ;
        RECT 130.140 53.850 130.550 54.270 ;
        RECT 130.750 53.850 131.160 54.270 ;
        RECT 131.360 53.850 131.775 54.270 ;
        RECT 133.185 53.850 133.605 54.270 ;
        RECT 133.795 53.850 134.215 54.270 ;
        RECT 134.405 53.850 134.920 54.270 ;
        RECT 143.220 53.850 143.735 54.270 ;
        RECT 143.925 53.850 144.345 54.270 ;
        RECT 144.535 53.850 144.955 54.270 ;
        RECT 145.145 53.850 145.565 54.270 ;
        RECT 146.620 53.850 147.040 54.270 ;
        RECT 147.230 53.850 147.650 54.270 ;
        RECT 147.840 53.850 148.260 54.270 ;
        RECT 148.450 53.850 148.870 54.270 ;
        RECT 149.060 53.850 149.480 54.270 ;
        RECT 150.545 53.850 150.965 54.270 ;
        RECT 151.155 53.850 151.575 54.270 ;
        RECT 151.765 53.850 152.185 54.270 ;
        RECT 152.375 53.850 152.890 54.270 ;
        RECT 159.640 53.850 160.050 54.270 ;
        RECT 160.250 53.850 160.660 54.270 ;
        RECT 160.860 53.850 161.275 54.270 ;
        RECT 162.685 53.850 163.105 54.270 ;
        RECT 163.295 53.850 163.715 54.270 ;
        RECT 163.905 53.850 164.420 54.270 ;
        RECT 172.615 53.965 172.785 54.135 ;
        RECT 172.975 53.965 173.145 54.135 ;
        RECT 173.335 53.965 173.505 54.135 ;
        RECT 173.695 53.965 173.865 54.135 ;
        RECT 174.055 53.965 174.225 54.135 ;
        RECT 175.745 53.505 175.915 53.675 ;
        RECT 176.105 53.505 176.275 53.675 ;
        RECT 176.465 53.505 176.635 53.675 ;
        RECT 176.825 53.505 176.995 53.675 ;
        RECT 177.185 53.505 177.355 53.675 ;
        RECT 3.675 48.410 4.095 48.830 ;
        RECT 4.285 48.410 4.705 48.830 ;
        RECT 4.895 48.410 5.315 48.830 ;
        RECT 6.730 48.410 7.140 48.830 ;
        RECT 7.340 48.410 7.750 48.830 ;
        RECT 7.950 48.410 8.460 48.830 ;
        RECT 14.500 48.410 15.015 48.830 ;
        RECT 15.205 48.410 15.625 48.830 ;
        RECT 15.815 48.410 16.235 48.830 ;
        RECT 16.425 48.410 16.845 48.830 ;
        RECT 17.910 48.410 18.330 48.830 ;
        RECT 18.520 48.410 18.940 48.830 ;
        RECT 19.130 48.410 19.550 48.830 ;
        RECT 19.740 48.410 20.160 48.830 ;
        RECT 20.350 48.410 20.770 48.830 ;
        RECT 21.825 48.410 22.245 48.830 ;
        RECT 22.435 48.410 22.855 48.830 ;
        RECT 23.045 48.410 23.465 48.830 ;
        RECT 23.655 48.410 24.170 48.830 ;
        RECT 33.175 48.410 33.595 48.830 ;
        RECT 33.785 48.410 34.205 48.830 ;
        RECT 34.395 48.410 34.815 48.830 ;
        RECT 36.230 48.410 36.640 48.830 ;
        RECT 36.840 48.410 37.250 48.830 ;
        RECT 37.450 48.410 37.960 48.830 ;
        RECT 44.000 48.410 44.515 48.830 ;
        RECT 44.705 48.410 45.125 48.830 ;
        RECT 45.315 48.410 45.735 48.830 ;
        RECT 45.925 48.410 46.345 48.830 ;
        RECT 47.410 48.410 47.830 48.830 ;
        RECT 48.020 48.410 48.440 48.830 ;
        RECT 48.630 48.410 49.050 48.830 ;
        RECT 49.240 48.410 49.660 48.830 ;
        RECT 49.850 48.410 50.270 48.830 ;
        RECT 51.325 48.410 51.745 48.830 ;
        RECT 51.935 48.410 52.355 48.830 ;
        RECT 52.545 48.410 52.965 48.830 ;
        RECT 53.155 48.410 53.670 48.830 ;
        RECT 62.675 48.410 63.095 48.830 ;
        RECT 63.285 48.410 63.705 48.830 ;
        RECT 63.895 48.410 64.315 48.830 ;
        RECT 65.730 48.410 66.140 48.830 ;
        RECT 66.340 48.410 66.750 48.830 ;
        RECT 66.950 48.410 67.460 48.830 ;
        RECT 73.500 48.410 74.015 48.830 ;
        RECT 74.205 48.410 74.625 48.830 ;
        RECT 74.815 48.410 75.235 48.830 ;
        RECT 75.425 48.410 75.845 48.830 ;
        RECT 76.910 48.410 77.330 48.830 ;
        RECT 77.520 48.410 77.940 48.830 ;
        RECT 78.130 48.410 78.550 48.830 ;
        RECT 78.740 48.410 79.160 48.830 ;
        RECT 79.350 48.410 79.770 48.830 ;
        RECT 80.825 48.410 81.245 48.830 ;
        RECT 81.435 48.410 81.855 48.830 ;
        RECT 82.045 48.410 82.465 48.830 ;
        RECT 82.655 48.410 83.170 48.830 ;
        RECT 92.175 48.410 92.595 48.830 ;
        RECT 92.785 48.410 93.205 48.830 ;
        RECT 93.395 48.410 93.815 48.830 ;
        RECT 95.230 48.410 95.640 48.830 ;
        RECT 95.840 48.410 96.250 48.830 ;
        RECT 96.450 48.410 96.960 48.830 ;
        RECT 103.000 48.410 103.515 48.830 ;
        RECT 103.705 48.410 104.125 48.830 ;
        RECT 104.315 48.410 104.735 48.830 ;
        RECT 104.925 48.410 105.345 48.830 ;
        RECT 106.410 48.410 106.830 48.830 ;
        RECT 107.020 48.410 107.440 48.830 ;
        RECT 107.630 48.410 108.050 48.830 ;
        RECT 108.240 48.410 108.660 48.830 ;
        RECT 108.850 48.410 109.270 48.830 ;
        RECT 110.325 48.410 110.745 48.830 ;
        RECT 110.935 48.410 111.355 48.830 ;
        RECT 111.545 48.410 111.965 48.830 ;
        RECT 112.155 48.410 112.670 48.830 ;
        RECT 121.675 48.410 122.095 48.830 ;
        RECT 122.285 48.410 122.705 48.830 ;
        RECT 122.895 48.410 123.315 48.830 ;
        RECT 124.730 48.410 125.140 48.830 ;
        RECT 125.340 48.410 125.750 48.830 ;
        RECT 125.950 48.410 126.460 48.830 ;
        RECT 132.500 48.410 133.015 48.830 ;
        RECT 133.205 48.410 133.625 48.830 ;
        RECT 133.815 48.410 134.235 48.830 ;
        RECT 134.425 48.410 134.845 48.830 ;
        RECT 135.910 48.410 136.330 48.830 ;
        RECT 136.520 48.410 136.940 48.830 ;
        RECT 137.130 48.410 137.550 48.830 ;
        RECT 137.740 48.410 138.160 48.830 ;
        RECT 138.350 48.410 138.770 48.830 ;
        RECT 139.825 48.410 140.245 48.830 ;
        RECT 140.435 48.410 140.855 48.830 ;
        RECT 141.045 48.410 141.465 48.830 ;
        RECT 141.655 48.410 142.170 48.830 ;
        RECT 151.175 48.410 151.595 48.830 ;
        RECT 151.785 48.410 152.205 48.830 ;
        RECT 152.395 48.410 152.815 48.830 ;
        RECT 154.230 48.410 154.640 48.830 ;
        RECT 154.840 48.410 155.250 48.830 ;
        RECT 155.450 48.410 155.960 48.830 ;
        RECT 162.000 48.410 162.515 48.830 ;
        RECT 162.705 48.410 163.125 48.830 ;
        RECT 163.315 48.410 163.735 48.830 ;
        RECT 163.925 48.410 164.345 48.830 ;
        RECT 165.410 48.410 165.830 48.830 ;
        RECT 166.020 48.410 166.440 48.830 ;
        RECT 166.630 48.410 167.050 48.830 ;
        RECT 167.240 48.410 167.660 48.830 ;
        RECT 167.850 48.410 168.270 48.830 ;
        RECT 169.325 48.410 169.745 48.830 ;
        RECT 169.935 48.410 170.355 48.830 ;
        RECT 170.545 48.410 170.965 48.830 ;
        RECT 171.155 48.410 171.670 48.830 ;
        RECT 5.415 38.735 6.035 39.455 ;
        RECT 10.900 38.800 11.930 39.390 ;
        RECT 12.120 38.800 12.570 39.390 ;
        RECT 29.060 38.620 30.070 39.560 ;
        RECT 34.915 38.735 35.535 39.455 ;
        RECT 40.400 38.800 41.430 39.390 ;
        RECT 41.620 38.800 42.070 39.390 ;
        RECT 58.560 38.620 59.570 39.560 ;
        RECT 64.415 38.735 65.035 39.455 ;
        RECT 69.900 38.800 70.930 39.390 ;
        RECT 71.120 38.800 71.570 39.390 ;
        RECT 88.060 38.620 89.070 39.560 ;
        RECT 93.915 38.735 94.535 39.455 ;
        RECT 99.400 38.800 100.430 39.390 ;
        RECT 100.620 38.800 101.070 39.390 ;
        RECT 117.560 38.620 118.570 39.560 ;
        RECT 123.415 38.735 124.035 39.455 ;
        RECT 128.900 38.800 129.930 39.390 ;
        RECT 130.120 38.800 130.570 39.390 ;
        RECT 147.060 38.620 148.070 39.560 ;
        RECT 152.915 38.735 153.535 39.455 ;
        RECT 158.400 38.800 159.430 39.390 ;
        RECT 159.620 38.800 160.070 39.390 ;
        RECT 176.560 38.620 177.570 39.560 ;
        RECT 7.355 32.090 7.775 32.510 ;
        RECT 7.965 32.090 8.385 32.510 ;
        RECT 8.575 32.090 8.995 32.510 ;
        RECT 9.185 32.090 9.700 32.510 ;
        RECT 10.500 32.090 11.015 32.510 ;
        RECT 11.205 32.090 11.625 32.510 ;
        RECT 11.815 32.090 12.235 32.510 ;
        RECT 12.425 32.090 12.845 32.510 ;
        RECT 21.150 32.090 21.665 32.510 ;
        RECT 21.855 32.090 22.275 32.510 ;
        RECT 22.465 32.090 22.885 32.510 ;
        RECT 23.075 32.090 23.495 32.510 ;
        RECT 24.550 32.090 24.970 32.510 ;
        RECT 25.160 32.090 25.580 32.510 ;
        RECT 25.770 32.090 26.190 32.510 ;
        RECT 26.380 32.090 26.800 32.510 ;
        RECT 26.990 32.090 27.410 32.510 ;
        RECT 28.475 32.090 28.895 32.510 ;
        RECT 29.085 32.090 29.505 32.510 ;
        RECT 29.695 32.090 30.115 32.510 ;
        RECT 30.305 32.090 30.820 32.510 ;
        RECT 36.855 32.090 37.275 32.510 ;
        RECT 37.465 32.090 37.885 32.510 ;
        RECT 38.075 32.090 38.495 32.510 ;
        RECT 38.685 32.090 39.200 32.510 ;
        RECT 40.000 32.090 40.515 32.510 ;
        RECT 40.705 32.090 41.125 32.510 ;
        RECT 41.315 32.090 41.735 32.510 ;
        RECT 41.925 32.090 42.345 32.510 ;
        RECT 50.650 32.090 51.165 32.510 ;
        RECT 51.355 32.090 51.775 32.510 ;
        RECT 51.965 32.090 52.385 32.510 ;
        RECT 52.575 32.090 52.995 32.510 ;
        RECT 54.050 32.090 54.470 32.510 ;
        RECT 54.660 32.090 55.080 32.510 ;
        RECT 55.270 32.090 55.690 32.510 ;
        RECT 55.880 32.090 56.300 32.510 ;
        RECT 56.490 32.090 56.910 32.510 ;
        RECT 57.975 32.090 58.395 32.510 ;
        RECT 58.585 32.090 59.005 32.510 ;
        RECT 59.195 32.090 59.615 32.510 ;
        RECT 59.805 32.090 60.320 32.510 ;
        RECT 66.355 32.090 66.775 32.510 ;
        RECT 66.965 32.090 67.385 32.510 ;
        RECT 67.575 32.090 67.995 32.510 ;
        RECT 68.185 32.090 68.700 32.510 ;
        RECT 69.500 32.090 70.015 32.510 ;
        RECT 70.205 32.090 70.625 32.510 ;
        RECT 70.815 32.090 71.235 32.510 ;
        RECT 71.425 32.090 71.845 32.510 ;
        RECT 80.150 32.090 80.665 32.510 ;
        RECT 80.855 32.090 81.275 32.510 ;
        RECT 81.465 32.090 81.885 32.510 ;
        RECT 82.075 32.090 82.495 32.510 ;
        RECT 83.550 32.090 83.970 32.510 ;
        RECT 84.160 32.090 84.580 32.510 ;
        RECT 84.770 32.090 85.190 32.510 ;
        RECT 85.380 32.090 85.800 32.510 ;
        RECT 85.990 32.090 86.410 32.510 ;
        RECT 87.475 32.090 87.895 32.510 ;
        RECT 88.085 32.090 88.505 32.510 ;
        RECT 88.695 32.090 89.115 32.510 ;
        RECT 89.305 32.090 89.820 32.510 ;
        RECT 95.855 32.090 96.275 32.510 ;
        RECT 96.465 32.090 96.885 32.510 ;
        RECT 97.075 32.090 97.495 32.510 ;
        RECT 97.685 32.090 98.200 32.510 ;
        RECT 99.000 32.090 99.515 32.510 ;
        RECT 99.705 32.090 100.125 32.510 ;
        RECT 100.315 32.090 100.735 32.510 ;
        RECT 100.925 32.090 101.345 32.510 ;
        RECT 109.650 32.090 110.165 32.510 ;
        RECT 110.355 32.090 110.775 32.510 ;
        RECT 110.965 32.090 111.385 32.510 ;
        RECT 111.575 32.090 111.995 32.510 ;
        RECT 113.050 32.090 113.470 32.510 ;
        RECT 113.660 32.090 114.080 32.510 ;
        RECT 114.270 32.090 114.690 32.510 ;
        RECT 114.880 32.090 115.300 32.510 ;
        RECT 115.490 32.090 115.910 32.510 ;
        RECT 116.975 32.090 117.395 32.510 ;
        RECT 117.585 32.090 118.005 32.510 ;
        RECT 118.195 32.090 118.615 32.510 ;
        RECT 118.805 32.090 119.320 32.510 ;
        RECT 125.355 32.090 125.775 32.510 ;
        RECT 125.965 32.090 126.385 32.510 ;
        RECT 126.575 32.090 126.995 32.510 ;
        RECT 127.185 32.090 127.700 32.510 ;
        RECT 128.500 32.090 129.015 32.510 ;
        RECT 129.205 32.090 129.625 32.510 ;
        RECT 129.815 32.090 130.235 32.510 ;
        RECT 130.425 32.090 130.845 32.510 ;
        RECT 139.150 32.090 139.665 32.510 ;
        RECT 139.855 32.090 140.275 32.510 ;
        RECT 140.465 32.090 140.885 32.510 ;
        RECT 141.075 32.090 141.495 32.510 ;
        RECT 142.550 32.090 142.970 32.510 ;
        RECT 143.160 32.090 143.580 32.510 ;
        RECT 143.770 32.090 144.190 32.510 ;
        RECT 144.380 32.090 144.800 32.510 ;
        RECT 144.990 32.090 145.410 32.510 ;
        RECT 146.475 32.090 146.895 32.510 ;
        RECT 147.085 32.090 147.505 32.510 ;
        RECT 147.695 32.090 148.115 32.510 ;
        RECT 148.305 32.090 148.820 32.510 ;
        RECT 154.855 32.090 155.275 32.510 ;
        RECT 155.465 32.090 155.885 32.510 ;
        RECT 156.075 32.090 156.495 32.510 ;
        RECT 156.685 32.090 157.200 32.510 ;
        RECT 158.000 32.090 158.515 32.510 ;
        RECT 158.705 32.090 159.125 32.510 ;
        RECT 159.315 32.090 159.735 32.510 ;
        RECT 159.925 32.090 160.345 32.510 ;
        RECT 168.650 32.090 169.165 32.510 ;
        RECT 169.355 32.090 169.775 32.510 ;
        RECT 169.965 32.090 170.385 32.510 ;
        RECT 170.575 32.090 170.995 32.510 ;
        RECT 172.050 32.090 172.470 32.510 ;
        RECT 172.660 32.090 173.080 32.510 ;
        RECT 173.270 32.090 173.690 32.510 ;
        RECT 173.880 32.090 174.300 32.510 ;
        RECT 174.490 32.090 174.910 32.510 ;
        RECT 175.975 32.090 176.395 32.510 ;
        RECT 176.585 32.090 177.005 32.510 ;
        RECT 177.195 32.090 177.615 32.510 ;
        RECT 177.805 32.090 178.320 32.510 ;
      LAYER met1 ;
        RECT 16.280 70.140 173.490 70.620 ;
        RECT 19.290 63.915 20.420 64.140 ;
        RECT 43.295 63.915 44.035 63.975 ;
        RECT 48.790 63.915 49.920 64.140 ;
        RECT 72.795 63.915 73.535 63.975 ;
        RECT 78.290 63.915 79.420 64.140 ;
        RECT 102.295 63.915 103.035 63.975 ;
        RECT 107.790 63.915 108.920 64.140 ;
        RECT 131.795 63.915 132.535 63.975 ;
        RECT 137.290 63.915 138.420 64.140 ;
        RECT 161.295 63.915 162.035 63.975 ;
        RECT 17.840 63.255 20.420 63.915 ;
        RECT 35.060 63.910 49.920 63.915 ;
        RECT 64.560 63.910 79.420 63.915 ;
        RECT 94.060 63.910 108.920 63.915 ;
        RECT 123.560 63.910 138.420 63.915 ;
        RECT 153.060 63.910 165.440 63.915 ;
        RECT 19.290 63.040 20.420 63.255 ;
        RECT 25.290 63.255 49.920 63.910 ;
        RECT 25.290 63.250 38.550 63.255 ;
        RECT 43.295 63.195 44.035 63.255 ;
        RECT 48.790 63.040 49.920 63.255 ;
        RECT 54.790 63.255 79.420 63.910 ;
        RECT 54.790 63.250 68.050 63.255 ;
        RECT 72.795 63.195 73.535 63.255 ;
        RECT 78.290 63.040 79.420 63.255 ;
        RECT 84.290 63.255 108.920 63.910 ;
        RECT 84.290 63.250 97.550 63.255 ;
        RECT 102.295 63.195 103.035 63.255 ;
        RECT 107.790 63.040 108.920 63.255 ;
        RECT 113.790 63.255 138.420 63.910 ;
        RECT 113.790 63.250 127.050 63.255 ;
        RECT 131.795 63.195 132.535 63.255 ;
        RECT 137.290 63.040 138.420 63.255 ;
        RECT 143.290 63.255 165.440 63.910 ;
        RECT 143.290 63.250 156.550 63.255 ;
        RECT 161.295 63.195 162.035 63.255 ;
        RECT 17.890 54.290 165.390 54.300 ;
        RECT 17.000 53.810 177.530 54.290 ;
        RECT 175.570 53.460 177.530 53.810 ;
        RECT 2.000 48.380 180.440 48.860 ;
        RECT 5.355 39.425 6.095 39.485 ;
        RECT 10.840 39.425 24.100 39.430 ;
        RECT 2.000 38.770 24.100 39.425 ;
        RECT 28.970 39.425 30.100 39.640 ;
        RECT 34.855 39.425 35.595 39.485 ;
        RECT 40.340 39.425 53.600 39.430 ;
        RECT 28.970 38.770 53.600 39.425 ;
        RECT 58.470 39.425 59.600 39.640 ;
        RECT 64.355 39.425 65.095 39.485 ;
        RECT 69.840 39.425 83.100 39.430 ;
        RECT 58.470 38.770 83.100 39.425 ;
        RECT 87.970 39.425 89.100 39.640 ;
        RECT 93.855 39.425 94.595 39.485 ;
        RECT 99.340 39.425 112.600 39.430 ;
        RECT 87.970 38.770 112.600 39.425 ;
        RECT 117.470 39.425 118.600 39.640 ;
        RECT 123.355 39.425 124.095 39.485 ;
        RECT 128.840 39.425 142.100 39.430 ;
        RECT 117.470 38.770 142.100 39.425 ;
        RECT 146.970 39.425 148.100 39.640 ;
        RECT 152.855 39.425 153.595 39.485 ;
        RECT 158.340 39.425 171.600 39.430 ;
        RECT 146.970 38.770 171.600 39.425 ;
        RECT 176.470 39.425 177.600 39.640 ;
        RECT 176.470 39.395 179.000 39.425 ;
        RECT 172.640 38.795 179.000 39.395 ;
        RECT 2.000 38.765 14.330 38.770 ;
        RECT 28.970 38.765 43.830 38.770 ;
        RECT 58.470 38.765 73.330 38.770 ;
        RECT 87.970 38.765 102.830 38.770 ;
        RECT 117.470 38.765 132.330 38.770 ;
        RECT 146.970 38.765 161.830 38.770 ;
        RECT 176.470 38.765 179.000 38.795 ;
        RECT 5.355 38.705 6.095 38.765 ;
        RECT 28.970 38.540 30.100 38.765 ;
        RECT 34.855 38.705 35.595 38.765 ;
        RECT 58.470 38.540 59.600 38.765 ;
        RECT 64.355 38.705 65.095 38.765 ;
        RECT 87.970 38.540 89.100 38.765 ;
        RECT 93.855 38.705 94.595 38.765 ;
        RECT 117.470 38.540 118.600 38.765 ;
        RECT 123.355 38.705 124.095 38.765 ;
        RECT 146.970 38.540 148.100 38.765 ;
        RECT 152.855 38.705 153.595 38.765 ;
        RECT 176.470 38.540 177.600 38.765 ;
        RECT 2.000 32.060 180.440 32.540 ;
      LAYER via ;
        RECT 39.000 70.240 39.260 70.500 ;
        RECT 39.370 70.240 39.630 70.500 ;
        RECT 39.740 70.240 40.000 70.500 ;
        RECT 70.000 70.240 70.260 70.500 ;
        RECT 70.370 70.240 70.630 70.500 ;
        RECT 70.740 70.240 71.000 70.500 ;
        RECT 112.000 70.240 112.260 70.500 ;
        RECT 112.370 70.240 112.630 70.500 ;
        RECT 112.740 70.240 113.000 70.500 ;
        RECT 143.000 70.240 143.260 70.500 ;
        RECT 143.370 70.240 143.630 70.500 ;
        RECT 143.740 70.240 144.000 70.500 ;
        RECT 172.490 70.250 172.750 70.510 ;
        RECT 172.810 70.250 173.070 70.510 ;
        RECT 173.130 70.250 173.390 70.510 ;
        RECT 18.045 63.295 18.625 63.875 ;
        RECT 164.480 63.295 165.380 63.875 ;
        RECT 39.000 53.920 39.260 54.180 ;
        RECT 39.370 53.920 39.630 54.180 ;
        RECT 39.740 53.920 40.000 54.180 ;
        RECT 70.000 53.920 70.260 54.180 ;
        RECT 70.370 53.920 70.630 54.180 ;
        RECT 70.740 53.920 71.000 54.180 ;
        RECT 112.000 53.920 112.260 54.180 ;
        RECT 112.370 53.920 112.630 54.180 ;
        RECT 112.740 53.920 113.000 54.180 ;
        RECT 143.000 53.920 143.260 54.180 ;
        RECT 143.370 53.920 143.630 54.180 ;
        RECT 143.740 53.920 144.000 54.180 ;
        RECT 172.470 53.950 172.730 54.210 ;
        RECT 172.830 53.950 173.090 54.210 ;
        RECT 173.190 53.950 173.450 54.210 ;
        RECT 173.550 53.950 173.810 54.210 ;
        RECT 173.920 53.950 174.180 54.210 ;
        RECT 174.280 53.950 174.540 54.210 ;
        RECT 174.660 53.950 174.920 54.210 ;
        RECT 175.035 53.950 175.295 54.210 ;
        RECT 175.415 53.950 175.675 54.210 ;
        RECT 175.790 53.950 176.050 54.210 ;
        RECT 176.165 53.950 176.425 54.210 ;
        RECT 176.535 53.950 176.795 54.210 ;
        RECT 176.915 53.950 177.175 54.210 ;
        RECT 39.000 48.480 39.260 48.740 ;
        RECT 39.370 48.480 39.630 48.740 ;
        RECT 39.740 48.480 40.000 48.740 ;
        RECT 70.000 48.480 70.260 48.740 ;
        RECT 70.370 48.480 70.630 48.740 ;
        RECT 70.740 48.480 71.000 48.740 ;
        RECT 112.000 48.480 112.260 48.740 ;
        RECT 112.370 48.480 112.630 48.740 ;
        RECT 112.740 48.480 113.000 48.740 ;
        RECT 143.000 48.480 143.260 48.740 ;
        RECT 143.370 48.480 143.630 48.740 ;
        RECT 143.740 48.480 144.000 48.740 ;
        RECT 179.465 48.490 179.725 48.750 ;
        RECT 179.785 48.490 180.045 48.750 ;
        RECT 180.105 48.490 180.365 48.750 ;
        RECT 4.055 38.805 4.635 39.385 ;
        RECT 172.760 38.805 173.340 39.385 ;
        RECT 39.000 32.160 39.260 32.420 ;
        RECT 39.370 32.160 39.630 32.420 ;
        RECT 39.740 32.160 40.000 32.420 ;
        RECT 70.000 32.160 70.260 32.420 ;
        RECT 70.370 32.160 70.630 32.420 ;
        RECT 70.740 32.160 71.000 32.420 ;
        RECT 112.000 32.160 112.260 32.420 ;
        RECT 112.370 32.160 112.630 32.420 ;
        RECT 112.740 32.160 113.000 32.420 ;
        RECT 143.000 32.160 143.260 32.420 ;
        RECT 143.370 32.160 143.630 32.420 ;
        RECT 143.740 32.160 144.000 32.420 ;
        RECT 179.475 32.170 179.735 32.430 ;
        RECT 179.795 32.170 180.055 32.430 ;
        RECT 180.115 32.170 180.375 32.430 ;
      LAYER met2 ;
        RECT 39.000 70.170 40.000 70.570 ;
        RECT 70.000 70.170 71.000 70.570 ;
        RECT 112.000 70.170 113.000 70.570 ;
        RECT 143.000 70.170 144.000 70.570 ;
        RECT 17.890 63.935 18.785 63.965 ;
        RECT 14.420 63.235 18.785 63.935 ;
        RECT 14.420 52.350 15.120 63.235 ;
        RECT 17.890 63.205 18.785 63.235 ;
        RECT 164.470 63.935 165.390 63.965 ;
        RECT 164.470 63.235 169.490 63.935 ;
        RECT 164.470 63.205 165.390 63.235 ;
        RECT 39.000 53.850 40.000 54.250 ;
        RECT 70.000 53.850 71.000 54.250 ;
        RECT 112.000 53.850 113.000 54.250 ;
        RECT 143.000 53.850 144.000 54.250 ;
        RECT 4.000 51.650 15.120 52.350 ;
        RECT 4.000 50.835 4.700 51.650 ;
        RECT 3.995 45.265 4.700 50.835 ;
        RECT 168.790 49.935 169.490 63.235 ;
        RECT 172.440 54.540 173.440 70.670 ;
        RECT 172.440 53.540 180.440 54.540 ;
        RECT 179.440 53.000 180.435 53.540 ;
        RECT 168.790 49.235 173.400 49.935 ;
        RECT 39.000 48.410 40.000 48.810 ;
        RECT 70.000 48.410 71.000 48.810 ;
        RECT 112.000 48.410 113.000 48.810 ;
        RECT 143.000 48.410 144.000 48.810 ;
        RECT 3.995 38.715 4.695 45.265 ;
        RECT 172.700 38.745 173.400 49.235 ;
        RECT 39.000 32.090 40.000 32.490 ;
        RECT 70.000 32.090 71.000 32.490 ;
        RECT 112.000 32.090 113.000 32.490 ;
        RECT 143.000 32.090 144.000 32.490 ;
        RECT 179.440 32.010 180.440 53.000 ;
      LAYER via2 ;
        RECT 39.100 70.220 39.400 70.520 ;
        RECT 39.600 70.220 39.900 70.520 ;
        RECT 70.100 70.220 70.400 70.520 ;
        RECT 70.600 70.220 70.900 70.520 ;
        RECT 112.100 70.220 112.400 70.520 ;
        RECT 112.600 70.220 112.900 70.520 ;
        RECT 143.100 70.220 143.400 70.520 ;
        RECT 143.600 70.220 143.900 70.520 ;
        RECT 39.100 53.900 39.400 54.200 ;
        RECT 39.600 53.900 39.900 54.200 ;
        RECT 70.100 53.900 70.400 54.200 ;
        RECT 70.600 53.900 70.900 54.200 ;
        RECT 112.100 53.900 112.400 54.200 ;
        RECT 112.600 53.900 112.900 54.200 ;
        RECT 143.100 53.900 143.400 54.200 ;
        RECT 143.600 53.900 143.900 54.200 ;
        RECT 179.750 51.400 180.150 51.800 ;
        RECT 179.750 50.870 180.150 51.270 ;
        RECT 39.100 48.460 39.400 48.760 ;
        RECT 39.600 48.460 39.900 48.760 ;
        RECT 70.100 48.460 70.400 48.760 ;
        RECT 70.600 48.460 70.900 48.760 ;
        RECT 112.100 48.460 112.400 48.760 ;
        RECT 112.600 48.460 112.900 48.760 ;
        RECT 143.100 48.460 143.400 48.760 ;
        RECT 143.600 48.460 143.900 48.760 ;
        RECT 39.100 32.140 39.400 32.440 ;
        RECT 39.600 32.140 39.900 32.440 ;
        RECT 70.100 32.140 70.400 32.440 ;
        RECT 70.600 32.140 70.900 32.440 ;
        RECT 112.100 32.140 112.400 32.440 ;
        RECT 112.600 32.140 112.900 32.440 ;
        RECT 143.100 32.140 143.400 32.440 ;
        RECT 143.600 32.140 143.900 32.440 ;
      LAYER met3 ;
        RECT 39.000 51.910 40.000 70.620 ;
        RECT 70.000 51.910 71.000 70.620 ;
        RECT 112.000 51.910 113.000 70.620 ;
        RECT 143.000 51.910 144.000 70.620 ;
        RECT 39.000 50.760 180.440 51.910 ;
        RECT 39.000 32.060 40.000 50.760 ;
        RECT 70.000 32.060 71.000 50.760 ;
        RECT 112.000 32.060 113.000 50.760 ;
        RECT 143.000 32.060 144.000 50.760 ;
  END
END vco_r100
END LIBRARY

