magic
tech sky130A
magscale 1 2
timestamp 1624033926
<< obsli1 >>
rect 1104 1445 178848 117521
<< obsm1 >>
rect 382 1368 179570 117768
<< metal2 >>
rect 386 119200 442 120000
rect 1214 119200 1270 120000
rect 2134 119200 2190 120000
rect 2962 119200 3018 120000
rect 3882 119200 3938 120000
rect 4802 119200 4858 120000
rect 5630 119200 5686 120000
rect 6550 119200 6606 120000
rect 7470 119200 7526 120000
rect 8298 119200 8354 120000
rect 9218 119200 9274 120000
rect 10138 119200 10194 120000
rect 10966 119200 11022 120000
rect 11886 119200 11942 120000
rect 12714 119200 12770 120000
rect 13634 119200 13690 120000
rect 14554 119200 14610 120000
rect 15382 119200 15438 120000
rect 16302 119200 16358 120000
rect 17222 119200 17278 120000
rect 18050 119200 18106 120000
rect 18970 119200 19026 120000
rect 19890 119200 19946 120000
rect 20718 119200 20774 120000
rect 21638 119200 21694 120000
rect 22558 119200 22614 120000
rect 23386 119200 23442 120000
rect 24306 119200 24362 120000
rect 25134 119200 25190 120000
rect 26054 119200 26110 120000
rect 26974 119200 27030 120000
rect 27802 119200 27858 120000
rect 28722 119200 28778 120000
rect 29642 119200 29698 120000
rect 30470 119200 30526 120000
rect 31390 119200 31446 120000
rect 32310 119200 32366 120000
rect 33138 119200 33194 120000
rect 34058 119200 34114 120000
rect 34886 119200 34942 120000
rect 35806 119200 35862 120000
rect 36726 119200 36782 120000
rect 37554 119200 37610 120000
rect 38474 119200 38530 120000
rect 39394 119200 39450 120000
rect 40222 119200 40278 120000
rect 41142 119200 41198 120000
rect 42062 119200 42118 120000
rect 42890 119200 42946 120000
rect 43810 119200 43866 120000
rect 44730 119200 44786 120000
rect 45558 119200 45614 120000
rect 46478 119200 46534 120000
rect 47306 119200 47362 120000
rect 48226 119200 48282 120000
rect 49146 119200 49202 120000
rect 49974 119200 50030 120000
rect 50894 119200 50950 120000
rect 51814 119200 51870 120000
rect 52642 119200 52698 120000
rect 53562 119200 53618 120000
rect 54482 119200 54538 120000
rect 55310 119200 55366 120000
rect 56230 119200 56286 120000
rect 57058 119200 57114 120000
rect 57978 119200 58034 120000
rect 58898 119200 58954 120000
rect 59726 119200 59782 120000
rect 60646 119200 60702 120000
rect 61566 119200 61622 120000
rect 62394 119200 62450 120000
rect 63314 119200 63370 120000
rect 64234 119200 64290 120000
rect 65062 119200 65118 120000
rect 65982 119200 66038 120000
rect 66902 119200 66958 120000
rect 67730 119200 67786 120000
rect 68650 119200 68706 120000
rect 69478 119200 69534 120000
rect 70398 119200 70454 120000
rect 71318 119200 71374 120000
rect 72146 119200 72202 120000
rect 73066 119200 73122 120000
rect 73986 119200 74042 120000
rect 74814 119200 74870 120000
rect 75734 119200 75790 120000
rect 76654 119200 76710 120000
rect 77482 119200 77538 120000
rect 78402 119200 78458 120000
rect 79230 119200 79286 120000
rect 80150 119200 80206 120000
rect 81070 119200 81126 120000
rect 81898 119200 81954 120000
rect 82818 119200 82874 120000
rect 83738 119200 83794 120000
rect 84566 119200 84622 120000
rect 85486 119200 85542 120000
rect 86406 119200 86462 120000
rect 87234 119200 87290 120000
rect 88154 119200 88210 120000
rect 89074 119200 89130 120000
rect 89902 119200 89958 120000
rect 90822 119200 90878 120000
rect 91650 119200 91706 120000
rect 92570 119200 92626 120000
rect 93490 119200 93546 120000
rect 94318 119200 94374 120000
rect 95238 119200 95294 120000
rect 96158 119200 96214 120000
rect 96986 119200 97042 120000
rect 97906 119200 97962 120000
rect 98826 119200 98882 120000
rect 99654 119200 99710 120000
rect 100574 119200 100630 120000
rect 101494 119200 101550 120000
rect 102322 119200 102378 120000
rect 103242 119200 103298 120000
rect 104070 119200 104126 120000
rect 104990 119200 105046 120000
rect 105910 119200 105966 120000
rect 106738 119200 106794 120000
rect 107658 119200 107714 120000
rect 108578 119200 108634 120000
rect 109406 119200 109462 120000
rect 110326 119200 110382 120000
rect 111246 119200 111302 120000
rect 112074 119200 112130 120000
rect 112994 119200 113050 120000
rect 113822 119200 113878 120000
rect 114742 119200 114798 120000
rect 115662 119200 115718 120000
rect 116490 119200 116546 120000
rect 117410 119200 117466 120000
rect 118330 119200 118386 120000
rect 119158 119200 119214 120000
rect 120078 119200 120134 120000
rect 120998 119200 121054 120000
rect 121826 119200 121882 120000
rect 122746 119200 122802 120000
rect 123666 119200 123722 120000
rect 124494 119200 124550 120000
rect 125414 119200 125470 120000
rect 126242 119200 126298 120000
rect 127162 119200 127218 120000
rect 128082 119200 128138 120000
rect 128910 119200 128966 120000
rect 129830 119200 129886 120000
rect 130750 119200 130806 120000
rect 131578 119200 131634 120000
rect 132498 119200 132554 120000
rect 133418 119200 133474 120000
rect 134246 119200 134302 120000
rect 135166 119200 135222 120000
rect 135994 119200 136050 120000
rect 136914 119200 136970 120000
rect 137834 119200 137890 120000
rect 138662 119200 138718 120000
rect 139582 119200 139638 120000
rect 140502 119200 140558 120000
rect 141330 119200 141386 120000
rect 142250 119200 142306 120000
rect 143170 119200 143226 120000
rect 143998 119200 144054 120000
rect 144918 119200 144974 120000
rect 145838 119200 145894 120000
rect 146666 119200 146722 120000
rect 147586 119200 147642 120000
rect 148414 119200 148470 120000
rect 149334 119200 149390 120000
rect 150254 119200 150310 120000
rect 151082 119200 151138 120000
rect 152002 119200 152058 120000
rect 152922 119200 152978 120000
rect 153750 119200 153806 120000
rect 154670 119200 154726 120000
rect 155590 119200 155646 120000
rect 156418 119200 156474 120000
rect 157338 119200 157394 120000
rect 158166 119200 158222 120000
rect 159086 119200 159142 120000
rect 160006 119200 160062 120000
rect 160834 119200 160890 120000
rect 161754 119200 161810 120000
rect 162674 119200 162730 120000
rect 163502 119200 163558 120000
rect 164422 119200 164478 120000
rect 165342 119200 165398 120000
rect 166170 119200 166226 120000
rect 167090 119200 167146 120000
rect 168010 119200 168066 120000
rect 168838 119200 168894 120000
rect 169758 119200 169814 120000
rect 170586 119200 170642 120000
rect 171506 119200 171562 120000
rect 172426 119200 172482 120000
rect 173254 119200 173310 120000
rect 174174 119200 174230 120000
rect 175094 119200 175150 120000
rect 175922 119200 175978 120000
rect 176842 119200 176898 120000
rect 177762 119200 177818 120000
rect 178590 119200 178646 120000
rect 179510 119200 179566 120000
rect 570 0 626 800
rect 1766 0 1822 800
rect 3054 0 3110 800
rect 4342 0 4398 800
rect 5630 0 5686 800
rect 6918 0 6974 800
rect 8206 0 8262 800
rect 9494 0 9550 800
rect 10782 0 10838 800
rect 12070 0 12126 800
rect 13358 0 13414 800
rect 14646 0 14702 800
rect 15934 0 15990 800
rect 17222 0 17278 800
rect 18510 0 18566 800
rect 19798 0 19854 800
rect 21086 0 21142 800
rect 22374 0 22430 800
rect 23662 0 23718 800
rect 24950 0 25006 800
rect 26238 0 26294 800
rect 27526 0 27582 800
rect 28814 0 28870 800
rect 30102 0 30158 800
rect 31390 0 31446 800
rect 32678 0 32734 800
rect 33966 0 34022 800
rect 35254 0 35310 800
rect 36542 0 36598 800
rect 37830 0 37886 800
rect 39118 0 39174 800
rect 40406 0 40462 800
rect 41694 0 41750 800
rect 42982 0 43038 800
rect 44270 0 44326 800
rect 45558 0 45614 800
rect 46846 0 46902 800
rect 48134 0 48190 800
rect 49422 0 49478 800
rect 50710 0 50766 800
rect 51998 0 52054 800
rect 53286 0 53342 800
rect 54574 0 54630 800
rect 55862 0 55918 800
rect 57150 0 57206 800
rect 58438 0 58494 800
rect 59726 0 59782 800
rect 60922 0 60978 800
rect 62210 0 62266 800
rect 63498 0 63554 800
rect 64786 0 64842 800
rect 66074 0 66130 800
rect 67362 0 67418 800
rect 68650 0 68706 800
rect 69938 0 69994 800
rect 71226 0 71282 800
rect 72514 0 72570 800
rect 73802 0 73858 800
rect 75090 0 75146 800
rect 76378 0 76434 800
rect 77666 0 77722 800
rect 78954 0 79010 800
rect 80242 0 80298 800
rect 81530 0 81586 800
rect 82818 0 82874 800
rect 84106 0 84162 800
rect 85394 0 85450 800
rect 86682 0 86738 800
rect 87970 0 88026 800
rect 89258 0 89314 800
rect 90546 0 90602 800
rect 91834 0 91890 800
rect 93122 0 93178 800
rect 94410 0 94466 800
rect 95698 0 95754 800
rect 96986 0 97042 800
rect 98274 0 98330 800
rect 99562 0 99618 800
rect 100850 0 100906 800
rect 102138 0 102194 800
rect 103426 0 103482 800
rect 104714 0 104770 800
rect 106002 0 106058 800
rect 107290 0 107346 800
rect 108578 0 108634 800
rect 109866 0 109922 800
rect 111154 0 111210 800
rect 112442 0 112498 800
rect 113730 0 113786 800
rect 115018 0 115074 800
rect 116306 0 116362 800
rect 117594 0 117650 800
rect 118882 0 118938 800
rect 120170 0 120226 800
rect 121366 0 121422 800
rect 122654 0 122710 800
rect 123942 0 123998 800
rect 125230 0 125286 800
rect 126518 0 126574 800
rect 127806 0 127862 800
rect 129094 0 129150 800
rect 130382 0 130438 800
rect 131670 0 131726 800
rect 132958 0 133014 800
rect 134246 0 134302 800
rect 135534 0 135590 800
rect 136822 0 136878 800
rect 138110 0 138166 800
rect 139398 0 139454 800
rect 140686 0 140742 800
rect 141974 0 142030 800
rect 143262 0 143318 800
rect 144550 0 144606 800
rect 145838 0 145894 800
rect 147126 0 147182 800
rect 148414 0 148470 800
rect 149702 0 149758 800
rect 150990 0 151046 800
rect 152278 0 152334 800
rect 153566 0 153622 800
rect 154854 0 154910 800
rect 156142 0 156198 800
rect 157430 0 157486 800
rect 158718 0 158774 800
rect 160006 0 160062 800
rect 161294 0 161350 800
rect 162582 0 162638 800
rect 163870 0 163926 800
rect 165158 0 165214 800
rect 166446 0 166502 800
rect 167734 0 167790 800
rect 169022 0 169078 800
rect 170310 0 170366 800
rect 171598 0 171654 800
rect 172886 0 172942 800
rect 174174 0 174230 800
rect 175462 0 175518 800
rect 176750 0 176806 800
rect 178038 0 178094 800
rect 179326 0 179382 800
<< obsm2 >>
rect 498 119144 1158 119785
rect 1326 119144 2078 119785
rect 2246 119144 2906 119785
rect 3074 119144 3826 119785
rect 3994 119144 4746 119785
rect 4914 119144 5574 119785
rect 5742 119144 6494 119785
rect 6662 119144 7414 119785
rect 7582 119144 8242 119785
rect 8410 119144 9162 119785
rect 9330 119144 10082 119785
rect 10250 119144 10910 119785
rect 11078 119144 11830 119785
rect 11998 119144 12658 119785
rect 12826 119144 13578 119785
rect 13746 119144 14498 119785
rect 14666 119144 15326 119785
rect 15494 119144 16246 119785
rect 16414 119144 17166 119785
rect 17334 119144 17994 119785
rect 18162 119144 18914 119785
rect 19082 119144 19834 119785
rect 20002 119144 20662 119785
rect 20830 119144 21582 119785
rect 21750 119144 22502 119785
rect 22670 119144 23330 119785
rect 23498 119144 24250 119785
rect 24418 119144 25078 119785
rect 25246 119144 25998 119785
rect 26166 119144 26918 119785
rect 27086 119144 27746 119785
rect 27914 119144 28666 119785
rect 28834 119144 29586 119785
rect 29754 119144 30414 119785
rect 30582 119144 31334 119785
rect 31502 119144 32254 119785
rect 32422 119144 33082 119785
rect 33250 119144 34002 119785
rect 34170 119144 34830 119785
rect 34998 119144 35750 119785
rect 35918 119144 36670 119785
rect 36838 119144 37498 119785
rect 37666 119144 38418 119785
rect 38586 119144 39338 119785
rect 39506 119144 40166 119785
rect 40334 119144 41086 119785
rect 41254 119144 42006 119785
rect 42174 119144 42834 119785
rect 43002 119144 43754 119785
rect 43922 119144 44674 119785
rect 44842 119144 45502 119785
rect 45670 119144 46422 119785
rect 46590 119144 47250 119785
rect 47418 119144 48170 119785
rect 48338 119144 49090 119785
rect 49258 119144 49918 119785
rect 50086 119144 50838 119785
rect 51006 119144 51758 119785
rect 51926 119144 52586 119785
rect 52754 119144 53506 119785
rect 53674 119144 54426 119785
rect 54594 119144 55254 119785
rect 55422 119144 56174 119785
rect 56342 119144 57002 119785
rect 57170 119144 57922 119785
rect 58090 119144 58842 119785
rect 59010 119144 59670 119785
rect 59838 119144 60590 119785
rect 60758 119144 61510 119785
rect 61678 119144 62338 119785
rect 62506 119144 63258 119785
rect 63426 119144 64178 119785
rect 64346 119144 65006 119785
rect 65174 119144 65926 119785
rect 66094 119144 66846 119785
rect 67014 119144 67674 119785
rect 67842 119144 68594 119785
rect 68762 119144 69422 119785
rect 69590 119144 70342 119785
rect 70510 119144 71262 119785
rect 71430 119144 72090 119785
rect 72258 119144 73010 119785
rect 73178 119144 73930 119785
rect 74098 119144 74758 119785
rect 74926 119144 75678 119785
rect 75846 119144 76598 119785
rect 76766 119144 77426 119785
rect 77594 119144 78346 119785
rect 78514 119144 79174 119785
rect 79342 119144 80094 119785
rect 80262 119144 81014 119785
rect 81182 119144 81842 119785
rect 82010 119144 82762 119785
rect 82930 119144 83682 119785
rect 83850 119144 84510 119785
rect 84678 119144 85430 119785
rect 85598 119144 86350 119785
rect 86518 119144 87178 119785
rect 87346 119144 88098 119785
rect 88266 119144 89018 119785
rect 89186 119144 89846 119785
rect 90014 119144 90766 119785
rect 90934 119144 91594 119785
rect 91762 119144 92514 119785
rect 92682 119144 93434 119785
rect 93602 119144 94262 119785
rect 94430 119144 95182 119785
rect 95350 119144 96102 119785
rect 96270 119144 96930 119785
rect 97098 119144 97850 119785
rect 98018 119144 98770 119785
rect 98938 119144 99598 119785
rect 99766 119144 100518 119785
rect 100686 119144 101438 119785
rect 101606 119144 102266 119785
rect 102434 119144 103186 119785
rect 103354 119144 104014 119785
rect 104182 119144 104934 119785
rect 105102 119144 105854 119785
rect 106022 119144 106682 119785
rect 106850 119144 107602 119785
rect 107770 119144 108522 119785
rect 108690 119144 109350 119785
rect 109518 119144 110270 119785
rect 110438 119144 111190 119785
rect 111358 119144 112018 119785
rect 112186 119144 112938 119785
rect 113106 119144 113766 119785
rect 113934 119144 114686 119785
rect 114854 119144 115606 119785
rect 115774 119144 116434 119785
rect 116602 119144 117354 119785
rect 117522 119144 118274 119785
rect 118442 119144 119102 119785
rect 119270 119144 120022 119785
rect 120190 119144 120942 119785
rect 121110 119144 121770 119785
rect 121938 119144 122690 119785
rect 122858 119144 123610 119785
rect 123778 119144 124438 119785
rect 124606 119144 125358 119785
rect 125526 119144 126186 119785
rect 126354 119144 127106 119785
rect 127274 119144 128026 119785
rect 128194 119144 128854 119785
rect 129022 119144 129774 119785
rect 129942 119144 130694 119785
rect 130862 119144 131522 119785
rect 131690 119144 132442 119785
rect 132610 119144 133362 119785
rect 133530 119144 134190 119785
rect 134358 119144 135110 119785
rect 135278 119144 135938 119785
rect 136106 119144 136858 119785
rect 137026 119144 137778 119785
rect 137946 119144 138606 119785
rect 138774 119144 139526 119785
rect 139694 119144 140446 119785
rect 140614 119144 141274 119785
rect 141442 119144 142194 119785
rect 142362 119144 143114 119785
rect 143282 119144 143942 119785
rect 144110 119144 144862 119785
rect 145030 119144 145782 119785
rect 145950 119144 146610 119785
rect 146778 119144 147530 119785
rect 147698 119144 148358 119785
rect 148526 119144 149278 119785
rect 149446 119144 150198 119785
rect 150366 119144 151026 119785
rect 151194 119144 151946 119785
rect 152114 119144 152866 119785
rect 153034 119144 153694 119785
rect 153862 119144 154614 119785
rect 154782 119144 155534 119785
rect 155702 119144 156362 119785
rect 156530 119144 157282 119785
rect 157450 119144 158110 119785
rect 158278 119144 159030 119785
rect 159198 119144 159950 119785
rect 160118 119144 160778 119785
rect 160946 119144 161698 119785
rect 161866 119144 162618 119785
rect 162786 119144 163446 119785
rect 163614 119144 164366 119785
rect 164534 119144 165286 119785
rect 165454 119144 166114 119785
rect 166282 119144 167034 119785
rect 167202 119144 167954 119785
rect 168122 119144 168782 119785
rect 168950 119144 169702 119785
rect 169870 119144 170530 119785
rect 170698 119144 171450 119785
rect 171618 119144 172370 119785
rect 172538 119144 173198 119785
rect 173366 119144 174118 119785
rect 174286 119144 175038 119785
rect 175206 119144 175866 119785
rect 176034 119144 176786 119785
rect 176954 119144 177706 119785
rect 177874 119144 178534 119785
rect 178702 119144 179454 119785
rect 388 856 179564 119144
rect 388 167 514 856
rect 682 167 1710 856
rect 1878 167 2998 856
rect 3166 167 4286 856
rect 4454 167 5574 856
rect 5742 167 6862 856
rect 7030 167 8150 856
rect 8318 167 9438 856
rect 9606 167 10726 856
rect 10894 167 12014 856
rect 12182 167 13302 856
rect 13470 167 14590 856
rect 14758 167 15878 856
rect 16046 167 17166 856
rect 17334 167 18454 856
rect 18622 167 19742 856
rect 19910 167 21030 856
rect 21198 167 22318 856
rect 22486 167 23606 856
rect 23774 167 24894 856
rect 25062 167 26182 856
rect 26350 167 27470 856
rect 27638 167 28758 856
rect 28926 167 30046 856
rect 30214 167 31334 856
rect 31502 167 32622 856
rect 32790 167 33910 856
rect 34078 167 35198 856
rect 35366 167 36486 856
rect 36654 167 37774 856
rect 37942 167 39062 856
rect 39230 167 40350 856
rect 40518 167 41638 856
rect 41806 167 42926 856
rect 43094 167 44214 856
rect 44382 167 45502 856
rect 45670 167 46790 856
rect 46958 167 48078 856
rect 48246 167 49366 856
rect 49534 167 50654 856
rect 50822 167 51942 856
rect 52110 167 53230 856
rect 53398 167 54518 856
rect 54686 167 55806 856
rect 55974 167 57094 856
rect 57262 167 58382 856
rect 58550 167 59670 856
rect 59838 167 60866 856
rect 61034 167 62154 856
rect 62322 167 63442 856
rect 63610 167 64730 856
rect 64898 167 66018 856
rect 66186 167 67306 856
rect 67474 167 68594 856
rect 68762 167 69882 856
rect 70050 167 71170 856
rect 71338 167 72458 856
rect 72626 167 73746 856
rect 73914 167 75034 856
rect 75202 167 76322 856
rect 76490 167 77610 856
rect 77778 167 78898 856
rect 79066 167 80186 856
rect 80354 167 81474 856
rect 81642 167 82762 856
rect 82930 167 84050 856
rect 84218 167 85338 856
rect 85506 167 86626 856
rect 86794 167 87914 856
rect 88082 167 89202 856
rect 89370 167 90490 856
rect 90658 167 91778 856
rect 91946 167 93066 856
rect 93234 167 94354 856
rect 94522 167 95642 856
rect 95810 167 96930 856
rect 97098 167 98218 856
rect 98386 167 99506 856
rect 99674 167 100794 856
rect 100962 167 102082 856
rect 102250 167 103370 856
rect 103538 167 104658 856
rect 104826 167 105946 856
rect 106114 167 107234 856
rect 107402 167 108522 856
rect 108690 167 109810 856
rect 109978 167 111098 856
rect 111266 167 112386 856
rect 112554 167 113674 856
rect 113842 167 114962 856
rect 115130 167 116250 856
rect 116418 167 117538 856
rect 117706 167 118826 856
rect 118994 167 120114 856
rect 120282 167 121310 856
rect 121478 167 122598 856
rect 122766 167 123886 856
rect 124054 167 125174 856
rect 125342 167 126462 856
rect 126630 167 127750 856
rect 127918 167 129038 856
rect 129206 167 130326 856
rect 130494 167 131614 856
rect 131782 167 132902 856
rect 133070 167 134190 856
rect 134358 167 135478 856
rect 135646 167 136766 856
rect 136934 167 138054 856
rect 138222 167 139342 856
rect 139510 167 140630 856
rect 140798 167 141918 856
rect 142086 167 143206 856
rect 143374 167 144494 856
rect 144662 167 145782 856
rect 145950 167 147070 856
rect 147238 167 148358 856
rect 148526 167 149646 856
rect 149814 167 150934 856
rect 151102 167 152222 856
rect 152390 167 153510 856
rect 153678 167 154798 856
rect 154966 167 156086 856
rect 156254 167 157374 856
rect 157542 167 158662 856
rect 158830 167 159950 856
rect 160118 167 161238 856
rect 161406 167 162526 856
rect 162694 167 163814 856
rect 163982 167 165102 856
rect 165270 167 166390 856
rect 166558 167 167678 856
rect 167846 167 168966 856
rect 169134 167 170254 856
rect 170422 167 171542 856
rect 171710 167 172830 856
rect 172998 167 174118 856
rect 174286 167 175406 856
rect 175574 167 176694 856
rect 176862 167 177982 856
rect 178150 167 179270 856
rect 179438 167 179564 856
<< metal3 >>
rect 0 119688 800 119808
rect 0 119416 800 119536
rect 0 119144 800 119264
rect 0 118872 800 118992
rect 0 118600 800 118720
rect 0 118328 800 118448
rect 0 117920 800 118040
rect 179200 117920 180000 118040
rect 0 117648 800 117768
rect 0 117376 800 117496
rect 0 117104 800 117224
rect 0 116832 800 116952
rect 0 116560 800 116680
rect 0 116152 800 116272
rect 0 115880 800 116000
rect 0 115608 800 115728
rect 0 115336 800 115456
rect 0 115064 800 115184
rect 0 114792 800 114912
rect 0 114384 800 114504
rect 0 114112 800 114232
rect 179200 114112 180000 114232
rect 0 113840 800 113960
rect 0 113568 800 113688
rect 0 113296 800 113416
rect 0 113024 800 113144
rect 0 112616 800 112736
rect 0 112344 800 112464
rect 0 112072 800 112192
rect 0 111800 800 111920
rect 0 111528 800 111648
rect 0 111256 800 111376
rect 0 110848 800 110968
rect 0 110576 800 110696
rect 0 110304 800 110424
rect 0 110032 800 110152
rect 179200 110168 180000 110288
rect 0 109760 800 109880
rect 0 109488 800 109608
rect 0 109216 800 109336
rect 0 108808 800 108928
rect 0 108536 800 108656
rect 0 108264 800 108384
rect 0 107992 800 108112
rect 0 107720 800 107840
rect 0 107448 800 107568
rect 0 107040 800 107160
rect 0 106768 800 106888
rect 0 106496 800 106616
rect 0 106224 800 106344
rect 179200 106360 180000 106480
rect 0 105952 800 106072
rect 0 105680 800 105800
rect 0 105272 800 105392
rect 0 105000 800 105120
rect 0 104728 800 104848
rect 0 104456 800 104576
rect 0 104184 800 104304
rect 0 103912 800 104032
rect 0 103504 800 103624
rect 0 103232 800 103352
rect 0 102960 800 103080
rect 0 102688 800 102808
rect 0 102416 800 102536
rect 179200 102416 180000 102536
rect 0 102144 800 102264
rect 0 101736 800 101856
rect 0 101464 800 101584
rect 0 101192 800 101312
rect 0 100920 800 101040
rect 0 100648 800 100768
rect 0 100376 800 100496
rect 0 100104 800 100224
rect 0 99696 800 99816
rect 0 99424 800 99544
rect 0 99152 800 99272
rect 0 98880 800 99000
rect 0 98608 800 98728
rect 179200 98608 180000 98728
rect 0 98336 800 98456
rect 0 97928 800 98048
rect 0 97656 800 97776
rect 0 97384 800 97504
rect 0 97112 800 97232
rect 0 96840 800 96960
rect 0 96568 800 96688
rect 0 96160 800 96280
rect 0 95888 800 96008
rect 0 95616 800 95736
rect 0 95344 800 95464
rect 0 95072 800 95192
rect 0 94800 800 94920
rect 179200 94664 180000 94784
rect 0 94392 800 94512
rect 0 94120 800 94240
rect 0 93848 800 93968
rect 0 93576 800 93696
rect 0 93304 800 93424
rect 0 93032 800 93152
rect 0 92624 800 92744
rect 0 92352 800 92472
rect 0 92080 800 92200
rect 0 91808 800 91928
rect 0 91536 800 91656
rect 0 91264 800 91384
rect 0 90856 800 90976
rect 179200 90856 180000 90976
rect 0 90584 800 90704
rect 0 90312 800 90432
rect 0 90040 800 90160
rect 0 89768 800 89888
rect 0 89496 800 89616
rect 0 89224 800 89344
rect 0 88816 800 88936
rect 0 88544 800 88664
rect 0 88272 800 88392
rect 0 88000 800 88120
rect 0 87728 800 87848
rect 0 87456 800 87576
rect 0 87048 800 87168
rect 0 86776 800 86896
rect 179200 86912 180000 87032
rect 0 86504 800 86624
rect 0 86232 800 86352
rect 0 85960 800 86080
rect 0 85688 800 85808
rect 0 85280 800 85400
rect 0 85008 800 85128
rect 0 84736 800 84856
rect 0 84464 800 84584
rect 0 84192 800 84312
rect 0 83920 800 84040
rect 0 83512 800 83632
rect 0 83240 800 83360
rect 0 82968 800 83088
rect 179200 83104 180000 83224
rect 0 82696 800 82816
rect 0 82424 800 82544
rect 0 82152 800 82272
rect 0 81744 800 81864
rect 0 81472 800 81592
rect 0 81200 800 81320
rect 0 80928 800 81048
rect 0 80656 800 80776
rect 0 80384 800 80504
rect 0 80112 800 80232
rect 0 79704 800 79824
rect 0 79432 800 79552
rect 0 79160 800 79280
rect 179200 79296 180000 79416
rect 0 78888 800 79008
rect 0 78616 800 78736
rect 0 78344 800 78464
rect 0 77936 800 78056
rect 0 77664 800 77784
rect 0 77392 800 77512
rect 0 77120 800 77240
rect 0 76848 800 76968
rect 0 76576 800 76696
rect 0 76168 800 76288
rect 0 75896 800 76016
rect 0 75624 800 75744
rect 0 75352 800 75472
rect 179200 75352 180000 75472
rect 0 75080 800 75200
rect 0 74808 800 74928
rect 0 74400 800 74520
rect 0 74128 800 74248
rect 0 73856 800 73976
rect 0 73584 800 73704
rect 0 73312 800 73432
rect 0 73040 800 73160
rect 0 72632 800 72752
rect 0 72360 800 72480
rect 0 72088 800 72208
rect 0 71816 800 71936
rect 0 71544 800 71664
rect 179200 71544 180000 71664
rect 0 71272 800 71392
rect 0 70864 800 70984
rect 0 70592 800 70712
rect 0 70320 800 70440
rect 0 70048 800 70168
rect 0 69776 800 69896
rect 0 69504 800 69624
rect 0 69232 800 69352
rect 0 68824 800 68944
rect 0 68552 800 68672
rect 0 68280 800 68400
rect 0 68008 800 68128
rect 0 67736 800 67856
rect 0 67464 800 67584
rect 179200 67600 180000 67720
rect 0 67056 800 67176
rect 0 66784 800 66904
rect 0 66512 800 66632
rect 0 66240 800 66360
rect 0 65968 800 66088
rect 0 65696 800 65816
rect 0 65288 800 65408
rect 0 65016 800 65136
rect 0 64744 800 64864
rect 0 64472 800 64592
rect 0 64200 800 64320
rect 0 63928 800 64048
rect 179200 63792 180000 63912
rect 0 63520 800 63640
rect 0 63248 800 63368
rect 0 62976 800 63096
rect 0 62704 800 62824
rect 0 62432 800 62552
rect 0 62160 800 62280
rect 0 61752 800 61872
rect 0 61480 800 61600
rect 0 61208 800 61328
rect 0 60936 800 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 0 59712 800 59832
rect 179200 59848 180000 59968
rect 0 59440 800 59560
rect 0 59168 800 59288
rect 0 58896 800 59016
rect 0 58624 800 58744
rect 0 58352 800 58472
rect 0 57944 800 58064
rect 0 57672 800 57792
rect 0 57400 800 57520
rect 0 57128 800 57248
rect 0 56856 800 56976
rect 0 56584 800 56704
rect 0 56176 800 56296
rect 0 55904 800 56024
rect 179200 56040 180000 56160
rect 0 55632 800 55752
rect 0 55360 800 55480
rect 0 55088 800 55208
rect 0 54816 800 54936
rect 0 54408 800 54528
rect 0 54136 800 54256
rect 0 53864 800 53984
rect 0 53592 800 53712
rect 0 53320 800 53440
rect 0 53048 800 53168
rect 0 52640 800 52760
rect 0 52368 800 52488
rect 0 52096 800 52216
rect 179200 52096 180000 52216
rect 0 51824 800 51944
rect 0 51552 800 51672
rect 0 51280 800 51400
rect 0 50872 800 50992
rect 0 50600 800 50720
rect 0 50328 800 50448
rect 0 50056 800 50176
rect 0 49784 800 49904
rect 0 49512 800 49632
rect 0 49240 800 49360
rect 0 48832 800 48952
rect 0 48560 800 48680
rect 0 48288 800 48408
rect 179200 48288 180000 48408
rect 0 48016 800 48136
rect 0 47744 800 47864
rect 0 47472 800 47592
rect 0 47064 800 47184
rect 0 46792 800 46912
rect 0 46520 800 46640
rect 0 46248 800 46368
rect 0 45976 800 46096
rect 0 45704 800 45824
rect 0 45296 800 45416
rect 0 45024 800 45144
rect 0 44752 800 44872
rect 0 44480 800 44600
rect 0 44208 800 44328
rect 179200 44344 180000 44464
rect 0 43936 800 44056
rect 0 43528 800 43648
rect 0 43256 800 43376
rect 0 42984 800 43104
rect 0 42712 800 42832
rect 0 42440 800 42560
rect 0 42168 800 42288
rect 0 41760 800 41880
rect 0 41488 800 41608
rect 0 41216 800 41336
rect 0 40944 800 41064
rect 0 40672 800 40792
rect 0 40400 800 40520
rect 179200 40536 180000 40656
rect 0 40128 800 40248
rect 0 39720 800 39840
rect 0 39448 800 39568
rect 0 39176 800 39296
rect 0 38904 800 39024
rect 0 38632 800 38752
rect 0 38360 800 38480
rect 0 37952 800 38072
rect 0 37680 800 37800
rect 0 37408 800 37528
rect 0 37136 800 37256
rect 0 36864 800 36984
rect 0 36592 800 36712
rect 179200 36728 180000 36848
rect 0 36184 800 36304
rect 0 35912 800 36032
rect 0 35640 800 35760
rect 0 35368 800 35488
rect 0 35096 800 35216
rect 0 34824 800 34944
rect 0 34416 800 34536
rect 0 34144 800 34264
rect 0 33872 800 33992
rect 0 33600 800 33720
rect 0 33328 800 33448
rect 0 33056 800 33176
rect 0 32648 800 32768
rect 179200 32784 180000 32904
rect 0 32376 800 32496
rect 0 32104 800 32224
rect 0 31832 800 31952
rect 0 31560 800 31680
rect 0 31288 800 31408
rect 0 30880 800 31000
rect 0 30608 800 30728
rect 0 30336 800 30456
rect 0 30064 800 30184
rect 0 29792 800 29912
rect 0 29520 800 29640
rect 0 29248 800 29368
rect 0 28840 800 28960
rect 179200 28976 180000 29096
rect 0 28568 800 28688
rect 0 28296 800 28416
rect 0 28024 800 28144
rect 0 27752 800 27872
rect 0 27480 800 27600
rect 0 27072 800 27192
rect 0 26800 800 26920
rect 0 26528 800 26648
rect 0 26256 800 26376
rect 0 25984 800 26104
rect 0 25712 800 25832
rect 0 25304 800 25424
rect 0 25032 800 25152
rect 179200 25032 180000 25152
rect 0 24760 800 24880
rect 0 24488 800 24608
rect 0 24216 800 24336
rect 0 23944 800 24064
rect 0 23536 800 23656
rect 0 23264 800 23384
rect 0 22992 800 23112
rect 0 22720 800 22840
rect 0 22448 800 22568
rect 0 22176 800 22296
rect 0 21768 800 21888
rect 0 21496 800 21616
rect 0 21224 800 21344
rect 179200 21224 180000 21344
rect 0 20952 800 21072
rect 0 20680 800 20800
rect 0 20408 800 20528
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19456 800 19576
rect 0 19184 800 19304
rect 0 18912 800 19032
rect 0 18640 800 18760
rect 0 18368 800 18488
rect 0 17960 800 18080
rect 0 17688 800 17808
rect 0 17416 800 17536
rect 0 17144 800 17264
rect 179200 17280 180000 17400
rect 0 16872 800 16992
rect 0 16600 800 16720
rect 0 16192 800 16312
rect 0 15920 800 16040
rect 0 15648 800 15768
rect 0 15376 800 15496
rect 0 15104 800 15224
rect 0 14832 800 14952
rect 0 14424 800 14544
rect 0 14152 800 14272
rect 0 13880 800 14000
rect 0 13608 800 13728
rect 0 13336 800 13456
rect 179200 13472 180000 13592
rect 0 13064 800 13184
rect 0 12656 800 12776
rect 0 12384 800 12504
rect 0 12112 800 12232
rect 0 11840 800 11960
rect 0 11568 800 11688
rect 0 11296 800 11416
rect 0 10888 800 11008
rect 0 10616 800 10736
rect 0 10344 800 10464
rect 0 10072 800 10192
rect 0 9800 800 9920
rect 0 9528 800 9648
rect 179200 9528 180000 9648
rect 0 9256 800 9376
rect 0 8848 800 8968
rect 0 8576 800 8696
rect 0 8304 800 8424
rect 0 8032 800 8152
rect 0 7760 800 7880
rect 0 7488 800 7608
rect 0 7080 800 7200
rect 0 6808 800 6928
rect 0 6536 800 6656
rect 0 6264 800 6384
rect 0 5992 800 6112
rect 0 5720 800 5840
rect 179200 5720 180000 5840
rect 0 5312 800 5432
rect 0 5040 800 5160
rect 0 4768 800 4888
rect 0 4496 800 4616
rect 0 4224 800 4344
rect 0 3952 800 4072
rect 0 3544 800 3664
rect 0 3272 800 3392
rect 0 3000 800 3120
rect 0 2728 800 2848
rect 0 2456 800 2576
rect 0 2184 800 2304
rect 0 1776 800 1896
rect 179200 1912 180000 2032
rect 0 1504 800 1624
rect 0 1232 800 1352
rect 0 960 800 1080
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
<< obsm3 >>
rect 880 118248 179200 119781
rect 800 118120 179200 118248
rect 880 117840 179120 118120
rect 880 116480 179200 117840
rect 800 116352 179200 116480
rect 880 114712 179200 116352
rect 800 114584 179200 114712
rect 880 114312 179200 114584
rect 880 114032 179120 114312
rect 880 112944 179200 114032
rect 800 112816 179200 112944
rect 880 111176 179200 112816
rect 800 111048 179200 111176
rect 880 110368 179200 111048
rect 880 110088 179120 110368
rect 880 109136 179200 110088
rect 800 109008 179200 109136
rect 880 107368 179200 109008
rect 800 107240 179200 107368
rect 880 106560 179200 107240
rect 880 106280 179120 106560
rect 880 105600 179200 106280
rect 800 105472 179200 105600
rect 880 103832 179200 105472
rect 800 103704 179200 103832
rect 880 102616 179200 103704
rect 880 102336 179120 102616
rect 880 102064 179200 102336
rect 800 101936 179200 102064
rect 880 100024 179200 101936
rect 800 99896 179200 100024
rect 880 98808 179200 99896
rect 880 98528 179120 98808
rect 880 98256 179200 98528
rect 800 98128 179200 98256
rect 880 96488 179200 98128
rect 800 96360 179200 96488
rect 880 94864 179200 96360
rect 880 94720 179120 94864
rect 800 94592 179120 94720
rect 880 94584 179120 94592
rect 880 92952 179200 94584
rect 800 92824 179200 92952
rect 880 91184 179200 92824
rect 800 91056 179200 91184
rect 880 90776 179120 91056
rect 880 89144 179200 90776
rect 800 89016 179200 89144
rect 880 87376 179200 89016
rect 800 87248 179200 87376
rect 880 87112 179200 87248
rect 880 86832 179120 87112
rect 880 85608 179200 86832
rect 800 85480 179200 85608
rect 880 83840 179200 85480
rect 800 83712 179200 83840
rect 880 83304 179200 83712
rect 880 83024 179120 83304
rect 880 82072 179200 83024
rect 800 81944 179200 82072
rect 880 80032 179200 81944
rect 800 79904 179200 80032
rect 880 79496 179200 79904
rect 880 79216 179120 79496
rect 880 78264 179200 79216
rect 800 78136 179200 78264
rect 880 76496 179200 78136
rect 800 76368 179200 76496
rect 880 75552 179200 76368
rect 880 75272 179120 75552
rect 880 74728 179200 75272
rect 800 74600 179200 74728
rect 880 72960 179200 74600
rect 800 72832 179200 72960
rect 880 71744 179200 72832
rect 880 71464 179120 71744
rect 880 71192 179200 71464
rect 800 71064 179200 71192
rect 880 69152 179200 71064
rect 800 69024 179200 69152
rect 880 67800 179200 69024
rect 880 67520 179120 67800
rect 880 67384 179200 67520
rect 800 67256 179200 67384
rect 880 65616 179200 67256
rect 800 65488 179200 65616
rect 880 63992 179200 65488
rect 880 63848 179120 63992
rect 800 63720 179120 63848
rect 880 63712 179120 63720
rect 880 62080 179200 63712
rect 800 61952 179200 62080
rect 880 60048 179200 61952
rect 880 60040 179120 60048
rect 800 59912 179120 60040
rect 880 59768 179120 59912
rect 880 58272 179200 59768
rect 800 58144 179200 58272
rect 880 56504 179200 58144
rect 800 56376 179200 56504
rect 880 56240 179200 56376
rect 880 55960 179120 56240
rect 880 54736 179200 55960
rect 800 54608 179200 54736
rect 880 52968 179200 54608
rect 800 52840 179200 52968
rect 880 52296 179200 52840
rect 880 52016 179120 52296
rect 880 51200 179200 52016
rect 800 51072 179200 51200
rect 880 49160 179200 51072
rect 800 49032 179200 49160
rect 880 48488 179200 49032
rect 880 48208 179120 48488
rect 880 47392 179200 48208
rect 800 47264 179200 47392
rect 880 45624 179200 47264
rect 800 45496 179200 45624
rect 880 44544 179200 45496
rect 880 44264 179120 44544
rect 880 43856 179200 44264
rect 800 43728 179200 43856
rect 880 42088 179200 43728
rect 800 41960 179200 42088
rect 880 40736 179200 41960
rect 880 40456 179120 40736
rect 880 40048 179200 40456
rect 800 39920 179200 40048
rect 880 38280 179200 39920
rect 800 38152 179200 38280
rect 880 36928 179200 38152
rect 880 36648 179120 36928
rect 880 36512 179200 36648
rect 800 36384 179200 36512
rect 880 34744 179200 36384
rect 800 34616 179200 34744
rect 880 32984 179200 34616
rect 880 32976 179120 32984
rect 800 32848 179120 32976
rect 880 32704 179120 32848
rect 880 31208 179200 32704
rect 800 31080 179200 31208
rect 880 29176 179200 31080
rect 880 29168 179120 29176
rect 800 29040 179120 29168
rect 880 28896 179120 29040
rect 880 27400 179200 28896
rect 800 27272 179200 27400
rect 880 25632 179200 27272
rect 800 25504 179200 25632
rect 880 25232 179200 25504
rect 880 24952 179120 25232
rect 880 23864 179200 24952
rect 800 23736 179200 23864
rect 880 22096 179200 23736
rect 800 21968 179200 22096
rect 880 21424 179200 21968
rect 880 21144 179120 21424
rect 880 20056 179200 21144
rect 800 19928 179200 20056
rect 880 18288 179200 19928
rect 800 18160 179200 18288
rect 880 17480 179200 18160
rect 880 17200 179120 17480
rect 880 16520 179200 17200
rect 800 16392 179200 16520
rect 880 14752 179200 16392
rect 800 14624 179200 14752
rect 880 13672 179200 14624
rect 880 13392 179120 13672
rect 880 12984 179200 13392
rect 800 12856 179200 12984
rect 880 11216 179200 12856
rect 800 11088 179200 11216
rect 880 9728 179200 11088
rect 880 9448 179120 9728
rect 880 9176 179200 9448
rect 800 9048 179200 9176
rect 880 7408 179200 9048
rect 800 7280 179200 7408
rect 880 5920 179200 7280
rect 880 5640 179120 5920
rect 800 5512 179200 5640
rect 880 3872 179200 5512
rect 800 3744 179200 3872
rect 880 2112 179200 3744
rect 880 2104 179120 2112
rect 800 1976 179120 2104
rect 880 1832 179120 1976
rect 880 171 179200 1832
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 85534 115907 96288 116789
rect 96768 115907 96948 116789
rect 97428 115907 97608 116789
rect 98088 115907 98268 116789
rect 98748 115907 111648 116789
rect 112128 115907 112308 116789
rect 112788 115907 112968 116789
rect 113448 115907 113628 116789
rect 114108 115907 119994 116789
<< obsm5 >>
rect 85492 116460 120036 116780
<< labels >>
rlabel metal2 s 115662 119200 115718 120000 6 adc_dat_i[0]
port 1 nsew signal input
rlabel metal2 s 124494 119200 124550 120000 6 adc_dat_i[10]
port 2 nsew signal input
rlabel metal2 s 125414 119200 125470 120000 6 adc_dat_i[11]
port 3 nsew signal input
rlabel metal2 s 126242 119200 126298 120000 6 adc_dat_i[12]
port 4 nsew signal input
rlabel metal2 s 127162 119200 127218 120000 6 adc_dat_i[13]
port 5 nsew signal input
rlabel metal2 s 128082 119200 128138 120000 6 adc_dat_i[14]
port 6 nsew signal input
rlabel metal2 s 128910 119200 128966 120000 6 adc_dat_i[15]
port 7 nsew signal input
rlabel metal2 s 129830 119200 129886 120000 6 adc_dat_i[16]
port 8 nsew signal input
rlabel metal2 s 130750 119200 130806 120000 6 adc_dat_i[17]
port 9 nsew signal input
rlabel metal2 s 131578 119200 131634 120000 6 adc_dat_i[18]
port 10 nsew signal input
rlabel metal2 s 132498 119200 132554 120000 6 adc_dat_i[19]
port 11 nsew signal input
rlabel metal2 s 116490 119200 116546 120000 6 adc_dat_i[1]
port 12 nsew signal input
rlabel metal2 s 133418 119200 133474 120000 6 adc_dat_i[20]
port 13 nsew signal input
rlabel metal2 s 134246 119200 134302 120000 6 adc_dat_i[21]
port 14 nsew signal input
rlabel metal2 s 135166 119200 135222 120000 6 adc_dat_i[22]
port 15 nsew signal input
rlabel metal2 s 135994 119200 136050 120000 6 adc_dat_i[23]
port 16 nsew signal input
rlabel metal2 s 136914 119200 136970 120000 6 adc_dat_i[24]
port 17 nsew signal input
rlabel metal2 s 137834 119200 137890 120000 6 adc_dat_i[25]
port 18 nsew signal input
rlabel metal2 s 138662 119200 138718 120000 6 adc_dat_i[26]
port 19 nsew signal input
rlabel metal2 s 139582 119200 139638 120000 6 adc_dat_i[27]
port 20 nsew signal input
rlabel metal2 s 140502 119200 140558 120000 6 adc_dat_i[28]
port 21 nsew signal input
rlabel metal2 s 141330 119200 141386 120000 6 adc_dat_i[29]
port 22 nsew signal input
rlabel metal2 s 117410 119200 117466 120000 6 adc_dat_i[2]
port 23 nsew signal input
rlabel metal2 s 142250 119200 142306 120000 6 adc_dat_i[30]
port 24 nsew signal input
rlabel metal2 s 143170 119200 143226 120000 6 adc_dat_i[31]
port 25 nsew signal input
rlabel metal2 s 118330 119200 118386 120000 6 adc_dat_i[3]
port 26 nsew signal input
rlabel metal2 s 119158 119200 119214 120000 6 adc_dat_i[4]
port 27 nsew signal input
rlabel metal2 s 120078 119200 120134 120000 6 adc_dat_i[5]
port 28 nsew signal input
rlabel metal2 s 120998 119200 121054 120000 6 adc_dat_i[6]
port 29 nsew signal input
rlabel metal2 s 121826 119200 121882 120000 6 adc_dat_i[7]
port 30 nsew signal input
rlabel metal2 s 122746 119200 122802 120000 6 adc_dat_i[8]
port 31 nsew signal input
rlabel metal2 s 123666 119200 123722 120000 6 adc_dat_i[9]
port 32 nsew signal input
rlabel metal2 s 114742 119200 114798 120000 6 adc_dvalid_i
port 33 nsew signal input
rlabel metal2 s 112994 119200 113050 120000 6 adc_sel_o[0]
port 34 nsew signal output
rlabel metal2 s 113822 119200 113878 120000 6 adc_sel_o[1]
port 35 nsew signal output
rlabel metal2 s 386 119200 442 120000 6 io_in[0]
port 36 nsew signal input
rlabel metal2 s 26974 119200 27030 120000 6 io_in[10]
port 37 nsew signal input
rlabel metal2 s 29642 119200 29698 120000 6 io_in[11]
port 38 nsew signal input
rlabel metal2 s 32310 119200 32366 120000 6 io_in[12]
port 39 nsew signal input
rlabel metal2 s 34886 119200 34942 120000 6 io_in[13]
port 40 nsew signal input
rlabel metal2 s 37554 119200 37610 120000 6 io_in[14]
port 41 nsew signal input
rlabel metal2 s 40222 119200 40278 120000 6 io_in[15]
port 42 nsew signal input
rlabel metal2 s 42890 119200 42946 120000 6 io_in[16]
port 43 nsew signal input
rlabel metal2 s 45558 119200 45614 120000 6 io_in[17]
port 44 nsew signal input
rlabel metal2 s 48226 119200 48282 120000 6 io_in[18]
port 45 nsew signal input
rlabel metal2 s 50894 119200 50950 120000 6 io_in[19]
port 46 nsew signal input
rlabel metal2 s 2962 119200 3018 120000 6 io_in[1]
port 47 nsew signal input
rlabel metal2 s 53562 119200 53618 120000 6 io_in[20]
port 48 nsew signal input
rlabel metal2 s 56230 119200 56286 120000 6 io_in[21]
port 49 nsew signal input
rlabel metal2 s 58898 119200 58954 120000 6 io_in[22]
port 50 nsew signal input
rlabel metal2 s 61566 119200 61622 120000 6 io_in[23]
port 51 nsew signal input
rlabel metal2 s 64234 119200 64290 120000 6 io_in[24]
port 52 nsew signal input
rlabel metal2 s 66902 119200 66958 120000 6 io_in[25]
port 53 nsew signal input
rlabel metal2 s 69478 119200 69534 120000 6 io_in[26]
port 54 nsew signal input
rlabel metal2 s 72146 119200 72202 120000 6 io_in[27]
port 55 nsew signal input
rlabel metal2 s 74814 119200 74870 120000 6 io_in[28]
port 56 nsew signal input
rlabel metal2 s 77482 119200 77538 120000 6 io_in[29]
port 57 nsew signal input
rlabel metal2 s 5630 119200 5686 120000 6 io_in[2]
port 58 nsew signal input
rlabel metal2 s 80150 119200 80206 120000 6 io_in[30]
port 59 nsew signal input
rlabel metal2 s 82818 119200 82874 120000 6 io_in[31]
port 60 nsew signal input
rlabel metal2 s 85486 119200 85542 120000 6 io_in[32]
port 61 nsew signal input
rlabel metal2 s 88154 119200 88210 120000 6 io_in[33]
port 62 nsew signal input
rlabel metal2 s 90822 119200 90878 120000 6 io_in[34]
port 63 nsew signal input
rlabel metal2 s 93490 119200 93546 120000 6 io_in[35]
port 64 nsew signal input
rlabel metal2 s 96158 119200 96214 120000 6 io_in[36]
port 65 nsew signal input
rlabel metal2 s 98826 119200 98882 120000 6 io_in[37]
port 66 nsew signal input
rlabel metal2 s 8298 119200 8354 120000 6 io_in[3]
port 67 nsew signal input
rlabel metal2 s 10966 119200 11022 120000 6 io_in[4]
port 68 nsew signal input
rlabel metal2 s 13634 119200 13690 120000 6 io_in[5]
port 69 nsew signal input
rlabel metal2 s 16302 119200 16358 120000 6 io_in[6]
port 70 nsew signal input
rlabel metal2 s 18970 119200 19026 120000 6 io_in[7]
port 71 nsew signal input
rlabel metal2 s 21638 119200 21694 120000 6 io_in[8]
port 72 nsew signal input
rlabel metal2 s 24306 119200 24362 120000 6 io_in[9]
port 73 nsew signal input
rlabel metal2 s 1214 119200 1270 120000 6 io_oeb[0]
port 74 nsew signal output
rlabel metal2 s 27802 119200 27858 120000 6 io_oeb[10]
port 75 nsew signal output
rlabel metal2 s 30470 119200 30526 120000 6 io_oeb[11]
port 76 nsew signal output
rlabel metal2 s 33138 119200 33194 120000 6 io_oeb[12]
port 77 nsew signal output
rlabel metal2 s 35806 119200 35862 120000 6 io_oeb[13]
port 78 nsew signal output
rlabel metal2 s 38474 119200 38530 120000 6 io_oeb[14]
port 79 nsew signal output
rlabel metal2 s 41142 119200 41198 120000 6 io_oeb[15]
port 80 nsew signal output
rlabel metal2 s 43810 119200 43866 120000 6 io_oeb[16]
port 81 nsew signal output
rlabel metal2 s 46478 119200 46534 120000 6 io_oeb[17]
port 82 nsew signal output
rlabel metal2 s 49146 119200 49202 120000 6 io_oeb[18]
port 83 nsew signal output
rlabel metal2 s 51814 119200 51870 120000 6 io_oeb[19]
port 84 nsew signal output
rlabel metal2 s 3882 119200 3938 120000 6 io_oeb[1]
port 85 nsew signal output
rlabel metal2 s 54482 119200 54538 120000 6 io_oeb[20]
port 86 nsew signal output
rlabel metal2 s 57058 119200 57114 120000 6 io_oeb[21]
port 87 nsew signal output
rlabel metal2 s 59726 119200 59782 120000 6 io_oeb[22]
port 88 nsew signal output
rlabel metal2 s 62394 119200 62450 120000 6 io_oeb[23]
port 89 nsew signal output
rlabel metal2 s 65062 119200 65118 120000 6 io_oeb[24]
port 90 nsew signal output
rlabel metal2 s 67730 119200 67786 120000 6 io_oeb[25]
port 91 nsew signal output
rlabel metal2 s 70398 119200 70454 120000 6 io_oeb[26]
port 92 nsew signal output
rlabel metal2 s 73066 119200 73122 120000 6 io_oeb[27]
port 93 nsew signal output
rlabel metal2 s 75734 119200 75790 120000 6 io_oeb[28]
port 94 nsew signal output
rlabel metal2 s 78402 119200 78458 120000 6 io_oeb[29]
port 95 nsew signal output
rlabel metal2 s 6550 119200 6606 120000 6 io_oeb[2]
port 96 nsew signal output
rlabel metal2 s 81070 119200 81126 120000 6 io_oeb[30]
port 97 nsew signal output
rlabel metal2 s 83738 119200 83794 120000 6 io_oeb[31]
port 98 nsew signal output
rlabel metal2 s 86406 119200 86462 120000 6 io_oeb[32]
port 99 nsew signal output
rlabel metal2 s 89074 119200 89130 120000 6 io_oeb[33]
port 100 nsew signal output
rlabel metal2 s 91650 119200 91706 120000 6 io_oeb[34]
port 101 nsew signal output
rlabel metal2 s 94318 119200 94374 120000 6 io_oeb[35]
port 102 nsew signal output
rlabel metal2 s 96986 119200 97042 120000 6 io_oeb[36]
port 103 nsew signal output
rlabel metal2 s 99654 119200 99710 120000 6 io_oeb[37]
port 104 nsew signal output
rlabel metal2 s 9218 119200 9274 120000 6 io_oeb[3]
port 105 nsew signal output
rlabel metal2 s 11886 119200 11942 120000 6 io_oeb[4]
port 106 nsew signal output
rlabel metal2 s 14554 119200 14610 120000 6 io_oeb[5]
port 107 nsew signal output
rlabel metal2 s 17222 119200 17278 120000 6 io_oeb[6]
port 108 nsew signal output
rlabel metal2 s 19890 119200 19946 120000 6 io_oeb[7]
port 109 nsew signal output
rlabel metal2 s 22558 119200 22614 120000 6 io_oeb[8]
port 110 nsew signal output
rlabel metal2 s 25134 119200 25190 120000 6 io_oeb[9]
port 111 nsew signal output
rlabel metal2 s 2134 119200 2190 120000 6 io_out[0]
port 112 nsew signal output
rlabel metal2 s 28722 119200 28778 120000 6 io_out[10]
port 113 nsew signal output
rlabel metal2 s 31390 119200 31446 120000 6 io_out[11]
port 114 nsew signal output
rlabel metal2 s 34058 119200 34114 120000 6 io_out[12]
port 115 nsew signal output
rlabel metal2 s 36726 119200 36782 120000 6 io_out[13]
port 116 nsew signal output
rlabel metal2 s 39394 119200 39450 120000 6 io_out[14]
port 117 nsew signal output
rlabel metal2 s 42062 119200 42118 120000 6 io_out[15]
port 118 nsew signal output
rlabel metal2 s 44730 119200 44786 120000 6 io_out[16]
port 119 nsew signal output
rlabel metal2 s 47306 119200 47362 120000 6 io_out[17]
port 120 nsew signal output
rlabel metal2 s 49974 119200 50030 120000 6 io_out[18]
port 121 nsew signal output
rlabel metal2 s 52642 119200 52698 120000 6 io_out[19]
port 122 nsew signal output
rlabel metal2 s 4802 119200 4858 120000 6 io_out[1]
port 123 nsew signal output
rlabel metal2 s 55310 119200 55366 120000 6 io_out[20]
port 124 nsew signal output
rlabel metal2 s 57978 119200 58034 120000 6 io_out[21]
port 125 nsew signal output
rlabel metal2 s 60646 119200 60702 120000 6 io_out[22]
port 126 nsew signal output
rlabel metal2 s 63314 119200 63370 120000 6 io_out[23]
port 127 nsew signal output
rlabel metal2 s 65982 119200 66038 120000 6 io_out[24]
port 128 nsew signal output
rlabel metal2 s 68650 119200 68706 120000 6 io_out[25]
port 129 nsew signal output
rlabel metal2 s 71318 119200 71374 120000 6 io_out[26]
port 130 nsew signal output
rlabel metal2 s 73986 119200 74042 120000 6 io_out[27]
port 131 nsew signal output
rlabel metal2 s 76654 119200 76710 120000 6 io_out[28]
port 132 nsew signal output
rlabel metal2 s 79230 119200 79286 120000 6 io_out[29]
port 133 nsew signal output
rlabel metal2 s 7470 119200 7526 120000 6 io_out[2]
port 134 nsew signal output
rlabel metal2 s 81898 119200 81954 120000 6 io_out[30]
port 135 nsew signal output
rlabel metal2 s 84566 119200 84622 120000 6 io_out[31]
port 136 nsew signal output
rlabel metal2 s 87234 119200 87290 120000 6 io_out[32]
port 137 nsew signal output
rlabel metal2 s 89902 119200 89958 120000 6 io_out[33]
port 138 nsew signal output
rlabel metal2 s 92570 119200 92626 120000 6 io_out[34]
port 139 nsew signal output
rlabel metal2 s 95238 119200 95294 120000 6 io_out[35]
port 140 nsew signal output
rlabel metal2 s 97906 119200 97962 120000 6 io_out[36]
port 141 nsew signal output
rlabel metal2 s 100574 119200 100630 120000 6 io_out[37]
port 142 nsew signal output
rlabel metal2 s 10138 119200 10194 120000 6 io_out[3]
port 143 nsew signal output
rlabel metal2 s 12714 119200 12770 120000 6 io_out[4]
port 144 nsew signal output
rlabel metal2 s 15382 119200 15438 120000 6 io_out[5]
port 145 nsew signal output
rlabel metal2 s 18050 119200 18106 120000 6 io_out[6]
port 146 nsew signal output
rlabel metal2 s 20718 119200 20774 120000 6 io_out[7]
port 147 nsew signal output
rlabel metal2 s 23386 119200 23442 120000 6 io_out[8]
port 148 nsew signal output
rlabel metal2 s 26054 119200 26110 120000 6 io_out[9]
port 149 nsew signal output
rlabel metal3 s 179200 1912 180000 2032 6 irq[0]
port 150 nsew signal output
rlabel metal2 s 149334 119200 149390 120000 6 irq[1]
port 151 nsew signal output
rlabel metal3 s 179200 9528 180000 9648 6 irq[2]
port 152 nsew signal output
rlabel metal3 s 0 144 800 264 6 la_data_in[0]
port 153 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 la_data_in[100]
port 154 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 la_data_in[101]
port 155 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 la_data_in[102]
port 156 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 la_data_in[103]
port 157 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 la_data_in[104]
port 158 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 la_data_in[105]
port 159 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 la_data_in[106]
port 160 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 la_data_in[107]
port 161 nsew signal input
rlabel metal3 s 0 95344 800 95464 6 la_data_in[108]
port 162 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 la_data_in[109]
port 163 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_data_in[10]
port 164 nsew signal input
rlabel metal3 s 0 97112 800 97232 6 la_data_in[110]
port 165 nsew signal input
rlabel metal3 s 0 97928 800 98048 6 la_data_in[111]
port 166 nsew signal input
rlabel metal3 s 0 98880 800 99000 6 la_data_in[112]
port 167 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 la_data_in[113]
port 168 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 la_data_in[114]
port 169 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 la_data_in[115]
port 170 nsew signal input
rlabel metal3 s 0 102416 800 102536 6 la_data_in[116]
port 171 nsew signal input
rlabel metal3 s 0 103232 800 103352 6 la_data_in[117]
port 172 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 la_data_in[118]
port 173 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 la_data_in[119]
port 174 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 la_data_in[11]
port 175 nsew signal input
rlabel metal3 s 0 105952 800 106072 6 la_data_in[120]
port 176 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 la_data_in[121]
port 177 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 la_data_in[122]
port 178 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 la_data_in[123]
port 179 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 la_data_in[124]
port 180 nsew signal input
rlabel metal3 s 0 110304 800 110424 6 la_data_in[125]
port 181 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 la_data_in[126]
port 182 nsew signal input
rlabel metal3 s 0 112072 800 112192 6 la_data_in[127]
port 183 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 la_data_in[12]
port 184 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_data_in[13]
port 185 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 la_data_in[14]
port 186 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 la_data_in[15]
port 187 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 la_data_in[16]
port 188 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 la_data_in[17]
port 189 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 la_data_in[18]
port 190 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 la_data_in[19]
port 191 nsew signal input
rlabel metal3 s 0 960 800 1080 6 la_data_in[1]
port 192 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 la_data_in[20]
port 193 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 la_data_in[21]
port 194 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 la_data_in[22]
port 195 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_data_in[23]
port 196 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 la_data_in[24]
port 197 nsew signal input
rlabel metal3 s 0 22176 800 22296 6 la_data_in[25]
port 198 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 la_data_in[26]
port 199 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 la_data_in[27]
port 200 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 la_data_in[28]
port 201 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 la_data_in[29]
port 202 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 la_data_in[2]
port 203 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 la_data_in[30]
port 204 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 la_data_in[31]
port 205 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 la_data_in[32]
port 206 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 la_data_in[33]
port 207 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 la_data_in[34]
port 208 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 la_data_in[35]
port 209 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 la_data_in[36]
port 210 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la_data_in[37]
port 211 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 la_data_in[38]
port 212 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 la_data_in[39]
port 213 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_data_in[3]
port 214 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 la_data_in[40]
port 215 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 la_data_in[41]
port 216 nsew signal input
rlabel metal3 s 0 37136 800 37256 6 la_data_in[42]
port 217 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 la_data_in[43]
port 218 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 la_data_in[44]
port 219 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 la_data_in[45]
port 220 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 la_data_in[46]
port 221 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 la_data_in[47]
port 222 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 la_data_in[48]
port 223 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 la_data_in[49]
port 224 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 la_data_in[4]
port 225 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 la_data_in[50]
port 226 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 la_data_in[51]
port 227 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 la_data_in[52]
port 228 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 la_data_in[53]
port 229 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 la_data_in[54]
port 230 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 la_data_in[55]
port 231 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 la_data_in[56]
port 232 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 la_data_in[57]
port 233 nsew signal input
rlabel metal3 s 0 51280 800 51400 6 la_data_in[58]
port 234 nsew signal input
rlabel metal3 s 0 52096 800 52216 6 la_data_in[59]
port 235 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 la_data_in[5]
port 236 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 la_data_in[60]
port 237 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 la_data_in[61]
port 238 nsew signal input
rlabel metal3 s 0 54816 800 54936 6 la_data_in[62]
port 239 nsew signal input
rlabel metal3 s 0 55632 800 55752 6 la_data_in[63]
port 240 nsew signal input
rlabel metal3 s 0 56584 800 56704 6 la_data_in[64]
port 241 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 la_data_in[65]
port 242 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 la_data_in[66]
port 243 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_data_in[67]
port 244 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 la_data_in[68]
port 245 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 la_data_in[69]
port 246 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 la_data_in[6]
port 247 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 la_data_in[70]
port 248 nsew signal input
rlabel metal3 s 0 62704 800 62824 6 la_data_in[71]
port 249 nsew signal input
rlabel metal3 s 0 63520 800 63640 6 la_data_in[72]
port 250 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 la_data_in[73]
port 251 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 la_data_in[74]
port 252 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 la_data_in[75]
port 253 nsew signal input
rlabel metal3 s 0 67056 800 67176 6 la_data_in[76]
port 254 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 la_data_in[77]
port 255 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 la_data_in[78]
port 256 nsew signal input
rlabel metal3 s 0 69776 800 69896 6 la_data_in[79]
port 257 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 la_data_in[7]
port 258 nsew signal input
rlabel metal3 s 0 70592 800 70712 6 la_data_in[80]
port 259 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 la_data_in[81]
port 260 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 la_data_in[82]
port 261 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 la_data_in[83]
port 262 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_data_in[84]
port 263 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 la_data_in[85]
port 264 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 la_data_in[86]
port 265 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 la_data_in[87]
port 266 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 la_data_in[88]
port 267 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 la_data_in[89]
port 268 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 la_data_in[8]
port 269 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 la_data_in[90]
port 270 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 la_data_in[91]
port 271 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 la_data_in[92]
port 272 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 la_data_in[93]
port 273 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 la_data_in[94]
port 274 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 la_data_in[95]
port 275 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 la_data_in[96]
port 276 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 la_data_in[97]
port 277 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 la_data_in[98]
port 278 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 la_data_in[99]
port 279 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 la_data_in[9]
port 280 nsew signal input
rlabel metal3 s 0 416 800 536 6 la_data_out[0]
port 281 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 la_data_out[100]
port 282 nsew signal output
rlabel metal3 s 0 89496 800 89616 6 la_data_out[101]
port 283 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 la_data_out[102]
port 284 nsew signal output
rlabel metal3 s 0 91264 800 91384 6 la_data_out[103]
port 285 nsew signal output
rlabel metal3 s 0 92080 800 92200 6 la_data_out[104]
port 286 nsew signal output
rlabel metal3 s 0 93032 800 93152 6 la_data_out[105]
port 287 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 la_data_out[106]
port 288 nsew signal output
rlabel metal3 s 0 94800 800 94920 6 la_data_out[107]
port 289 nsew signal output
rlabel metal3 s 0 95616 800 95736 6 la_data_out[108]
port 290 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 la_data_out[109]
port 291 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 la_data_out[10]
port 292 nsew signal output
rlabel metal3 s 0 97384 800 97504 6 la_data_out[110]
port 293 nsew signal output
rlabel metal3 s 0 98336 800 98456 6 la_data_out[111]
port 294 nsew signal output
rlabel metal3 s 0 99152 800 99272 6 la_data_out[112]
port 295 nsew signal output
rlabel metal3 s 0 100104 800 100224 6 la_data_out[113]
port 296 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 la_data_out[114]
port 297 nsew signal output
rlabel metal3 s 0 101736 800 101856 6 la_data_out[115]
port 298 nsew signal output
rlabel metal3 s 0 102688 800 102808 6 la_data_out[116]
port 299 nsew signal output
rlabel metal3 s 0 103504 800 103624 6 la_data_out[117]
port 300 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 la_data_out[118]
port 301 nsew signal output
rlabel metal3 s 0 105272 800 105392 6 la_data_out[119]
port 302 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 la_data_out[11]
port 303 nsew signal output
rlabel metal3 s 0 106224 800 106344 6 la_data_out[120]
port 304 nsew signal output
rlabel metal3 s 0 107040 800 107160 6 la_data_out[121]
port 305 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 la_data_out[122]
port 306 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 la_data_out[123]
port 307 nsew signal output
rlabel metal3 s 0 109760 800 109880 6 la_data_out[124]
port 308 nsew signal output
rlabel metal3 s 0 110576 800 110696 6 la_data_out[125]
port 309 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 la_data_out[126]
port 310 nsew signal output
rlabel metal3 s 0 112344 800 112464 6 la_data_out[127]
port 311 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 la_data_out[12]
port 312 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 la_data_out[13]
port 313 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 la_data_out[14]
port 314 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 la_data_out[15]
port 315 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 la_data_out[16]
port 316 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 la_data_out[17]
port 317 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 la_data_out[18]
port 318 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 la_data_out[19]
port 319 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 la_data_out[1]
port 320 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 la_data_out[20]
port 321 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 la_data_out[21]
port 322 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[22]
port 323 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 la_data_out[23]
port 324 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 la_data_out[24]
port 325 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 la_data_out[25]
port 326 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 la_data_out[26]
port 327 nsew signal output
rlabel metal3 s 0 24216 800 24336 6 la_data_out[27]
port 328 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 la_data_out[28]
port 329 nsew signal output
rlabel metal3 s 0 25984 800 26104 6 la_data_out[29]
port 330 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 la_data_out[2]
port 331 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 la_data_out[30]
port 332 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 la_data_out[31]
port 333 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 la_data_out[32]
port 334 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 la_data_out[33]
port 335 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 la_data_out[34]
port 336 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 la_data_out[35]
port 337 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 la_data_out[36]
port 338 nsew signal output
rlabel metal3 s 0 33056 800 33176 6 la_data_out[37]
port 339 nsew signal output
rlabel metal3 s 0 33872 800 33992 6 la_data_out[38]
port 340 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 la_data_out[39]
port 341 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 la_data_out[3]
port 342 nsew signal output
rlabel metal3 s 0 35640 800 35760 6 la_data_out[40]
port 343 nsew signal output
rlabel metal3 s 0 36592 800 36712 6 la_data_out[41]
port 344 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 la_data_out[42]
port 345 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 la_data_out[43]
port 346 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 la_data_out[44]
port 347 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 la_data_out[45]
port 348 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 la_data_out[46]
port 349 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 la_data_out[47]
port 350 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 la_data_out[48]
port 351 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 la_data_out[49]
port 352 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 la_data_out[4]
port 353 nsew signal output
rlabel metal3 s 0 44480 800 44600 6 la_data_out[50]
port 354 nsew signal output
rlabel metal3 s 0 45296 800 45416 6 la_data_out[51]
port 355 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 la_data_out[52]
port 356 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 la_data_out[53]
port 357 nsew signal output
rlabel metal3 s 0 48016 800 48136 6 la_data_out[54]
port 358 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 la_data_out[55]
port 359 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 la_data_out[56]
port 360 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 la_data_out[57]
port 361 nsew signal output
rlabel metal3 s 0 51552 800 51672 6 la_data_out[58]
port 362 nsew signal output
rlabel metal3 s 0 52368 800 52488 6 la_data_out[59]
port 363 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 la_data_out[5]
port 364 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 la_data_out[60]
port 365 nsew signal output
rlabel metal3 s 0 54136 800 54256 6 la_data_out[61]
port 366 nsew signal output
rlabel metal3 s 0 55088 800 55208 6 la_data_out[62]
port 367 nsew signal output
rlabel metal3 s 0 55904 800 56024 6 la_data_out[63]
port 368 nsew signal output
rlabel metal3 s 0 56856 800 56976 6 la_data_out[64]
port 369 nsew signal output
rlabel metal3 s 0 57672 800 57792 6 la_data_out[65]
port 370 nsew signal output
rlabel metal3 s 0 58624 800 58744 6 la_data_out[66]
port 371 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 la_data_out[67]
port 372 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 la_data_out[68]
port 373 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 la_data_out[69]
port 374 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 la_data_out[6]
port 375 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 la_data_out[70]
port 376 nsew signal output
rlabel metal3 s 0 62976 800 63096 6 la_data_out[71]
port 377 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 la_data_out[72]
port 378 nsew signal output
rlabel metal3 s 0 64744 800 64864 6 la_data_out[73]
port 379 nsew signal output
rlabel metal3 s 0 65696 800 65816 6 la_data_out[74]
port 380 nsew signal output
rlabel metal3 s 0 66512 800 66632 6 la_data_out[75]
port 381 nsew signal output
rlabel metal3 s 0 67464 800 67584 6 la_data_out[76]
port 382 nsew signal output
rlabel metal3 s 0 68280 800 68400 6 la_data_out[77]
port 383 nsew signal output
rlabel metal3 s 0 69232 800 69352 6 la_data_out[78]
port 384 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 la_data_out[79]
port 385 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 la_data_out[7]
port 386 nsew signal output
rlabel metal3 s 0 70864 800 70984 6 la_data_out[80]
port 387 nsew signal output
rlabel metal3 s 0 71816 800 71936 6 la_data_out[81]
port 388 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 la_data_out[82]
port 389 nsew signal output
rlabel metal3 s 0 73584 800 73704 6 la_data_out[83]
port 390 nsew signal output
rlabel metal3 s 0 74400 800 74520 6 la_data_out[84]
port 391 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 la_data_out[85]
port 392 nsew signal output
rlabel metal3 s 0 76168 800 76288 6 la_data_out[86]
port 393 nsew signal output
rlabel metal3 s 0 77120 800 77240 6 la_data_out[87]
port 394 nsew signal output
rlabel metal3 s 0 77936 800 78056 6 la_data_out[88]
port 395 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 la_data_out[89]
port 396 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 la_data_out[8]
port 397 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 la_data_out[90]
port 398 nsew signal output
rlabel metal3 s 0 80656 800 80776 6 la_data_out[91]
port 399 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 la_data_out[92]
port 400 nsew signal output
rlabel metal3 s 0 82424 800 82544 6 la_data_out[93]
port 401 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 la_data_out[94]
port 402 nsew signal output
rlabel metal3 s 0 84192 800 84312 6 la_data_out[95]
port 403 nsew signal output
rlabel metal3 s 0 85008 800 85128 6 la_data_out[96]
port 404 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 la_data_out[97]
port 405 nsew signal output
rlabel metal3 s 0 86776 800 86896 6 la_data_out[98]
port 406 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 la_data_out[99]
port 407 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 la_data_out[9]
port 408 nsew signal output
rlabel metal3 s 0 688 800 808 6 la_oenb[0]
port 409 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 la_oenb[100]
port 410 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 la_oenb[101]
port 411 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 la_oenb[102]
port 412 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 la_oenb[103]
port 413 nsew signal input
rlabel metal3 s 0 92352 800 92472 6 la_oenb[104]
port 414 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 la_oenb[105]
port 415 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 la_oenb[106]
port 416 nsew signal input
rlabel metal3 s 0 95072 800 95192 6 la_oenb[107]
port 417 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 la_oenb[108]
port 418 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 la_oenb[109]
port 419 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 la_oenb[10]
port 420 nsew signal input
rlabel metal3 s 0 97656 800 97776 6 la_oenb[110]
port 421 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 la_oenb[111]
port 422 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 la_oenb[112]
port 423 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 la_oenb[113]
port 424 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 la_oenb[114]
port 425 nsew signal input
rlabel metal3 s 0 102144 800 102264 6 la_oenb[115]
port 426 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 la_oenb[116]
port 427 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 la_oenb[117]
port 428 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_oenb[118]
port 429 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 la_oenb[119]
port 430 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 la_oenb[11]
port 431 nsew signal input
rlabel metal3 s 0 106496 800 106616 6 la_oenb[120]
port 432 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 la_oenb[121]
port 433 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 la_oenb[122]
port 434 nsew signal input
rlabel metal3 s 0 109216 800 109336 6 la_oenb[123]
port 435 nsew signal input
rlabel metal3 s 0 110032 800 110152 6 la_oenb[124]
port 436 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 la_oenb[125]
port 437 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 la_oenb[126]
port 438 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 la_oenb[127]
port 439 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 la_oenb[12]
port 440 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 la_oenb[13]
port 441 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 la_oenb[14]
port 442 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 la_oenb[15]
port 443 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 la_oenb[16]
port 444 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_oenb[17]
port 445 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 la_oenb[18]
port 446 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 la_oenb[19]
port 447 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 la_oenb[1]
port 448 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 la_oenb[20]
port 449 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 la_oenb[21]
port 450 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 la_oenb[22]
port 451 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 la_oenb[23]
port 452 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 la_oenb[24]
port 453 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 la_oenb[25]
port 454 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 la_oenb[26]
port 455 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 la_oenb[27]
port 456 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 la_oenb[28]
port 457 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 la_oenb[29]
port 458 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 la_oenb[2]
port 459 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 la_oenb[30]
port 460 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 la_oenb[31]
port 461 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 la_oenb[32]
port 462 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 la_oenb[33]
port 463 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 la_oenb[34]
port 464 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 la_oenb[35]
port 465 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 la_oenb[36]
port 466 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 la_oenb[37]
port 467 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 la_oenb[38]
port 468 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 la_oenb[39]
port 469 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 la_oenb[3]
port 470 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 la_oenb[40]
port 471 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 la_oenb[41]
port 472 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 la_oenb[42]
port 473 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 la_oenb[43]
port 474 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_oenb[44]
port 475 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 la_oenb[45]
port 476 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 la_oenb[46]
port 477 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 la_oenb[47]
port 478 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 la_oenb[48]
port 479 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 la_oenb[49]
port 480 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 la_oenb[4]
port 481 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 la_oenb[50]
port 482 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 la_oenb[51]
port 483 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 la_oenb[52]
port 484 nsew signal input
rlabel metal3 s 0 47472 800 47592 6 la_oenb[53]
port 485 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 la_oenb[54]
port 486 nsew signal input
rlabel metal3 s 0 49240 800 49360 6 la_oenb[55]
port 487 nsew signal input
rlabel metal3 s 0 50056 800 50176 6 la_oenb[56]
port 488 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 la_oenb[57]
port 489 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 la_oenb[58]
port 490 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 la_oenb[59]
port 491 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 la_oenb[5]
port 492 nsew signal input
rlabel metal3 s 0 53592 800 53712 6 la_oenb[60]
port 493 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_oenb[61]
port 494 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 la_oenb[62]
port 495 nsew signal input
rlabel metal3 s 0 56176 800 56296 6 la_oenb[63]
port 496 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 la_oenb[64]
port 497 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 la_oenb[65]
port 498 nsew signal input
rlabel metal3 s 0 58896 800 59016 6 la_oenb[66]
port 499 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 la_oenb[67]
port 500 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 la_oenb[68]
port 501 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 la_oenb[69]
port 502 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 la_oenb[6]
port 503 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 la_oenb[70]
port 504 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_oenb[71]
port 505 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 la_oenb[72]
port 506 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 la_oenb[73]
port 507 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 la_oenb[74]
port 508 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 la_oenb[75]
port 509 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 la_oenb[76]
port 510 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 la_oenb[77]
port 511 nsew signal input
rlabel metal3 s 0 69504 800 69624 6 la_oenb[78]
port 512 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 la_oenb[79]
port 513 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_oenb[7]
port 514 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 la_oenb[80]
port 515 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 la_oenb[81]
port 516 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 la_oenb[82]
port 517 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 la_oenb[83]
port 518 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 la_oenb[84]
port 519 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 la_oenb[85]
port 520 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 la_oenb[86]
port 521 nsew signal input
rlabel metal3 s 0 77392 800 77512 6 la_oenb[87]
port 522 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 la_oenb[88]
port 523 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 la_oenb[89]
port 524 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 la_oenb[8]
port 525 nsew signal input
rlabel metal3 s 0 80112 800 80232 6 la_oenb[90]
port 526 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 la_oenb[91]
port 527 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 la_oenb[92]
port 528 nsew signal input
rlabel metal3 s 0 82696 800 82816 6 la_oenb[93]
port 529 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 la_oenb[94]
port 530 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 la_oenb[95]
port 531 nsew signal input
rlabel metal3 s 0 85280 800 85400 6 la_oenb[96]
port 532 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 la_oenb[97]
port 533 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 la_oenb[98]
port 534 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 la_oenb[99]
port 535 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 la_oenb[9]
port 536 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 mem1_data_i[0]
port 537 nsew signal input
rlabel metal2 s 157430 0 157486 800 6 mem1_data_i[10]
port 538 nsew signal input
rlabel metal3 s 179200 71544 180000 71664 6 mem1_data_i[11]
port 539 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 mem1_data_i[12]
port 540 nsew signal input
rlabel metal3 s 179200 75352 180000 75472 6 mem1_data_i[13]
port 541 nsew signal input
rlabel metal3 s 0 117376 800 117496 6 mem1_data_i[14]
port 542 nsew signal input
rlabel metal2 s 161754 119200 161810 120000 6 mem1_data_i[15]
port 543 nsew signal input
rlabel metal2 s 165158 0 165214 800 6 mem1_data_i[16]
port 544 nsew signal input
rlabel metal2 s 165342 119200 165398 120000 6 mem1_data_i[17]
port 545 nsew signal input
rlabel metal2 s 166446 0 166502 800 6 mem1_data_i[18]
port 546 nsew signal input
rlabel metal3 s 0 118600 800 118720 6 mem1_data_i[19]
port 547 nsew signal input
rlabel metal2 s 150254 119200 150310 120000 6 mem1_data_i[1]
port 548 nsew signal input
rlabel metal2 s 168838 119200 168894 120000 6 mem1_data_i[20]
port 549 nsew signal input
rlabel metal3 s 179200 83104 180000 83224 6 mem1_data_i[21]
port 550 nsew signal input
rlabel metal3 s 179200 86912 180000 87032 6 mem1_data_i[22]
port 551 nsew signal input
rlabel metal2 s 171506 119200 171562 120000 6 mem1_data_i[23]
port 552 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 mem1_data_i[24]
port 553 nsew signal input
rlabel metal3 s 179200 98608 180000 98728 6 mem1_data_i[25]
port 554 nsew signal input
rlabel metal2 s 175094 119200 175150 120000 6 mem1_data_i[26]
port 555 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 mem1_data_i[27]
port 556 nsew signal input
rlabel metal3 s 179200 110168 180000 110288 6 mem1_data_i[28]
port 557 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 mem1_data_i[29]
port 558 nsew signal input
rlabel metal2 s 144550 0 144606 800 6 mem1_data_i[2]
port 559 nsew signal input
rlabel metal2 s 176842 119200 176898 120000 6 mem1_data_i[30]
port 560 nsew signal input
rlabel metal2 s 178590 119200 178646 120000 6 mem1_data_i[31]
port 561 nsew signal input
rlabel metal3 s 179200 25032 180000 25152 6 mem1_data_i[3]
port 562 nsew signal input
rlabel metal2 s 154670 119200 154726 120000 6 mem1_data_i[4]
port 563 nsew signal input
rlabel metal3 s 179200 44344 180000 44464 6 mem1_data_i[5]
port 564 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 mem1_data_i[6]
port 565 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 mem1_data_i[7]
port 566 nsew signal input
rlabel metal3 s 179200 63792 180000 63912 6 mem1_data_i[8]
port 567 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 mem1_data_i[9]
port 568 nsew signal input
rlabel metal2 s 138110 0 138166 800 6 mem_data2_i[0]
port 569 nsew signal input
rlabel metal2 s 158718 0 158774 800 6 mem_data2_i[10]
port 570 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 mem_data2_i[11]
port 571 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 mem_data2_i[12]
port 572 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 mem_data2_i[13]
port 573 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 mem_data2_i[14]
port 574 nsew signal input
rlabel metal2 s 162674 119200 162730 120000 6 mem_data2_i[15]
port 575 nsew signal input
rlabel metal2 s 163502 119200 163558 120000 6 mem_data2_i[16]
port 576 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 mem_data2_i[17]
port 577 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 mem_data2_i[18]
port 578 nsew signal input
rlabel metal2 s 167734 0 167790 800 6 mem_data2_i[19]
port 579 nsew signal input
rlabel metal3 s 0 113024 800 113144 6 mem_data2_i[1]
port 580 nsew signal input
rlabel metal2 s 169758 119200 169814 120000 6 mem_data2_i[20]
port 581 nsew signal input
rlabel metal2 s 170586 119200 170642 120000 6 mem_data2_i[21]
port 582 nsew signal input
rlabel metal3 s 179200 90856 180000 90976 6 mem_data2_i[22]
port 583 nsew signal input
rlabel metal2 s 172426 119200 172482 120000 6 mem_data2_i[23]
port 584 nsew signal input
rlabel metal2 s 174174 119200 174230 120000 6 mem_data2_i[24]
port 585 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 mem_data2_i[25]
port 586 nsew signal input
rlabel metal2 s 172886 0 172942 800 6 mem_data2_i[26]
port 587 nsew signal input
rlabel metal2 s 175922 119200 175978 120000 6 mem_data2_i[27]
port 588 nsew signal input
rlabel metal2 s 175462 0 175518 800 6 mem_data2_i[28]
port 589 nsew signal input
rlabel metal3 s 179200 117920 180000 118040 6 mem_data2_i[29]
port 590 nsew signal input
rlabel metal2 s 145838 0 145894 800 6 mem_data2_i[2]
port 591 nsew signal input
rlabel metal2 s 178038 0 178094 800 6 mem_data2_i[30]
port 592 nsew signal input
rlabel metal2 s 179510 119200 179566 120000 6 mem_data2_i[31]
port 593 nsew signal input
rlabel metal3 s 179200 28976 180000 29096 6 mem_data2_i[3]
port 594 nsew signal input
rlabel metal3 s 179200 36728 180000 36848 6 mem_data2_i[4]
port 595 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 mem_data2_i[5]
port 596 nsew signal input
rlabel metal2 s 156418 119200 156474 120000 6 mem_data2_i[6]
port 597 nsew signal input
rlabel metal3 s 179200 52096 180000 52216 6 mem_data2_i[7]
port 598 nsew signal input
rlabel metal2 s 157338 119200 157394 120000 6 mem_data2_i[8]
port 599 nsew signal input
rlabel metal2 s 160006 119200 160062 120000 6 mem_data2_i[9]
port 600 nsew signal input
rlabel metal2 s 146666 119200 146722 120000 6 mem_data_i[0]
port 601 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 mem_data_i[10]
port 602 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 mem_data_i[11]
port 603 nsew signal input
rlabel metal3 s 0 116832 800 116952 6 mem_data_i[12]
port 604 nsew signal input
rlabel metal3 s 179200 79296 180000 79416 6 mem_data_i[13]
port 605 nsew signal input
rlabel metal2 s 163870 0 163926 800 6 mem_data_i[14]
port 606 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 mem_data_i[15]
port 607 nsew signal input
rlabel metal2 s 164422 119200 164478 120000 6 mem_data_i[16]
port 608 nsew signal input
rlabel metal2 s 166170 119200 166226 120000 6 mem_data_i[17]
port 609 nsew signal input
rlabel metal2 s 167090 119200 167146 120000 6 mem_data_i[18]
port 610 nsew signal input
rlabel metal2 s 168010 119200 168066 120000 6 mem_data_i[19]
port 611 nsew signal input
rlabel metal2 s 141974 0 142030 800 6 mem_data_i[1]
port 612 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 mem_data_i[20]
port 613 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 mem_data_i[21]
port 614 nsew signal input
rlabel metal3 s 179200 94664 180000 94784 6 mem_data_i[22]
port 615 nsew signal input
rlabel metal2 s 173254 119200 173310 120000 6 mem_data_i[23]
port 616 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 mem_data_i[24]
port 617 nsew signal input
rlabel metal2 s 171598 0 171654 800 6 mem_data_i[25]
port 618 nsew signal input
rlabel metal3 s 179200 102416 180000 102536 6 mem_data_i[26]
port 619 nsew signal input
rlabel metal3 s 179200 106360 180000 106480 6 mem_data_i[27]
port 620 nsew signal input
rlabel metal3 s 179200 114112 180000 114232 6 mem_data_i[28]
port 621 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 mem_data_i[29]
port 622 nsew signal input
rlabel metal3 s 179200 13472 180000 13592 6 mem_data_i[2]
port 623 nsew signal input
rlabel metal2 s 177762 119200 177818 120000 6 mem_data_i[30]
port 624 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 mem_data_i[31]
port 625 nsew signal input
rlabel metal3 s 179200 32784 180000 32904 6 mem_data_i[3]
port 626 nsew signal input
rlabel metal3 s 179200 40536 180000 40656 6 mem_data_i[4]
port 627 nsew signal input
rlabel metal2 s 155590 119200 155646 120000 6 mem_data_i[5]
port 628 nsew signal input
rlabel metal2 s 152278 0 152334 800 6 mem_data_i[6]
port 629 nsew signal input
rlabel metal3 s 0 115336 800 115456 6 mem_data_i[7]
port 630 nsew signal input
rlabel metal2 s 154854 0 154910 800 6 mem_data_i[8]
port 631 nsew signal input
rlabel metal3 s 179200 67600 180000 67720 6 mem_data_i[9]
port 632 nsew signal input
rlabel metal3 s 179200 5720 180000 5840 6 mem_raddr_o[0]
port 633 nsew signal output
rlabel metal2 s 151082 119200 151138 120000 6 mem_raddr_o[1]
port 634 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 mem_raddr_o[2]
port 635 nsew signal output
rlabel metal2 s 153750 119200 153806 120000 6 mem_raddr_o[3]
port 636 nsew signal output
rlabel metal2 s 148414 0 148470 800 6 mem_raddr_o[4]
port 637 nsew signal output
rlabel metal3 s 179200 48288 180000 48408 6 mem_raddr_o[5]
port 638 nsew signal output
rlabel metal2 s 153566 0 153622 800 6 mem_raddr_o[6]
port 639 nsew signal output
rlabel metal3 s 179200 56040 180000 56160 6 mem_raddr_o[7]
port 640 nsew signal output
rlabel metal2 s 158166 119200 158222 120000 6 mem_raddr_o[8]
port 641 nsew signal output
rlabel metal2 s 160834 119200 160890 120000 6 mem_raddr_o[9]
port 642 nsew signal output
rlabel metal2 s 147586 119200 147642 120000 6 mem_renb_o[0]
port 643 nsew signal output
rlabel metal2 s 152002 119200 152058 120000 6 mem_renb_o[1]
port 644 nsew signal output
rlabel metal2 s 148414 119200 148470 120000 6 mem_waddr_o[0]
port 645 nsew signal output
rlabel metal2 s 143262 0 143318 800 6 mem_waddr_o[1]
port 646 nsew signal output
rlabel metal3 s 179200 17280 180000 17400 6 mem_waddr_o[2]
port 647 nsew signal output
rlabel metal3 s 0 113840 800 113960 6 mem_waddr_o[3]
port 648 nsew signal output
rlabel metal3 s 0 114112 800 114232 6 mem_waddr_o[4]
port 649 nsew signal output
rlabel metal2 s 149702 0 149758 800 6 mem_waddr_o[5]
port 650 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 mem_waddr_o[6]
port 651 nsew signal output
rlabel metal3 s 179200 59848 180000 59968 6 mem_waddr_o[7]
port 652 nsew signal output
rlabel metal2 s 159086 119200 159142 120000 6 mem_waddr_o[8]
port 653 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 mem_waddr_o[9]
port 654 nsew signal output
rlabel metal2 s 139398 0 139454 800 6 mem_wenb_o[0]
port 655 nsew signal output
rlabel metal2 s 152922 119200 152978 120000 6 mem_wenb_o[1]
port 656 nsew signal output
rlabel metal2 s 101494 119200 101550 120000 6 oversample_o[0]
port 657 nsew signal output
rlabel metal2 s 102322 119200 102378 120000 6 oversample_o[1]
port 658 nsew signal output
rlabel metal2 s 103242 119200 103298 120000 6 oversample_o[2]
port 659 nsew signal output
rlabel metal2 s 104070 119200 104126 120000 6 oversample_o[3]
port 660 nsew signal output
rlabel metal2 s 104990 119200 105046 120000 6 oversample_o[4]
port 661 nsew signal output
rlabel metal2 s 105910 119200 105966 120000 6 oversample_o[5]
port 662 nsew signal output
rlabel metal2 s 106738 119200 106794 120000 6 oversample_o[6]
port 663 nsew signal output
rlabel metal2 s 107658 119200 107714 120000 6 oversample_o[7]
port 664 nsew signal output
rlabel metal2 s 108578 119200 108634 120000 6 oversample_o[8]
port 665 nsew signal output
rlabel metal2 s 109406 119200 109462 120000 6 oversample_o[9]
port 666 nsew signal output
rlabel metal2 s 110326 119200 110382 120000 6 sinc3_en_o[0]
port 667 nsew signal output
rlabel metal2 s 111246 119200 111302 120000 6 sinc3_en_o[1]
port 668 nsew signal output
rlabel metal2 s 112074 119200 112130 120000 6 sinc3_en_o[2]
port 669 nsew signal output
rlabel metal2 s 143998 119200 144054 120000 6 vco_enb_o[0]
port 670 nsew signal output
rlabel metal2 s 144918 119200 144974 120000 6 vco_enb_o[1]
port 671 nsew signal output
rlabel metal2 s 145838 119200 145894 120000 6 vco_enb_o[2]
port 672 nsew signal output
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 673 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wb_rst_i
port 674 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_ack_o
port 675 nsew signal output
rlabel metal2 s 8206 0 8262 800 6 wbs_adr_i[0]
port 676 nsew signal input
rlabel metal2 s 51998 0 52054 800 6 wbs_adr_i[10]
port 677 nsew signal input
rlabel metal2 s 55862 0 55918 800 6 wbs_adr_i[11]
port 678 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_adr_i[12]
port 679 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 wbs_adr_i[13]
port 680 nsew signal input
rlabel metal2 s 67362 0 67418 800 6 wbs_adr_i[14]
port 681 nsew signal input
rlabel metal2 s 71226 0 71282 800 6 wbs_adr_i[15]
port 682 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 wbs_adr_i[16]
port 683 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_adr_i[17]
port 684 nsew signal input
rlabel metal2 s 82818 0 82874 800 6 wbs_adr_i[18]
port 685 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 wbs_adr_i[19]
port 686 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wbs_adr_i[1]
port 687 nsew signal input
rlabel metal2 s 90546 0 90602 800 6 wbs_adr_i[20]
port 688 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 wbs_adr_i[21]
port 689 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 wbs_adr_i[22]
port 690 nsew signal input
rlabel metal2 s 102138 0 102194 800 6 wbs_adr_i[23]
port 691 nsew signal input
rlabel metal2 s 106002 0 106058 800 6 wbs_adr_i[24]
port 692 nsew signal input
rlabel metal2 s 109866 0 109922 800 6 wbs_adr_i[25]
port 693 nsew signal input
rlabel metal2 s 113730 0 113786 800 6 wbs_adr_i[26]
port 694 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 wbs_adr_i[27]
port 695 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 wbs_adr_i[28]
port 696 nsew signal input
rlabel metal2 s 125230 0 125286 800 6 wbs_adr_i[29]
port 697 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 wbs_adr_i[2]
port 698 nsew signal input
rlabel metal2 s 129094 0 129150 800 6 wbs_adr_i[30]
port 699 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 wbs_adr_i[31]
port 700 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 wbs_adr_i[3]
port 701 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_adr_i[4]
port 702 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wbs_adr_i[5]
port 703 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wbs_adr_i[6]
port 704 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 wbs_adr_i[7]
port 705 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_adr_i[8]
port 706 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 wbs_adr_i[9]
port 707 nsew signal input
rlabel metal2 s 4342 0 4398 800 6 wbs_cyc_i
port 708 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wbs_dat_i[0]
port 709 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 wbs_dat_i[10]
port 710 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 wbs_dat_i[11]
port 711 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 wbs_dat_i[12]
port 712 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_i[13]
port 713 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 wbs_dat_i[14]
port 714 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 wbs_dat_i[15]
port 715 nsew signal input
rlabel metal2 s 76378 0 76434 800 6 wbs_dat_i[16]
port 716 nsew signal input
rlabel metal2 s 80242 0 80298 800 6 wbs_dat_i[17]
port 717 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 wbs_dat_i[18]
port 718 nsew signal input
rlabel metal2 s 87970 0 88026 800 6 wbs_dat_i[19]
port 719 nsew signal input
rlabel metal2 s 14646 0 14702 800 6 wbs_dat_i[1]
port 720 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 wbs_dat_i[20]
port 721 nsew signal input
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_i[21]
port 722 nsew signal input
rlabel metal2 s 99562 0 99618 800 6 wbs_dat_i[22]
port 723 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 wbs_dat_i[23]
port 724 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 wbs_dat_i[24]
port 725 nsew signal input
rlabel metal2 s 111154 0 111210 800 6 wbs_dat_i[25]
port 726 nsew signal input
rlabel metal2 s 115018 0 115074 800 6 wbs_dat_i[26]
port 727 nsew signal input
rlabel metal2 s 118882 0 118938 800 6 wbs_dat_i[27]
port 728 nsew signal input
rlabel metal2 s 122654 0 122710 800 6 wbs_dat_i[28]
port 729 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_i[29]
port 730 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_i[2]
port 731 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 wbs_dat_i[30]
port 732 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 wbs_dat_i[31]
port 733 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[3]
port 734 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 wbs_dat_i[4]
port 735 nsew signal input
rlabel metal2 s 33966 0 34022 800 6 wbs_dat_i[5]
port 736 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_dat_i[6]
port 737 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 wbs_dat_i[7]
port 738 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_i[8]
port 739 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 wbs_dat_i[9]
port 740 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_o[0]
port 741 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 wbs_dat_o[10]
port 742 nsew signal output
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_o[11]
port 743 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 wbs_dat_o[12]
port 744 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 wbs_dat_o[13]
port 745 nsew signal output
rlabel metal2 s 69938 0 69994 800 6 wbs_dat_o[14]
port 746 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 wbs_dat_o[15]
port 747 nsew signal output
rlabel metal2 s 77666 0 77722 800 6 wbs_dat_o[16]
port 748 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_o[17]
port 749 nsew signal output
rlabel metal2 s 85394 0 85450 800 6 wbs_dat_o[18]
port 750 nsew signal output
rlabel metal2 s 89258 0 89314 800 6 wbs_dat_o[19]
port 751 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_o[1]
port 752 nsew signal output
rlabel metal2 s 93122 0 93178 800 6 wbs_dat_o[20]
port 753 nsew signal output
rlabel metal2 s 96986 0 97042 800 6 wbs_dat_o[21]
port 754 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 wbs_dat_o[22]
port 755 nsew signal output
rlabel metal2 s 104714 0 104770 800 6 wbs_dat_o[23]
port 756 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 wbs_dat_o[24]
port 757 nsew signal output
rlabel metal2 s 112442 0 112498 800 6 wbs_dat_o[25]
port 758 nsew signal output
rlabel metal2 s 116306 0 116362 800 6 wbs_dat_o[26]
port 759 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 wbs_dat_o[27]
port 760 nsew signal output
rlabel metal2 s 123942 0 123998 800 6 wbs_dat_o[28]
port 761 nsew signal output
rlabel metal2 s 127806 0 127862 800 6 wbs_dat_o[29]
port 762 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_o[2]
port 763 nsew signal output
rlabel metal2 s 131670 0 131726 800 6 wbs_dat_o[30]
port 764 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 wbs_dat_o[31]
port 765 nsew signal output
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_o[3]
port 766 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 wbs_dat_o[4]
port 767 nsew signal output
rlabel metal2 s 35254 0 35310 800 6 wbs_dat_o[5]
port 768 nsew signal output
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_o[6]
port 769 nsew signal output
rlabel metal2 s 42982 0 43038 800 6 wbs_dat_o[7]
port 770 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_o[8]
port 771 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 wbs_dat_o[9]
port 772 nsew signal output
rlabel metal2 s 12070 0 12126 800 6 wbs_sel_i[0]
port 773 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_sel_i[1]
port 774 nsew signal input
rlabel metal2 s 22374 0 22430 800 6 wbs_sel_i[2]
port 775 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_sel_i[3]
port 776 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_stb_i
port 777 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_we_i
port 778 nsew signal input
rlabel metal2 s 140686 0 140742 800 6 wmask_o[0]
port 779 nsew signal output
rlabel metal3 s 0 113296 800 113416 6 wmask_o[1]
port 780 nsew signal output
rlabel metal3 s 179200 21224 180000 21344 6 wmask_o[2]
port 781 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 wmask_o[3]
port 782 nsew signal output
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 783 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 784 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 785 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 786 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 787 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 788 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 789 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 790 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 791 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 792 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 793 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 794 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 795 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 796 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 797 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 798 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 799 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 800 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 801 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 802 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 803 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 804 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 805 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 806 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 807 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 808 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 809 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 810 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 811 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 812 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 813 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 814 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 815 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 816 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 817 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 818 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 819 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 820 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 821 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 822 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 823 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 824 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 825 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 826 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 827 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 828 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 829 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 830 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 8835230
string GDS_START 598470
<< end >>

