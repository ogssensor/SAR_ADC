VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ring_osc_3-1
  CLASS BLOCK ;
  FOREIGN ring_osc_3-1 ;
  ORIGIN 0.000 1.290 ;
  SIZE 181.500 BY 40.660 ;
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 133.300 9.880 134.500 10.460 ;
        RECT 132.500 9.760 134.500 9.880 ;
        RECT 151.270 9.820 152.450 10.100 ;
        RECT 132.500 9.160 136.500 9.760 ;
        RECT 150.770 9.220 152.450 9.820 ;
        RECT 151.270 9.020 152.450 9.220 ;
        RECT 154.935 8.730 155.435 9.880 ;
        RECT 157.450 8.730 157.745 12.995 ;
        RECT 164.600 10.460 164.890 15.790 ;
        RECT 168.780 10.460 169.070 15.790 ;
        RECT 164.600 10.170 169.070 10.460 ;
        RECT 167.030 8.730 167.530 10.170 ;
        RECT 154.935 8.230 167.530 8.730 ;
        RECT 157.455 0.550 157.750 8.230 ;
        RECT 164.600 3.230 164.890 8.230 ;
      LAYER mcon ;
        RECT 132.560 9.220 133.200 9.850 ;
        RECT 133.400 9.160 134.100 9.850 ;
        RECT 134.300 9.160 134.900 9.760 ;
        RECT 135.100 9.160 135.700 9.760 ;
        RECT 135.900 9.160 136.500 9.760 ;
        RECT 150.820 9.270 151.220 9.770 ;
        RECT 151.420 9.270 152.370 9.770 ;
        RECT 154.935 9.220 155.435 9.820 ;
      LAYER met1 ;
        RECT 132.500 9.820 136.600 9.880 ;
        RECT 154.905 9.820 155.465 9.880 ;
        RECT 132.500 9.220 155.465 9.820 ;
        RECT 132.500 9.160 136.600 9.220 ;
        RECT 154.905 9.160 155.465 9.220 ;
        RECT 133.300 9.130 136.600 9.160 ;
      LAYER via ;
        RECT 149.000 9.220 149.600 9.820 ;
        RECT 149.740 9.220 150.340 9.820 ;
      LAYER met2 ;
        RECT 149.000 9.190 150.340 9.870 ;
        RECT 149.270 -1.290 150.070 9.190 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 103.800 9.880 105.000 10.460 ;
        RECT 103.000 9.760 105.000 9.880 ;
        RECT 121.770 9.820 122.950 10.100 ;
        RECT 103.000 9.160 107.000 9.760 ;
        RECT 121.270 9.220 122.950 9.820 ;
        RECT 121.770 9.020 122.950 9.220 ;
        RECT 125.435 8.730 125.935 9.880 ;
        RECT 127.950 8.730 128.245 12.995 ;
        RECT 135.100 10.460 135.390 15.790 ;
        RECT 139.280 10.460 139.570 15.790 ;
        RECT 135.100 10.170 139.570 10.460 ;
        RECT 137.530 8.730 138.030 10.170 ;
        RECT 125.435 8.230 138.030 8.730 ;
        RECT 127.955 0.550 128.250 8.230 ;
        RECT 135.100 3.230 135.390 8.230 ;
      LAYER mcon ;
        RECT 103.060 9.220 103.700 9.850 ;
        RECT 103.900 9.160 104.600 9.850 ;
        RECT 104.800 9.160 105.400 9.760 ;
        RECT 105.600 9.160 106.200 9.760 ;
        RECT 106.400 9.160 107.000 9.760 ;
        RECT 121.320 9.270 121.720 9.770 ;
        RECT 121.920 9.270 122.870 9.770 ;
        RECT 125.435 9.220 125.935 9.820 ;
      LAYER met1 ;
        RECT 103.000 9.820 107.100 9.880 ;
        RECT 125.405 9.820 125.965 9.880 ;
        RECT 103.000 9.220 125.965 9.820 ;
        RECT 103.000 9.160 107.100 9.220 ;
        RECT 125.405 9.160 125.965 9.220 ;
        RECT 103.800 9.130 107.100 9.160 ;
      LAYER via ;
        RECT 119.500 9.220 120.100 9.820 ;
        RECT 120.240 9.220 120.840 9.820 ;
      LAYER met2 ;
        RECT 119.500 9.190 120.840 9.870 ;
        RECT 119.770 -1.290 120.570 9.190 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 74.300 9.880 75.500 10.460 ;
        RECT 73.500 9.760 75.500 9.880 ;
        RECT 92.270 9.820 93.450 10.100 ;
        RECT 73.500 9.160 77.500 9.760 ;
        RECT 91.770 9.220 93.450 9.820 ;
        RECT 92.270 9.020 93.450 9.220 ;
        RECT 95.935 8.730 96.435 9.880 ;
        RECT 98.450 8.730 98.745 12.995 ;
        RECT 105.600 10.460 105.890 15.790 ;
        RECT 109.780 10.460 110.070 15.790 ;
        RECT 105.600 10.170 110.070 10.460 ;
        RECT 108.030 8.730 108.530 10.170 ;
        RECT 95.935 8.230 108.530 8.730 ;
        RECT 98.455 0.550 98.750 8.230 ;
        RECT 105.600 3.230 105.890 8.230 ;
      LAYER mcon ;
        RECT 73.560 9.220 74.200 9.850 ;
        RECT 74.400 9.160 75.100 9.850 ;
        RECT 75.300 9.160 75.900 9.760 ;
        RECT 76.100 9.160 76.700 9.760 ;
        RECT 76.900 9.160 77.500 9.760 ;
        RECT 91.820 9.270 92.220 9.770 ;
        RECT 92.420 9.270 93.370 9.770 ;
        RECT 95.935 9.220 96.435 9.820 ;
      LAYER met1 ;
        RECT 73.500 9.820 77.600 9.880 ;
        RECT 95.905 9.820 96.465 9.880 ;
        RECT 73.500 9.220 96.465 9.820 ;
        RECT 73.500 9.160 77.600 9.220 ;
        RECT 95.905 9.160 96.465 9.220 ;
        RECT 74.300 9.130 77.600 9.160 ;
      LAYER via ;
        RECT 90.000 9.220 90.600 9.820 ;
        RECT 90.740 9.220 91.340 9.820 ;
      LAYER met2 ;
        RECT 90.000 9.190 91.340 9.870 ;
        RECT 90.270 -1.290 91.070 9.190 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 44.800 9.880 46.000 10.460 ;
        RECT 44.000 9.760 46.000 9.880 ;
        RECT 62.770 9.820 63.950 10.100 ;
        RECT 44.000 9.160 48.000 9.760 ;
        RECT 62.270 9.220 63.950 9.820 ;
        RECT 62.770 9.020 63.950 9.220 ;
        RECT 66.435 8.730 66.935 9.880 ;
        RECT 68.950 8.730 69.245 12.995 ;
        RECT 76.100 10.460 76.390 15.790 ;
        RECT 80.280 10.460 80.570 15.790 ;
        RECT 76.100 10.170 80.570 10.460 ;
        RECT 78.530 8.730 79.030 10.170 ;
        RECT 66.435 8.230 79.030 8.730 ;
        RECT 68.955 0.550 69.250 8.230 ;
        RECT 76.100 3.230 76.390 8.230 ;
      LAYER mcon ;
        RECT 44.060 9.220 44.700 9.850 ;
        RECT 44.900 9.160 45.600 9.850 ;
        RECT 45.800 9.160 46.400 9.760 ;
        RECT 46.600 9.160 47.200 9.760 ;
        RECT 47.400 9.160 48.000 9.760 ;
        RECT 62.320 9.270 62.720 9.770 ;
        RECT 62.920 9.270 63.870 9.770 ;
        RECT 66.435 9.220 66.935 9.820 ;
      LAYER met1 ;
        RECT 44.000 9.820 48.100 9.880 ;
        RECT 66.405 9.820 66.965 9.880 ;
        RECT 44.000 9.220 66.965 9.820 ;
        RECT 44.000 9.160 48.100 9.220 ;
        RECT 66.405 9.160 66.965 9.220 ;
        RECT 44.800 9.130 48.100 9.160 ;
      LAYER via ;
        RECT 60.500 9.220 61.100 9.820 ;
        RECT 61.240 9.220 61.840 9.820 ;
      LAYER met2 ;
        RECT 60.500 9.190 61.840 9.870 ;
        RECT 60.770 -1.290 61.570 9.190 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 15.300 9.880 16.500 10.460 ;
        RECT 14.500 9.760 16.500 9.880 ;
        RECT 33.270 9.820 34.450 10.100 ;
        RECT 14.500 9.160 18.500 9.760 ;
        RECT 32.770 9.220 34.450 9.820 ;
        RECT 33.270 9.020 34.450 9.220 ;
        RECT 36.935 8.730 37.435 9.880 ;
        RECT 39.450 8.730 39.745 12.995 ;
        RECT 46.600 10.460 46.890 15.790 ;
        RECT 50.780 10.460 51.070 15.790 ;
        RECT 46.600 10.170 51.070 10.460 ;
        RECT 49.030 8.730 49.530 10.170 ;
        RECT 36.935 8.230 49.530 8.730 ;
        RECT 39.455 0.550 39.750 8.230 ;
        RECT 46.600 3.230 46.890 8.230 ;
      LAYER mcon ;
        RECT 14.560 9.220 15.200 9.850 ;
        RECT 15.400 9.160 16.100 9.850 ;
        RECT 16.300 9.160 16.900 9.760 ;
        RECT 17.100 9.160 17.700 9.760 ;
        RECT 17.900 9.160 18.500 9.760 ;
        RECT 32.820 9.270 33.220 9.770 ;
        RECT 33.420 9.270 34.370 9.770 ;
        RECT 36.935 9.220 37.435 9.820 ;
      LAYER met1 ;
        RECT 14.500 9.820 18.600 9.880 ;
        RECT 36.905 9.820 37.465 9.880 ;
        RECT 14.500 9.220 37.465 9.820 ;
        RECT 14.500 9.160 18.600 9.220 ;
        RECT 36.905 9.160 37.465 9.220 ;
        RECT 15.300 9.130 18.600 9.160 ;
      LAYER via ;
        RECT 31.000 9.220 31.600 9.820 ;
        RECT 31.740 9.220 32.340 9.820 ;
      LAYER met2 ;
        RECT 31.000 9.190 32.340 9.870 ;
        RECT 31.270 -1.290 32.070 9.190 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 30.890 28.320 34.890 28.920 ;
        RECT 32.890 28.200 34.890 28.320 ;
        RECT 32.890 27.620 34.090 28.200 ;
        RECT 3.770 9.820 4.950 10.100 ;
        RECT 3.270 9.220 4.950 9.820 ;
        RECT 3.770 9.020 4.950 9.220 ;
        RECT 7.435 8.730 7.935 9.880 ;
        RECT 9.950 8.730 10.245 12.995 ;
        RECT 17.100 10.460 17.390 15.790 ;
        RECT 21.280 10.460 21.570 15.790 ;
        RECT 17.100 10.170 21.570 10.460 ;
        RECT 19.530 8.730 20.030 10.170 ;
        RECT 7.435 8.230 20.030 8.730 ;
        RECT 9.955 0.550 10.250 8.230 ;
        RECT 17.100 3.230 17.390 8.230 ;
      LAYER mcon ;
        RECT 30.890 28.320 31.490 28.920 ;
        RECT 31.690 28.320 32.290 28.920 ;
        RECT 32.490 28.320 33.090 28.920 ;
        RECT 33.290 28.230 33.990 28.920 ;
        RECT 34.190 28.230 34.830 28.860 ;
        RECT 3.320 9.270 3.720 9.770 ;
        RECT 3.920 9.270 4.870 9.770 ;
        RECT 7.435 9.220 7.935 9.820 ;
      LAYER met1 ;
        RECT 30.790 28.920 34.090 28.950 ;
        RECT 30.790 28.860 34.890 28.920 ;
        RECT 17.840 28.260 34.890 28.860 ;
        RECT 30.790 28.200 34.890 28.260 ;
        RECT 7.405 9.820 7.965 9.880 ;
        RECT 2.000 9.220 7.965 9.820 ;
        RECT 7.405 9.160 7.965 9.220 ;
      LAYER via ;
        RECT 17.890 28.260 18.865 28.860 ;
        RECT 6.705 9.220 7.405 9.820 ;
      LAYER met2 ;
        RECT 17.120 28.210 18.865 28.910 ;
        RECT 17.120 17.350 17.820 28.210 ;
        RECT 6.705 16.650 17.820 17.350 ;
        RECT 6.705 9.170 7.405 16.650 ;
        RECT 13.270 -1.290 14.070 16.650 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 32.000 29.850 32.290 34.850 ;
        RECT 39.140 29.850 39.435 37.530 ;
        RECT 29.360 29.350 41.955 29.850 ;
        RECT 29.360 27.910 29.860 29.350 ;
        RECT 27.820 27.620 32.290 27.910 ;
        RECT 27.820 22.290 28.110 27.620 ;
        RECT 32.000 22.290 32.290 27.620 ;
        RECT 39.145 25.085 39.440 29.350 ;
        RECT 41.455 28.200 41.955 29.350 ;
        RECT 44.440 28.860 45.620 29.060 ;
        RECT 44.440 28.260 46.120 28.860 ;
        RECT 60.390 28.320 64.390 28.920 ;
        RECT 44.440 27.980 45.620 28.260 ;
        RECT 62.390 28.200 64.390 28.320 ;
        RECT 62.390 27.620 63.590 28.200 ;
      LAYER mcon ;
        RECT 41.455 28.260 41.955 28.860 ;
        RECT 44.520 28.310 45.470 28.810 ;
        RECT 45.670 28.310 46.070 28.810 ;
        RECT 60.390 28.320 60.990 28.920 ;
        RECT 61.190 28.320 61.790 28.920 ;
        RECT 61.990 28.320 62.590 28.920 ;
        RECT 62.790 28.230 63.490 28.920 ;
        RECT 63.690 28.230 64.330 28.860 ;
      LAYER met1 ;
        RECT 60.290 28.920 63.590 28.950 ;
        RECT 41.425 28.860 41.985 28.920 ;
        RECT 60.290 28.860 64.390 28.920 ;
        RECT 41.425 28.260 64.390 28.860 ;
        RECT 41.425 28.200 41.985 28.260 ;
        RECT 60.290 28.200 64.390 28.260 ;
      LAYER via ;
        RECT 46.550 28.260 47.150 28.860 ;
        RECT 47.290 28.260 47.890 28.860 ;
      LAYER met2 ;
        RECT 46.820 28.920 47.620 39.370 ;
        RECT 46.550 28.210 47.890 28.920 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 61.500 29.850 61.790 34.850 ;
        RECT 68.640 29.850 68.935 37.530 ;
        RECT 58.860 29.350 71.455 29.850 ;
        RECT 58.860 27.910 59.360 29.350 ;
        RECT 57.320 27.620 61.790 27.910 ;
        RECT 57.320 22.290 57.610 27.620 ;
        RECT 61.500 22.290 61.790 27.620 ;
        RECT 68.645 25.085 68.940 29.350 ;
        RECT 70.955 28.200 71.455 29.350 ;
        RECT 73.940 28.860 75.120 29.060 ;
        RECT 73.940 28.260 75.620 28.860 ;
        RECT 89.890 28.320 93.890 28.920 ;
        RECT 73.940 27.980 75.120 28.260 ;
        RECT 91.890 28.200 93.890 28.320 ;
        RECT 91.890 27.620 93.090 28.200 ;
      LAYER mcon ;
        RECT 70.955 28.260 71.455 28.860 ;
        RECT 74.020 28.310 74.970 28.810 ;
        RECT 75.170 28.310 75.570 28.810 ;
        RECT 89.890 28.320 90.490 28.920 ;
        RECT 90.690 28.320 91.290 28.920 ;
        RECT 91.490 28.320 92.090 28.920 ;
        RECT 92.290 28.230 92.990 28.920 ;
        RECT 93.190 28.230 93.830 28.860 ;
      LAYER met1 ;
        RECT 89.790 28.920 93.090 28.950 ;
        RECT 70.925 28.860 71.485 28.920 ;
        RECT 89.790 28.860 93.890 28.920 ;
        RECT 70.925 28.260 93.890 28.860 ;
        RECT 70.925 28.200 71.485 28.260 ;
        RECT 89.790 28.200 93.890 28.260 ;
      LAYER via ;
        RECT 76.050 28.260 76.650 28.860 ;
        RECT 76.790 28.260 77.390 28.860 ;
      LAYER met2 ;
        RECT 76.320 28.920 77.120 39.370 ;
        RECT 76.050 28.210 77.390 28.920 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 91.000 29.850 91.290 34.850 ;
        RECT 98.140 29.850 98.435 37.530 ;
        RECT 88.360 29.350 100.955 29.850 ;
        RECT 88.360 27.910 88.860 29.350 ;
        RECT 86.820 27.620 91.290 27.910 ;
        RECT 86.820 22.290 87.110 27.620 ;
        RECT 91.000 22.290 91.290 27.620 ;
        RECT 98.145 25.085 98.440 29.350 ;
        RECT 100.455 28.200 100.955 29.350 ;
        RECT 103.440 28.860 104.620 29.060 ;
        RECT 103.440 28.260 105.120 28.860 ;
        RECT 119.390 28.320 123.390 28.920 ;
        RECT 103.440 27.980 104.620 28.260 ;
        RECT 121.390 28.200 123.390 28.320 ;
        RECT 121.390 27.620 122.590 28.200 ;
      LAYER mcon ;
        RECT 100.455 28.260 100.955 28.860 ;
        RECT 103.520 28.310 104.470 28.810 ;
        RECT 104.670 28.310 105.070 28.810 ;
        RECT 119.390 28.320 119.990 28.920 ;
        RECT 120.190 28.320 120.790 28.920 ;
        RECT 120.990 28.320 121.590 28.920 ;
        RECT 121.790 28.230 122.490 28.920 ;
        RECT 122.690 28.230 123.330 28.860 ;
      LAYER met1 ;
        RECT 119.290 28.920 122.590 28.950 ;
        RECT 100.425 28.860 100.985 28.920 ;
        RECT 119.290 28.860 123.390 28.920 ;
        RECT 100.425 28.260 123.390 28.860 ;
        RECT 100.425 28.200 100.985 28.260 ;
        RECT 119.290 28.200 123.390 28.260 ;
      LAYER via ;
        RECT 105.550 28.260 106.150 28.860 ;
        RECT 106.290 28.260 106.890 28.860 ;
      LAYER met2 ;
        RECT 105.820 28.920 106.620 39.370 ;
        RECT 105.550 28.210 106.890 28.920 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 120.500 29.850 120.790 34.850 ;
        RECT 127.640 29.850 127.935 37.530 ;
        RECT 117.860 29.350 130.455 29.850 ;
        RECT 117.860 27.910 118.360 29.350 ;
        RECT 116.320 27.620 120.790 27.910 ;
        RECT 116.320 22.290 116.610 27.620 ;
        RECT 120.500 22.290 120.790 27.620 ;
        RECT 127.645 25.085 127.940 29.350 ;
        RECT 129.955 28.200 130.455 29.350 ;
        RECT 132.940 28.860 134.120 29.060 ;
        RECT 132.940 28.260 134.620 28.860 ;
        RECT 148.890 28.320 152.890 28.920 ;
        RECT 132.940 27.980 134.120 28.260 ;
        RECT 150.890 28.200 152.890 28.320 ;
        RECT 150.890 27.620 152.090 28.200 ;
      LAYER mcon ;
        RECT 129.955 28.260 130.455 28.860 ;
        RECT 133.020 28.310 133.970 28.810 ;
        RECT 134.170 28.310 134.570 28.810 ;
        RECT 148.890 28.320 149.490 28.920 ;
        RECT 149.690 28.320 150.290 28.920 ;
        RECT 150.490 28.320 151.090 28.920 ;
        RECT 151.290 28.230 151.990 28.920 ;
        RECT 152.190 28.230 152.830 28.860 ;
      LAYER met1 ;
        RECT 148.790 28.920 152.090 28.950 ;
        RECT 129.925 28.860 130.485 28.920 ;
        RECT 148.790 28.860 152.890 28.920 ;
        RECT 129.925 28.260 152.890 28.860 ;
        RECT 129.925 28.200 130.485 28.260 ;
        RECT 148.790 28.200 152.890 28.260 ;
      LAYER via ;
        RECT 135.050 28.260 135.650 28.860 ;
        RECT 135.790 28.260 136.390 28.860 ;
      LAYER met2 ;
        RECT 135.320 28.920 136.120 39.370 ;
        RECT 135.050 28.210 136.390 28.920 ;
    END
  END p[9]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 150.000 29.850 150.290 34.850 ;
        RECT 157.140 29.850 157.435 37.530 ;
        RECT 147.360 29.350 159.955 29.850 ;
        RECT 147.360 27.910 147.860 29.350 ;
        RECT 145.820 27.620 150.290 27.910 ;
        RECT 145.820 22.290 146.110 27.620 ;
        RECT 150.000 22.290 150.290 27.620 ;
        RECT 157.145 25.085 157.440 29.350 ;
        RECT 159.455 28.200 159.955 29.350 ;
        RECT 162.440 28.860 163.620 29.060 ;
        RECT 162.440 28.260 164.120 28.860 ;
        RECT 162.440 27.980 163.620 28.260 ;
        RECT 162.800 9.880 164.000 10.460 ;
        RECT 162.000 9.760 164.000 9.880 ;
        RECT 162.000 9.160 166.000 9.760 ;
      LAYER mcon ;
        RECT 159.455 28.260 159.955 28.860 ;
        RECT 162.520 28.310 163.470 28.810 ;
        RECT 163.670 28.310 164.070 28.810 ;
        RECT 162.060 9.220 162.700 9.850 ;
        RECT 162.900 9.160 163.600 9.850 ;
        RECT 163.800 9.160 164.400 9.760 ;
        RECT 164.600 9.160 165.200 9.760 ;
        RECT 165.400 9.160 166.000 9.760 ;
      LAYER met1 ;
        RECT 159.425 28.860 159.985 28.920 ;
        RECT 159.425 28.260 165.440 28.860 ;
        RECT 159.425 28.200 159.985 28.260 ;
        RECT 162.000 9.820 166.100 9.880 ;
        RECT 162.000 9.220 179.000 9.820 ;
        RECT 162.000 9.160 166.100 9.220 ;
        RECT 162.800 9.130 166.100 9.160 ;
      LAYER via ;
        RECT 164.450 28.260 165.390 28.860 ;
        RECT 166.090 9.220 166.790 9.820 ;
        RECT 166.860 9.220 167.460 9.820 ;
      LAYER met2 ;
        RECT 164.450 28.210 166.790 28.910 ;
        RECT 166.090 9.870 166.790 28.210 ;
        RECT 166.090 9.140 167.460 9.870 ;
        RECT 166.360 -1.290 167.160 9.140 ;
    END
  END p[10]
  PIN input_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 175.550 25.740 177.550 25.910 ;
        RECT 175.630 25.710 177.470 25.740 ;
      LAYER met1 ;
        RECT 175.520 25.680 177.580 25.940 ;
      LAYER via ;
        RECT 175.570 25.680 177.530 25.940 ;
      LAYER met2 ;
        RECT 175.570 25.390 181.500 26.190 ;
        RECT 176.150 25.200 177.530 25.390 ;
    END
  END input_analog
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 2.790 2.495 6.550 7.770 ;
        RECT 14.320 2.445 20.170 8.300 ;
        RECT 32.290 2.495 36.050 7.770 ;
        RECT 43.820 2.445 49.670 8.300 ;
        RECT 61.790 2.495 65.550 7.770 ;
        RECT 73.320 2.445 79.170 8.300 ;
        RECT 91.290 2.495 95.050 7.770 ;
        RECT 102.820 2.445 108.670 8.300 ;
        RECT 120.790 2.495 124.550 7.770 ;
        RECT 132.320 2.445 138.170 8.300 ;
        RECT 150.290 2.495 154.050 7.770 ;
        RECT 161.820 2.445 167.670 8.300 ;
      LAYER li1 ;
        RECT 2.970 2.960 3.140 7.375 ;
        RECT 3.480 2.960 3.770 7.370 ;
        RECT 2.970 2.930 5.065 2.960 ;
        RECT 2.970 2.845 5.220 2.930 ;
        RECT 6.200 2.845 6.370 5.820 ;
        RECT 2.970 2.675 6.370 2.845 ;
        RECT 14.500 2.960 14.670 7.560 ;
        RECT 15.010 2.960 15.300 7.790 ;
        RECT 19.190 2.960 19.480 7.790 ;
        RECT 19.820 2.960 19.990 7.620 ;
        RECT 14.500 2.795 16.845 2.960 ;
        RECT 17.645 2.795 19.990 2.960 ;
        RECT 2.970 2.510 5.220 2.675 ;
        RECT 14.500 2.625 19.990 2.795 ;
        RECT 2.970 2.480 5.065 2.510 ;
        RECT 14.500 2.480 16.845 2.625 ;
        RECT 17.645 2.480 19.990 2.625 ;
        RECT 32.470 2.960 32.640 7.375 ;
        RECT 32.980 2.960 33.270 7.370 ;
        RECT 32.470 2.930 34.565 2.960 ;
        RECT 32.470 2.845 34.720 2.930 ;
        RECT 35.700 2.845 35.870 5.820 ;
        RECT 32.470 2.675 35.870 2.845 ;
        RECT 44.000 2.960 44.170 7.560 ;
        RECT 44.510 2.960 44.800 7.790 ;
        RECT 48.690 2.960 48.980 7.790 ;
        RECT 49.320 2.960 49.490 7.620 ;
        RECT 44.000 2.795 46.345 2.960 ;
        RECT 47.145 2.795 49.490 2.960 ;
        RECT 32.470 2.510 34.720 2.675 ;
        RECT 44.000 2.625 49.490 2.795 ;
        RECT 32.470 2.480 34.565 2.510 ;
        RECT 44.000 2.480 46.345 2.625 ;
        RECT 47.145 2.480 49.490 2.625 ;
        RECT 61.970 2.960 62.140 7.375 ;
        RECT 62.480 2.960 62.770 7.370 ;
        RECT 61.970 2.930 64.065 2.960 ;
        RECT 61.970 2.845 64.220 2.930 ;
        RECT 65.200 2.845 65.370 5.820 ;
        RECT 61.970 2.675 65.370 2.845 ;
        RECT 73.500 2.960 73.670 7.560 ;
        RECT 74.010 2.960 74.300 7.790 ;
        RECT 78.190 2.960 78.480 7.790 ;
        RECT 78.820 2.960 78.990 7.620 ;
        RECT 73.500 2.795 75.845 2.960 ;
        RECT 76.645 2.795 78.990 2.960 ;
        RECT 61.970 2.510 64.220 2.675 ;
        RECT 73.500 2.625 78.990 2.795 ;
        RECT 61.970 2.480 64.065 2.510 ;
        RECT 73.500 2.480 75.845 2.625 ;
        RECT 76.645 2.480 78.990 2.625 ;
        RECT 91.470 2.960 91.640 7.375 ;
        RECT 91.980 2.960 92.270 7.370 ;
        RECT 91.470 2.930 93.565 2.960 ;
        RECT 91.470 2.845 93.720 2.930 ;
        RECT 94.700 2.845 94.870 5.820 ;
        RECT 91.470 2.675 94.870 2.845 ;
        RECT 103.000 2.960 103.170 7.560 ;
        RECT 103.510 2.960 103.800 7.790 ;
        RECT 107.690 2.960 107.980 7.790 ;
        RECT 108.320 2.960 108.490 7.620 ;
        RECT 103.000 2.795 105.345 2.960 ;
        RECT 106.145 2.795 108.490 2.960 ;
        RECT 91.470 2.510 93.720 2.675 ;
        RECT 103.000 2.625 108.490 2.795 ;
        RECT 91.470 2.480 93.565 2.510 ;
        RECT 103.000 2.480 105.345 2.625 ;
        RECT 106.145 2.480 108.490 2.625 ;
        RECT 120.970 2.960 121.140 7.375 ;
        RECT 121.480 2.960 121.770 7.370 ;
        RECT 120.970 2.930 123.065 2.960 ;
        RECT 120.970 2.845 123.220 2.930 ;
        RECT 124.200 2.845 124.370 5.820 ;
        RECT 120.970 2.675 124.370 2.845 ;
        RECT 132.500 2.960 132.670 7.560 ;
        RECT 133.010 2.960 133.300 7.790 ;
        RECT 137.190 2.960 137.480 7.790 ;
        RECT 137.820 2.960 137.990 7.620 ;
        RECT 132.500 2.795 134.845 2.960 ;
        RECT 135.645 2.795 137.990 2.960 ;
        RECT 120.970 2.510 123.220 2.675 ;
        RECT 132.500 2.625 137.990 2.795 ;
        RECT 120.970 2.480 123.065 2.510 ;
        RECT 132.500 2.480 134.845 2.625 ;
        RECT 135.645 2.480 137.990 2.625 ;
        RECT 150.470 2.960 150.640 7.375 ;
        RECT 150.980 2.960 151.270 7.370 ;
        RECT 150.470 2.930 152.565 2.960 ;
        RECT 150.470 2.845 152.720 2.930 ;
        RECT 153.700 2.845 153.870 5.820 ;
        RECT 150.470 2.675 153.870 2.845 ;
        RECT 162.000 2.960 162.170 7.560 ;
        RECT 162.510 2.960 162.800 7.790 ;
        RECT 166.690 2.960 166.980 7.790 ;
        RECT 167.320 2.960 167.490 7.620 ;
        RECT 162.000 2.795 164.345 2.960 ;
        RECT 165.145 2.795 167.490 2.960 ;
        RECT 150.470 2.510 152.720 2.675 ;
        RECT 162.000 2.625 167.490 2.795 ;
        RECT 150.470 2.480 152.565 2.510 ;
        RECT 162.000 2.480 164.345 2.625 ;
        RECT 165.145 2.480 167.490 2.625 ;
      LAYER mcon ;
        RECT 3.580 2.510 4.000 2.930 ;
        RECT 4.190 2.510 4.610 2.930 ;
        RECT 4.800 2.510 5.220 2.930 ;
        RECT 14.500 2.510 15.015 2.930 ;
        RECT 15.205 2.510 15.625 2.930 ;
        RECT 15.815 2.510 16.235 2.930 ;
        RECT 16.425 2.510 16.845 2.930 ;
        RECT 17.645 2.510 18.065 2.930 ;
        RECT 18.255 2.510 18.675 2.930 ;
        RECT 18.865 2.510 19.285 2.930 ;
        RECT 19.475 2.510 19.990 2.930 ;
        RECT 33.080 2.510 33.500 2.930 ;
        RECT 33.690 2.510 34.110 2.930 ;
        RECT 34.300 2.510 34.720 2.930 ;
        RECT 44.000 2.510 44.515 2.930 ;
        RECT 44.705 2.510 45.125 2.930 ;
        RECT 45.315 2.510 45.735 2.930 ;
        RECT 45.925 2.510 46.345 2.930 ;
        RECT 47.145 2.510 47.565 2.930 ;
        RECT 47.755 2.510 48.175 2.930 ;
        RECT 48.365 2.510 48.785 2.930 ;
        RECT 48.975 2.510 49.490 2.930 ;
        RECT 62.580 2.510 63.000 2.930 ;
        RECT 63.190 2.510 63.610 2.930 ;
        RECT 63.800 2.510 64.220 2.930 ;
        RECT 73.500 2.510 74.015 2.930 ;
        RECT 74.205 2.510 74.625 2.930 ;
        RECT 74.815 2.510 75.235 2.930 ;
        RECT 75.425 2.510 75.845 2.930 ;
        RECT 76.645 2.510 77.065 2.930 ;
        RECT 77.255 2.510 77.675 2.930 ;
        RECT 77.865 2.510 78.285 2.930 ;
        RECT 78.475 2.510 78.990 2.930 ;
        RECT 92.080 2.510 92.500 2.930 ;
        RECT 92.690 2.510 93.110 2.930 ;
        RECT 93.300 2.510 93.720 2.930 ;
        RECT 103.000 2.510 103.515 2.930 ;
        RECT 103.705 2.510 104.125 2.930 ;
        RECT 104.315 2.510 104.735 2.930 ;
        RECT 104.925 2.510 105.345 2.930 ;
        RECT 106.145 2.510 106.565 2.930 ;
        RECT 106.755 2.510 107.175 2.930 ;
        RECT 107.365 2.510 107.785 2.930 ;
        RECT 107.975 2.510 108.490 2.930 ;
        RECT 121.580 2.510 122.000 2.930 ;
        RECT 122.190 2.510 122.610 2.930 ;
        RECT 122.800 2.510 123.220 2.930 ;
        RECT 132.500 2.510 133.015 2.930 ;
        RECT 133.205 2.510 133.625 2.930 ;
        RECT 133.815 2.510 134.235 2.930 ;
        RECT 134.425 2.510 134.845 2.930 ;
        RECT 135.645 2.510 136.065 2.930 ;
        RECT 136.255 2.510 136.675 2.930 ;
        RECT 136.865 2.510 137.285 2.930 ;
        RECT 137.475 2.510 137.990 2.930 ;
        RECT 151.080 2.510 151.500 2.930 ;
        RECT 151.690 2.510 152.110 2.930 ;
        RECT 152.300 2.510 152.720 2.930 ;
        RECT 162.000 2.510 162.515 2.930 ;
        RECT 162.705 2.510 163.125 2.930 ;
        RECT 163.315 2.510 163.735 2.930 ;
        RECT 163.925 2.510 164.345 2.930 ;
        RECT 165.145 2.510 165.565 2.930 ;
        RECT 165.755 2.510 166.175 2.930 ;
        RECT 166.365 2.510 166.785 2.930 ;
        RECT 166.975 2.510 167.490 2.930 ;
      LAYER met1 ;
        RECT 0.000 2.480 179.440 2.960 ;
    END
    PORT
      LAYER nwell ;
        RECT 9.265 8.520 13.025 13.830 ;
        RECT 25.150 7.960 31.000 13.835 ;
        RECT 38.765 8.520 42.525 13.830 ;
        RECT 54.650 7.960 60.500 13.835 ;
        RECT 68.265 8.520 72.025 13.830 ;
        RECT 84.150 7.960 90.000 13.835 ;
        RECT 97.765 8.520 101.525 13.830 ;
        RECT 113.650 7.960 119.500 13.835 ;
        RECT 127.265 8.520 131.025 13.830 ;
        RECT 143.150 7.960 149.000 13.835 ;
        RECT 156.765 8.520 160.525 13.830 ;
        RECT 172.650 7.960 178.500 13.835 ;
      LAYER li1 ;
        RECT 10.750 13.810 12.845 13.840 ;
        RECT 25.330 13.810 27.675 13.840 ;
        RECT 10.595 13.650 12.845 13.810 ;
        RECT 9.445 13.480 12.845 13.650 ;
        RECT 9.445 9.445 9.615 13.480 ;
        RECT 10.595 13.390 12.845 13.480 ;
        RECT 25.150 13.655 27.675 13.810 ;
        RECT 28.475 13.655 30.820 13.840 ;
        RECT 40.250 13.810 42.345 13.840 ;
        RECT 54.830 13.810 57.175 13.840 ;
        RECT 25.150 13.485 30.820 13.655 ;
        RECT 40.095 13.650 42.345 13.810 ;
        RECT 25.150 13.390 27.675 13.485 ;
        RECT 10.750 13.360 12.845 13.390 ;
        RECT 12.045 9.290 12.335 13.360 ;
        RECT 12.675 9.435 12.845 13.360 ;
        RECT 25.330 13.360 27.675 13.390 ;
        RECT 28.475 13.360 30.820 13.485 ;
        RECT 25.330 8.505 25.500 13.360 ;
        RECT 25.840 8.510 26.130 13.360 ;
        RECT 30.020 8.510 30.310 13.360 ;
        RECT 30.650 8.505 30.820 13.360 ;
        RECT 38.945 13.480 42.345 13.650 ;
        RECT 38.945 9.445 39.115 13.480 ;
        RECT 40.095 13.390 42.345 13.480 ;
        RECT 54.650 13.655 57.175 13.810 ;
        RECT 57.975 13.655 60.320 13.840 ;
        RECT 69.750 13.810 71.845 13.840 ;
        RECT 84.330 13.810 86.675 13.840 ;
        RECT 54.650 13.485 60.320 13.655 ;
        RECT 69.595 13.650 71.845 13.810 ;
        RECT 54.650 13.390 57.175 13.485 ;
        RECT 40.250 13.360 42.345 13.390 ;
        RECT 41.545 9.290 41.835 13.360 ;
        RECT 42.175 9.435 42.345 13.360 ;
        RECT 54.830 13.360 57.175 13.390 ;
        RECT 57.975 13.360 60.320 13.485 ;
        RECT 54.830 8.505 55.000 13.360 ;
        RECT 55.340 8.510 55.630 13.360 ;
        RECT 59.520 8.510 59.810 13.360 ;
        RECT 60.150 8.505 60.320 13.360 ;
        RECT 68.445 13.480 71.845 13.650 ;
        RECT 68.445 9.445 68.615 13.480 ;
        RECT 69.595 13.390 71.845 13.480 ;
        RECT 84.150 13.655 86.675 13.810 ;
        RECT 87.475 13.655 89.820 13.840 ;
        RECT 99.250 13.810 101.345 13.840 ;
        RECT 113.830 13.810 116.175 13.840 ;
        RECT 84.150 13.485 89.820 13.655 ;
        RECT 99.095 13.650 101.345 13.810 ;
        RECT 84.150 13.390 86.675 13.485 ;
        RECT 69.750 13.360 71.845 13.390 ;
        RECT 71.045 9.290 71.335 13.360 ;
        RECT 71.675 9.435 71.845 13.360 ;
        RECT 84.330 13.360 86.675 13.390 ;
        RECT 87.475 13.360 89.820 13.485 ;
        RECT 84.330 8.505 84.500 13.360 ;
        RECT 84.840 8.510 85.130 13.360 ;
        RECT 89.020 8.510 89.310 13.360 ;
        RECT 89.650 8.505 89.820 13.360 ;
        RECT 97.945 13.480 101.345 13.650 ;
        RECT 97.945 9.445 98.115 13.480 ;
        RECT 99.095 13.390 101.345 13.480 ;
        RECT 113.650 13.655 116.175 13.810 ;
        RECT 116.975 13.655 119.320 13.840 ;
        RECT 128.750 13.810 130.845 13.840 ;
        RECT 143.330 13.810 145.675 13.840 ;
        RECT 113.650 13.485 119.320 13.655 ;
        RECT 128.595 13.650 130.845 13.810 ;
        RECT 113.650 13.390 116.175 13.485 ;
        RECT 99.250 13.360 101.345 13.390 ;
        RECT 100.545 9.290 100.835 13.360 ;
        RECT 101.175 9.435 101.345 13.360 ;
        RECT 113.830 13.360 116.175 13.390 ;
        RECT 116.975 13.360 119.320 13.485 ;
        RECT 113.830 8.505 114.000 13.360 ;
        RECT 114.340 8.510 114.630 13.360 ;
        RECT 118.520 8.510 118.810 13.360 ;
        RECT 119.150 8.505 119.320 13.360 ;
        RECT 127.445 13.480 130.845 13.650 ;
        RECT 127.445 9.445 127.615 13.480 ;
        RECT 128.595 13.390 130.845 13.480 ;
        RECT 143.150 13.655 145.675 13.810 ;
        RECT 146.475 13.655 148.820 13.840 ;
        RECT 158.250 13.810 160.345 13.840 ;
        RECT 172.830 13.810 175.175 13.840 ;
        RECT 143.150 13.485 148.820 13.655 ;
        RECT 158.095 13.650 160.345 13.810 ;
        RECT 143.150 13.390 145.675 13.485 ;
        RECT 128.750 13.360 130.845 13.390 ;
        RECT 130.045 9.290 130.335 13.360 ;
        RECT 130.675 9.435 130.845 13.360 ;
        RECT 143.330 13.360 145.675 13.390 ;
        RECT 146.475 13.360 148.820 13.485 ;
        RECT 143.330 8.505 143.500 13.360 ;
        RECT 143.840 8.510 144.130 13.360 ;
        RECT 148.020 8.510 148.310 13.360 ;
        RECT 148.650 8.505 148.820 13.360 ;
        RECT 156.945 13.480 160.345 13.650 ;
        RECT 156.945 9.445 157.115 13.480 ;
        RECT 158.095 13.390 160.345 13.480 ;
        RECT 172.650 13.655 175.175 13.810 ;
        RECT 175.975 13.655 178.320 13.840 ;
        RECT 172.650 13.485 178.320 13.655 ;
        RECT 172.650 13.390 175.175 13.485 ;
        RECT 158.250 13.360 160.345 13.390 ;
        RECT 159.545 9.290 159.835 13.360 ;
        RECT 160.175 9.435 160.345 13.360 ;
        RECT 172.830 13.360 175.175 13.390 ;
        RECT 175.975 13.360 178.320 13.485 ;
        RECT 172.830 8.505 173.000 13.360 ;
        RECT 173.340 8.510 173.630 13.360 ;
        RECT 177.520 8.510 177.810 13.360 ;
        RECT 178.150 8.505 178.320 13.360 ;
      LAYER mcon ;
        RECT 11.205 13.390 11.625 13.810 ;
        RECT 11.815 13.390 12.235 13.810 ;
        RECT 12.425 13.390 12.845 13.810 ;
        RECT 25.855 13.390 26.275 13.810 ;
        RECT 26.465 13.390 26.885 13.810 ;
        RECT 27.075 13.390 27.495 13.810 ;
        RECT 28.475 13.390 28.895 13.810 ;
        RECT 29.085 13.390 29.505 13.810 ;
        RECT 29.695 13.390 30.115 13.810 ;
        RECT 30.305 13.390 30.820 13.810 ;
        RECT 40.705 13.390 41.125 13.810 ;
        RECT 41.315 13.390 41.735 13.810 ;
        RECT 41.925 13.390 42.345 13.810 ;
        RECT 55.355 13.390 55.775 13.810 ;
        RECT 55.965 13.390 56.385 13.810 ;
        RECT 56.575 13.390 56.995 13.810 ;
        RECT 57.975 13.390 58.395 13.810 ;
        RECT 58.585 13.390 59.005 13.810 ;
        RECT 59.195 13.390 59.615 13.810 ;
        RECT 59.805 13.390 60.320 13.810 ;
        RECT 70.205 13.390 70.625 13.810 ;
        RECT 70.815 13.390 71.235 13.810 ;
        RECT 71.425 13.390 71.845 13.810 ;
        RECT 84.855 13.390 85.275 13.810 ;
        RECT 85.465 13.390 85.885 13.810 ;
        RECT 86.075 13.390 86.495 13.810 ;
        RECT 87.475 13.390 87.895 13.810 ;
        RECT 88.085 13.390 88.505 13.810 ;
        RECT 88.695 13.390 89.115 13.810 ;
        RECT 89.305 13.390 89.820 13.810 ;
        RECT 99.705 13.390 100.125 13.810 ;
        RECT 100.315 13.390 100.735 13.810 ;
        RECT 100.925 13.390 101.345 13.810 ;
        RECT 114.355 13.390 114.775 13.810 ;
        RECT 114.965 13.390 115.385 13.810 ;
        RECT 115.575 13.390 115.995 13.810 ;
        RECT 116.975 13.390 117.395 13.810 ;
        RECT 117.585 13.390 118.005 13.810 ;
        RECT 118.195 13.390 118.615 13.810 ;
        RECT 118.805 13.390 119.320 13.810 ;
        RECT 129.205 13.390 129.625 13.810 ;
        RECT 129.815 13.390 130.235 13.810 ;
        RECT 130.425 13.390 130.845 13.810 ;
        RECT 143.855 13.390 144.275 13.810 ;
        RECT 144.465 13.390 144.885 13.810 ;
        RECT 145.075 13.390 145.495 13.810 ;
        RECT 146.475 13.390 146.895 13.810 ;
        RECT 147.085 13.390 147.505 13.810 ;
        RECT 147.695 13.390 148.115 13.810 ;
        RECT 148.305 13.390 148.820 13.810 ;
        RECT 158.705 13.390 159.125 13.810 ;
        RECT 159.315 13.390 159.735 13.810 ;
        RECT 159.925 13.390 160.345 13.810 ;
        RECT 173.355 13.390 173.775 13.810 ;
        RECT 173.965 13.390 174.385 13.810 ;
        RECT 174.575 13.390 174.995 13.810 ;
        RECT 175.975 13.390 176.395 13.810 ;
        RECT 176.585 13.390 177.005 13.810 ;
        RECT 177.195 13.390 177.615 13.810 ;
        RECT 177.805 13.390 178.320 13.810 ;
      LAYER met1 ;
        RECT 0.000 13.360 179.440 13.840 ;
    END
    PORT
      LAYER nwell ;
        RECT 18.390 24.245 24.240 30.120 ;
        RECT 36.365 24.250 40.125 29.560 ;
        RECT 47.890 24.245 53.740 30.120 ;
        RECT 65.865 24.250 69.625 29.560 ;
        RECT 77.390 24.245 83.240 30.120 ;
        RECT 95.365 24.250 99.125 29.560 ;
        RECT 106.890 24.245 112.740 30.120 ;
        RECT 124.865 24.250 128.625 29.560 ;
        RECT 136.390 24.245 142.240 30.120 ;
        RECT 154.365 24.250 158.125 29.560 ;
      LAYER li1 ;
        RECT 18.570 24.720 18.740 29.575 ;
        RECT 19.080 24.720 19.370 29.570 ;
        RECT 23.260 24.720 23.550 29.570 ;
        RECT 23.890 24.720 24.060 29.575 ;
        RECT 18.570 24.595 20.915 24.720 ;
        RECT 21.715 24.690 24.060 24.720 ;
        RECT 36.545 24.720 36.715 28.645 ;
        RECT 37.055 24.720 37.345 28.790 ;
        RECT 36.545 24.690 38.640 24.720 ;
        RECT 21.715 24.595 24.240 24.690 ;
        RECT 18.570 24.425 24.240 24.595 ;
        RECT 18.570 24.240 20.915 24.425 ;
        RECT 21.715 24.270 24.240 24.425 ;
        RECT 36.545 24.600 38.795 24.690 ;
        RECT 39.775 24.600 39.945 28.635 ;
        RECT 36.545 24.430 39.945 24.600 ;
        RECT 48.070 24.720 48.240 29.575 ;
        RECT 48.580 24.720 48.870 29.570 ;
        RECT 52.760 24.720 53.050 29.570 ;
        RECT 53.390 24.720 53.560 29.575 ;
        RECT 48.070 24.595 50.415 24.720 ;
        RECT 51.215 24.690 53.560 24.720 ;
        RECT 66.045 24.720 66.215 28.645 ;
        RECT 66.555 24.720 66.845 28.790 ;
        RECT 66.045 24.690 68.140 24.720 ;
        RECT 51.215 24.595 53.740 24.690 ;
        RECT 36.545 24.270 38.795 24.430 ;
        RECT 48.070 24.425 53.740 24.595 ;
        RECT 21.715 24.240 24.060 24.270 ;
        RECT 36.545 24.240 38.640 24.270 ;
        RECT 48.070 24.240 50.415 24.425 ;
        RECT 51.215 24.270 53.740 24.425 ;
        RECT 66.045 24.600 68.295 24.690 ;
        RECT 69.275 24.600 69.445 28.635 ;
        RECT 66.045 24.430 69.445 24.600 ;
        RECT 77.570 24.720 77.740 29.575 ;
        RECT 78.080 24.720 78.370 29.570 ;
        RECT 82.260 24.720 82.550 29.570 ;
        RECT 82.890 24.720 83.060 29.575 ;
        RECT 77.570 24.595 79.915 24.720 ;
        RECT 80.715 24.690 83.060 24.720 ;
        RECT 95.545 24.720 95.715 28.645 ;
        RECT 96.055 24.720 96.345 28.790 ;
        RECT 95.545 24.690 97.640 24.720 ;
        RECT 80.715 24.595 83.240 24.690 ;
        RECT 66.045 24.270 68.295 24.430 ;
        RECT 77.570 24.425 83.240 24.595 ;
        RECT 51.215 24.240 53.560 24.270 ;
        RECT 66.045 24.240 68.140 24.270 ;
        RECT 77.570 24.240 79.915 24.425 ;
        RECT 80.715 24.270 83.240 24.425 ;
        RECT 95.545 24.600 97.795 24.690 ;
        RECT 98.775 24.600 98.945 28.635 ;
        RECT 95.545 24.430 98.945 24.600 ;
        RECT 107.070 24.720 107.240 29.575 ;
        RECT 107.580 24.720 107.870 29.570 ;
        RECT 111.760 24.720 112.050 29.570 ;
        RECT 112.390 24.720 112.560 29.575 ;
        RECT 107.070 24.595 109.415 24.720 ;
        RECT 110.215 24.690 112.560 24.720 ;
        RECT 125.045 24.720 125.215 28.645 ;
        RECT 125.555 24.720 125.845 28.790 ;
        RECT 125.045 24.690 127.140 24.720 ;
        RECT 110.215 24.595 112.740 24.690 ;
        RECT 95.545 24.270 97.795 24.430 ;
        RECT 107.070 24.425 112.740 24.595 ;
        RECT 80.715 24.240 83.060 24.270 ;
        RECT 95.545 24.240 97.640 24.270 ;
        RECT 107.070 24.240 109.415 24.425 ;
        RECT 110.215 24.270 112.740 24.425 ;
        RECT 125.045 24.600 127.295 24.690 ;
        RECT 128.275 24.600 128.445 28.635 ;
        RECT 125.045 24.430 128.445 24.600 ;
        RECT 136.570 24.720 136.740 29.575 ;
        RECT 137.080 24.720 137.370 29.570 ;
        RECT 141.260 24.720 141.550 29.570 ;
        RECT 141.890 24.720 142.060 29.575 ;
        RECT 136.570 24.595 138.915 24.720 ;
        RECT 139.715 24.690 142.060 24.720 ;
        RECT 154.545 24.720 154.715 28.645 ;
        RECT 155.055 24.720 155.345 28.790 ;
        RECT 154.545 24.690 156.640 24.720 ;
        RECT 139.715 24.595 142.240 24.690 ;
        RECT 125.045 24.270 127.295 24.430 ;
        RECT 136.570 24.425 142.240 24.595 ;
        RECT 110.215 24.240 112.560 24.270 ;
        RECT 125.045 24.240 127.140 24.270 ;
        RECT 136.570 24.240 138.915 24.425 ;
        RECT 139.715 24.270 142.240 24.425 ;
        RECT 154.545 24.600 156.795 24.690 ;
        RECT 157.775 24.600 157.945 28.635 ;
        RECT 154.545 24.430 157.945 24.600 ;
        RECT 154.545 24.270 156.795 24.430 ;
        RECT 139.715 24.240 142.060 24.270 ;
        RECT 154.545 24.240 156.640 24.270 ;
      LAYER mcon ;
        RECT 18.570 24.270 19.085 24.690 ;
        RECT 19.275 24.270 19.695 24.690 ;
        RECT 19.885 24.270 20.305 24.690 ;
        RECT 20.495 24.270 20.915 24.690 ;
        RECT 21.895 24.270 22.315 24.690 ;
        RECT 22.505 24.270 22.925 24.690 ;
        RECT 23.115 24.270 23.535 24.690 ;
        RECT 23.725 24.270 24.240 24.690 ;
        RECT 37.155 24.270 37.575 24.690 ;
        RECT 37.765 24.270 38.185 24.690 ;
        RECT 38.375 24.270 38.795 24.690 ;
        RECT 48.070 24.270 48.585 24.690 ;
        RECT 48.775 24.270 49.195 24.690 ;
        RECT 49.385 24.270 49.805 24.690 ;
        RECT 49.995 24.270 50.415 24.690 ;
        RECT 51.395 24.270 51.815 24.690 ;
        RECT 52.005 24.270 52.425 24.690 ;
        RECT 52.615 24.270 53.035 24.690 ;
        RECT 53.225 24.270 53.740 24.690 ;
        RECT 66.655 24.270 67.075 24.690 ;
        RECT 67.265 24.270 67.685 24.690 ;
        RECT 67.875 24.270 68.295 24.690 ;
        RECT 77.570 24.270 78.085 24.690 ;
        RECT 78.275 24.270 78.695 24.690 ;
        RECT 78.885 24.270 79.305 24.690 ;
        RECT 79.495 24.270 79.915 24.690 ;
        RECT 80.895 24.270 81.315 24.690 ;
        RECT 81.505 24.270 81.925 24.690 ;
        RECT 82.115 24.270 82.535 24.690 ;
        RECT 82.725 24.270 83.240 24.690 ;
        RECT 96.155 24.270 96.575 24.690 ;
        RECT 96.765 24.270 97.185 24.690 ;
        RECT 97.375 24.270 97.795 24.690 ;
        RECT 107.070 24.270 107.585 24.690 ;
        RECT 107.775 24.270 108.195 24.690 ;
        RECT 108.385 24.270 108.805 24.690 ;
        RECT 108.995 24.270 109.415 24.690 ;
        RECT 110.395 24.270 110.815 24.690 ;
        RECT 111.005 24.270 111.425 24.690 ;
        RECT 111.615 24.270 112.035 24.690 ;
        RECT 112.225 24.270 112.740 24.690 ;
        RECT 125.655 24.270 126.075 24.690 ;
        RECT 126.265 24.270 126.685 24.690 ;
        RECT 126.875 24.270 127.295 24.690 ;
        RECT 136.570 24.270 137.085 24.690 ;
        RECT 137.275 24.270 137.695 24.690 ;
        RECT 137.885 24.270 138.305 24.690 ;
        RECT 138.495 24.270 138.915 24.690 ;
        RECT 139.895 24.270 140.315 24.690 ;
        RECT 140.505 24.270 140.925 24.690 ;
        RECT 141.115 24.270 141.535 24.690 ;
        RECT 141.725 24.270 142.240 24.690 ;
        RECT 155.155 24.270 155.575 24.690 ;
        RECT 155.765 24.270 156.185 24.690 ;
        RECT 156.375 24.270 156.795 24.690 ;
      LAYER met1 ;
        RECT 0.000 24.240 172.440 24.720 ;
    END
    PORT
      LAYER nwell ;
        RECT 29.220 29.780 35.070 35.635 ;
        RECT 42.840 30.310 46.600 35.585 ;
        RECT 58.720 29.780 64.570 35.635 ;
        RECT 72.340 30.310 76.100 35.585 ;
        RECT 88.220 29.780 94.070 35.635 ;
        RECT 101.840 30.310 105.600 35.585 ;
        RECT 117.720 29.780 123.570 35.635 ;
        RECT 131.340 30.310 135.100 35.585 ;
        RECT 147.220 29.780 153.070 35.635 ;
        RECT 160.840 30.310 164.600 35.585 ;
      LAYER li1 ;
        RECT 29.400 35.455 31.745 35.600 ;
        RECT 32.545 35.455 34.890 35.600 ;
        RECT 44.325 35.570 46.420 35.600 ;
        RECT 29.400 35.285 34.890 35.455 ;
        RECT 44.170 35.405 46.420 35.570 ;
        RECT 29.400 35.120 31.745 35.285 ;
        RECT 32.545 35.120 34.890 35.285 ;
        RECT 29.400 30.460 29.570 35.120 ;
        RECT 29.910 30.290 30.200 35.120 ;
        RECT 34.090 30.290 34.380 35.120 ;
        RECT 34.720 30.520 34.890 35.120 ;
        RECT 43.020 35.235 46.420 35.405 ;
        RECT 43.020 32.260 43.190 35.235 ;
        RECT 44.170 35.150 46.420 35.235 ;
        RECT 44.325 35.120 46.420 35.150 ;
        RECT 45.620 30.710 45.910 35.120 ;
        RECT 46.250 30.705 46.420 35.120 ;
        RECT 58.900 35.455 61.245 35.600 ;
        RECT 62.045 35.455 64.390 35.600 ;
        RECT 73.825 35.570 75.920 35.600 ;
        RECT 58.900 35.285 64.390 35.455 ;
        RECT 73.670 35.405 75.920 35.570 ;
        RECT 58.900 35.120 61.245 35.285 ;
        RECT 62.045 35.120 64.390 35.285 ;
        RECT 58.900 30.460 59.070 35.120 ;
        RECT 59.410 30.290 59.700 35.120 ;
        RECT 63.590 30.290 63.880 35.120 ;
        RECT 64.220 30.520 64.390 35.120 ;
        RECT 72.520 35.235 75.920 35.405 ;
        RECT 72.520 32.260 72.690 35.235 ;
        RECT 73.670 35.150 75.920 35.235 ;
        RECT 73.825 35.120 75.920 35.150 ;
        RECT 75.120 30.710 75.410 35.120 ;
        RECT 75.750 30.705 75.920 35.120 ;
        RECT 88.400 35.455 90.745 35.600 ;
        RECT 91.545 35.455 93.890 35.600 ;
        RECT 103.325 35.570 105.420 35.600 ;
        RECT 88.400 35.285 93.890 35.455 ;
        RECT 103.170 35.405 105.420 35.570 ;
        RECT 88.400 35.120 90.745 35.285 ;
        RECT 91.545 35.120 93.890 35.285 ;
        RECT 88.400 30.460 88.570 35.120 ;
        RECT 88.910 30.290 89.200 35.120 ;
        RECT 93.090 30.290 93.380 35.120 ;
        RECT 93.720 30.520 93.890 35.120 ;
        RECT 102.020 35.235 105.420 35.405 ;
        RECT 102.020 32.260 102.190 35.235 ;
        RECT 103.170 35.150 105.420 35.235 ;
        RECT 103.325 35.120 105.420 35.150 ;
        RECT 104.620 30.710 104.910 35.120 ;
        RECT 105.250 30.705 105.420 35.120 ;
        RECT 117.900 35.455 120.245 35.600 ;
        RECT 121.045 35.455 123.390 35.600 ;
        RECT 132.825 35.570 134.920 35.600 ;
        RECT 117.900 35.285 123.390 35.455 ;
        RECT 132.670 35.405 134.920 35.570 ;
        RECT 117.900 35.120 120.245 35.285 ;
        RECT 121.045 35.120 123.390 35.285 ;
        RECT 117.900 30.460 118.070 35.120 ;
        RECT 118.410 30.290 118.700 35.120 ;
        RECT 122.590 30.290 122.880 35.120 ;
        RECT 123.220 30.520 123.390 35.120 ;
        RECT 131.520 35.235 134.920 35.405 ;
        RECT 131.520 32.260 131.690 35.235 ;
        RECT 132.670 35.150 134.920 35.235 ;
        RECT 132.825 35.120 134.920 35.150 ;
        RECT 134.120 30.710 134.410 35.120 ;
        RECT 134.750 30.705 134.920 35.120 ;
        RECT 147.400 35.455 149.745 35.600 ;
        RECT 150.545 35.455 152.890 35.600 ;
        RECT 162.325 35.570 164.420 35.600 ;
        RECT 147.400 35.285 152.890 35.455 ;
        RECT 162.170 35.405 164.420 35.570 ;
        RECT 147.400 35.120 149.745 35.285 ;
        RECT 150.545 35.120 152.890 35.285 ;
        RECT 147.400 30.460 147.570 35.120 ;
        RECT 147.910 30.290 148.200 35.120 ;
        RECT 152.090 30.290 152.380 35.120 ;
        RECT 152.720 30.520 152.890 35.120 ;
        RECT 161.020 35.235 164.420 35.405 ;
        RECT 161.020 32.260 161.190 35.235 ;
        RECT 162.170 35.150 164.420 35.235 ;
        RECT 162.325 35.120 164.420 35.150 ;
        RECT 163.620 30.710 163.910 35.120 ;
        RECT 164.250 30.705 164.420 35.120 ;
      LAYER mcon ;
        RECT 29.400 35.150 29.915 35.570 ;
        RECT 30.105 35.150 30.525 35.570 ;
        RECT 30.715 35.150 31.135 35.570 ;
        RECT 31.325 35.150 31.745 35.570 ;
        RECT 32.545 35.150 32.965 35.570 ;
        RECT 33.155 35.150 33.575 35.570 ;
        RECT 33.765 35.150 34.185 35.570 ;
        RECT 34.375 35.150 34.890 35.570 ;
        RECT 44.780 35.150 45.200 35.570 ;
        RECT 45.390 35.150 45.810 35.570 ;
        RECT 46.000 35.150 46.420 35.570 ;
        RECT 58.900 35.150 59.415 35.570 ;
        RECT 59.605 35.150 60.025 35.570 ;
        RECT 60.215 35.150 60.635 35.570 ;
        RECT 60.825 35.150 61.245 35.570 ;
        RECT 62.045 35.150 62.465 35.570 ;
        RECT 62.655 35.150 63.075 35.570 ;
        RECT 63.265 35.150 63.685 35.570 ;
        RECT 63.875 35.150 64.390 35.570 ;
        RECT 74.280 35.150 74.700 35.570 ;
        RECT 74.890 35.150 75.310 35.570 ;
        RECT 75.500 35.150 75.920 35.570 ;
        RECT 88.400 35.150 88.915 35.570 ;
        RECT 89.105 35.150 89.525 35.570 ;
        RECT 89.715 35.150 90.135 35.570 ;
        RECT 90.325 35.150 90.745 35.570 ;
        RECT 91.545 35.150 91.965 35.570 ;
        RECT 92.155 35.150 92.575 35.570 ;
        RECT 92.765 35.150 93.185 35.570 ;
        RECT 93.375 35.150 93.890 35.570 ;
        RECT 103.780 35.150 104.200 35.570 ;
        RECT 104.390 35.150 104.810 35.570 ;
        RECT 105.000 35.150 105.420 35.570 ;
        RECT 117.900 35.150 118.415 35.570 ;
        RECT 118.605 35.150 119.025 35.570 ;
        RECT 119.215 35.150 119.635 35.570 ;
        RECT 119.825 35.150 120.245 35.570 ;
        RECT 121.045 35.150 121.465 35.570 ;
        RECT 121.655 35.150 122.075 35.570 ;
        RECT 122.265 35.150 122.685 35.570 ;
        RECT 122.875 35.150 123.390 35.570 ;
        RECT 133.280 35.150 133.700 35.570 ;
        RECT 133.890 35.150 134.310 35.570 ;
        RECT 134.500 35.150 134.920 35.570 ;
        RECT 147.400 35.150 147.915 35.570 ;
        RECT 148.105 35.150 148.525 35.570 ;
        RECT 148.715 35.150 149.135 35.570 ;
        RECT 149.325 35.150 149.745 35.570 ;
        RECT 150.545 35.150 150.965 35.570 ;
        RECT 151.155 35.150 151.575 35.570 ;
        RECT 151.765 35.150 152.185 35.570 ;
        RECT 152.375 35.150 152.890 35.570 ;
        RECT 162.780 35.150 163.200 35.570 ;
        RECT 163.390 35.150 163.810 35.570 ;
        RECT 164.000 35.150 164.420 35.570 ;
      LAYER met1 ;
        RECT 0.000 35.120 172.440 35.600 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER li1 ;
        RECT 172.420 26.200 174.420 26.370 ;
        RECT 172.500 26.170 174.340 26.200 ;
      LAYER met1 ;
        RECT 0.000 26.960 174.400 27.440 ;
        RECT 172.440 26.140 174.400 26.960 ;
    END
  END vssd1
  OBS
      LAYER pwell ;
        RECT 18.390 32.310 28.420 38.370 ;
        RECT 36.365 32.270 42.215 38.370 ;
        RECT 47.890 32.310 57.920 38.370 ;
        RECT 65.865 32.270 71.715 38.370 ;
        RECT 77.390 32.310 87.420 38.370 ;
        RECT 95.365 32.270 101.215 38.370 ;
        RECT 106.890 32.310 116.920 38.370 ;
        RECT 124.865 32.270 130.715 38.370 ;
        RECT 136.390 32.310 146.420 38.370 ;
        RECT 154.365 32.270 160.215 38.370 ;
        RECT 25.040 21.460 35.070 27.860 ;
        RECT 40.745 26.625 46.595 27.565 ;
        RECT 40.745 26.575 46.600 26.625 ;
        RECT 40.750 21.465 46.600 26.575 ;
        RECT 54.540 21.460 64.570 27.860 ;
        RECT 70.245 26.625 76.095 27.565 ;
        RECT 70.245 26.575 76.100 26.625 ;
        RECT 70.250 21.465 76.100 26.575 ;
        RECT 84.040 21.460 94.070 27.860 ;
        RECT 99.745 26.625 105.595 27.565 ;
        RECT 99.745 26.575 105.600 26.625 ;
        RECT 99.750 21.465 105.600 26.575 ;
        RECT 113.540 21.460 123.570 27.860 ;
        RECT 129.245 26.625 135.095 27.565 ;
        RECT 129.245 26.575 135.100 26.625 ;
        RECT 129.250 21.465 135.100 26.575 ;
        RECT 143.040 21.460 153.070 27.860 ;
        RECT 158.745 26.625 164.595 27.565 ;
        RECT 158.745 26.575 164.600 26.625 ;
        RECT 158.750 21.465 164.600 26.575 ;
      LAYER nwell ;
        RECT 171.590 20.280 178.380 27.280 ;
      LAYER pwell ;
        RECT 2.790 11.505 8.640 16.615 ;
        RECT 2.790 11.455 8.645 11.505 ;
        RECT 2.795 10.515 8.645 11.455 ;
        RECT 14.320 10.220 24.350 16.620 ;
        RECT 32.290 11.505 38.140 16.615 ;
        RECT 32.290 11.455 38.145 11.505 ;
        RECT 32.295 10.515 38.145 11.455 ;
        RECT 43.820 10.220 53.850 16.620 ;
        RECT 61.790 11.505 67.640 16.615 ;
        RECT 61.790 11.455 67.645 11.505 ;
        RECT 61.795 10.515 67.645 11.455 ;
        RECT 73.320 10.220 83.350 16.620 ;
        RECT 91.290 11.505 97.140 16.615 ;
        RECT 91.290 11.455 97.145 11.505 ;
        RECT 91.295 10.515 97.145 11.455 ;
        RECT 102.820 10.220 112.850 16.620 ;
        RECT 120.790 11.505 126.640 16.615 ;
        RECT 120.790 11.455 126.645 11.505 ;
        RECT 120.795 10.515 126.645 11.455 ;
        RECT 132.320 10.220 142.350 16.620 ;
        RECT 150.290 11.505 156.140 16.615 ;
        RECT 150.290 11.455 156.145 11.505 ;
        RECT 150.295 10.515 156.145 11.455 ;
        RECT 161.820 10.220 171.850 16.620 ;
        RECT 7.175 -0.290 13.025 5.810 ;
        RECT 20.970 -0.290 31.000 5.770 ;
        RECT 36.675 -0.290 42.525 5.810 ;
        RECT 50.470 -0.290 60.500 5.770 ;
        RECT 66.175 -0.290 72.025 5.810 ;
        RECT 79.970 -0.290 90.000 5.770 ;
        RECT 95.675 -0.290 101.525 5.810 ;
        RECT 109.470 -0.290 119.500 5.770 ;
        RECT 125.175 -0.290 131.025 5.810 ;
        RECT 138.970 -0.290 149.000 5.770 ;
        RECT 154.675 -0.290 160.525 5.810 ;
        RECT 168.470 -0.290 178.500 5.770 ;
      LAYER li1 ;
        RECT 18.570 38.190 20.915 38.320 ;
        RECT 21.980 38.190 24.840 38.320 ;
        RECT 25.895 38.190 28.240 38.320 ;
        RECT 18.570 38.020 28.240 38.190 ;
        RECT 18.570 37.840 20.915 38.020 ;
        RECT 21.980 37.840 24.840 38.020 ;
        RECT 25.895 37.840 28.240 38.020 ;
        RECT 18.570 33.190 18.740 37.840 ;
        RECT 19.080 33.245 19.370 37.840 ;
        RECT 19.140 33.000 19.310 33.245 ;
        RECT 19.290 30.790 20.420 31.790 ;
        RECT 21.170 31.480 21.460 37.540 ;
        RECT 23.260 33.245 23.550 37.840 ;
        RECT 23.320 33.000 23.490 33.245 ;
        RECT 25.350 31.580 25.640 37.540 ;
        RECT 27.440 33.245 27.730 37.840 ;
        RECT 27.500 33.235 27.695 33.245 ;
        RECT 27.500 33.000 27.670 33.235 ;
        RECT 28.070 33.090 28.240 37.840 ;
        RECT 36.545 38.180 38.890 38.320 ;
        RECT 39.690 38.180 42.035 38.320 ;
        RECT 36.545 38.010 42.035 38.180 ;
        RECT 36.545 37.840 38.890 38.010 ;
        RECT 39.690 37.840 42.035 38.010 ;
        RECT 36.545 33.485 36.715 37.840 ;
        RECT 37.055 33.490 37.345 37.840 ;
        RECT 41.235 33.490 41.525 37.840 ;
        RECT 41.865 33.485 42.035 37.840 ;
        RECT 48.070 38.190 50.415 38.320 ;
        RECT 51.480 38.190 54.340 38.320 ;
        RECT 55.395 38.190 57.740 38.320 ;
        RECT 48.070 38.020 57.740 38.190 ;
        RECT 48.070 37.840 50.415 38.020 ;
        RECT 51.480 37.840 54.340 38.020 ;
        RECT 55.395 37.840 57.740 38.020 ;
        RECT 37.290 31.580 38.490 31.890 ;
        RECT 43.525 31.675 43.820 34.750 ;
        RECT 48.070 33.190 48.240 37.840 ;
        RECT 48.580 33.245 48.870 37.840 ;
        RECT 48.640 33.000 48.810 33.245 ;
        RECT 25.350 31.480 26.170 31.580 ;
        RECT 21.170 30.980 26.170 31.480 ;
        RECT 21.170 25.030 21.460 30.980 ;
        RECT 36.790 30.960 38.490 31.580 ;
        RECT 37.290 30.760 38.490 30.960 ;
        RECT 43.295 30.895 44.035 31.675 ;
        RECT 25.220 22.000 25.390 26.740 ;
        RECT 25.790 26.595 25.960 26.830 ;
        RECT 25.765 26.585 25.960 26.595 ;
        RECT 29.970 26.585 30.140 26.810 ;
        RECT 34.150 26.585 34.320 26.810 ;
        RECT 25.730 22.000 26.020 26.585 ;
        RECT 29.910 22.000 30.200 26.585 ;
        RECT 34.090 22.000 34.380 26.585 ;
        RECT 34.720 22.000 34.890 26.640 ;
        RECT 25.220 21.810 27.565 22.000 ;
        RECT 28.620 21.810 31.480 22.000 ;
        RECT 32.545 21.810 34.890 22.000 ;
        RECT 25.220 21.640 34.890 21.810 ;
        RECT 25.220 21.520 27.565 21.640 ;
        RECT 28.620 21.520 31.480 21.640 ;
        RECT 32.545 21.520 34.890 21.640 ;
        RECT 40.930 22.000 41.100 26.350 ;
        RECT 41.440 22.000 41.730 26.345 ;
        RECT 43.525 22.305 43.820 30.895 ;
        RECT 48.790 30.790 49.920 31.790 ;
        RECT 50.670 31.480 50.960 37.540 ;
        RECT 52.760 33.245 53.050 37.840 ;
        RECT 52.820 33.000 52.990 33.245 ;
        RECT 54.850 31.580 55.140 37.540 ;
        RECT 56.940 33.245 57.230 37.840 ;
        RECT 57.000 33.235 57.195 33.245 ;
        RECT 57.000 33.000 57.170 33.235 ;
        RECT 57.570 33.090 57.740 37.840 ;
        RECT 66.045 38.180 68.390 38.320 ;
        RECT 69.190 38.180 71.535 38.320 ;
        RECT 66.045 38.010 71.535 38.180 ;
        RECT 66.045 37.840 68.390 38.010 ;
        RECT 69.190 37.840 71.535 38.010 ;
        RECT 66.045 33.485 66.215 37.840 ;
        RECT 66.555 33.490 66.845 37.840 ;
        RECT 70.735 33.490 71.025 37.840 ;
        RECT 71.365 33.485 71.535 37.840 ;
        RECT 77.570 38.190 79.915 38.320 ;
        RECT 80.980 38.190 83.840 38.320 ;
        RECT 84.895 38.190 87.240 38.320 ;
        RECT 77.570 38.020 87.240 38.190 ;
        RECT 77.570 37.840 79.915 38.020 ;
        RECT 80.980 37.840 83.840 38.020 ;
        RECT 84.895 37.840 87.240 38.020 ;
        RECT 66.790 31.580 67.990 31.890 ;
        RECT 73.025 31.675 73.320 34.750 ;
        RECT 77.570 33.190 77.740 37.840 ;
        RECT 78.080 33.245 78.370 37.840 ;
        RECT 78.140 33.000 78.310 33.245 ;
        RECT 54.850 31.480 55.670 31.580 ;
        RECT 50.670 30.980 55.670 31.480 ;
        RECT 45.620 22.000 45.910 26.345 ;
        RECT 46.250 22.000 46.420 26.350 ;
        RECT 50.670 25.030 50.960 30.980 ;
        RECT 66.290 30.960 67.990 31.580 ;
        RECT 66.790 30.760 67.990 30.960 ;
        RECT 72.795 30.895 73.535 31.675 ;
        RECT 40.930 21.825 43.275 22.000 ;
        RECT 44.075 21.825 46.420 22.000 ;
        RECT 40.930 21.655 46.420 21.825 ;
        RECT 40.930 21.520 43.275 21.655 ;
        RECT 44.075 21.520 46.420 21.655 ;
        RECT 54.720 22.000 54.890 26.740 ;
        RECT 55.290 26.595 55.460 26.830 ;
        RECT 55.265 26.585 55.460 26.595 ;
        RECT 59.470 26.585 59.640 26.810 ;
        RECT 63.650 26.585 63.820 26.810 ;
        RECT 55.230 22.000 55.520 26.585 ;
        RECT 59.410 22.000 59.700 26.585 ;
        RECT 63.590 22.000 63.880 26.585 ;
        RECT 64.220 22.000 64.390 26.640 ;
        RECT 54.720 21.810 57.065 22.000 ;
        RECT 58.120 21.810 60.980 22.000 ;
        RECT 62.045 21.810 64.390 22.000 ;
        RECT 54.720 21.640 64.390 21.810 ;
        RECT 54.720 21.520 57.065 21.640 ;
        RECT 58.120 21.520 60.980 21.640 ;
        RECT 62.045 21.520 64.390 21.640 ;
        RECT 70.430 22.000 70.600 26.350 ;
        RECT 70.940 22.000 71.230 26.345 ;
        RECT 73.025 22.305 73.320 30.895 ;
        RECT 78.290 30.790 79.420 31.790 ;
        RECT 80.170 31.480 80.460 37.540 ;
        RECT 82.260 33.245 82.550 37.840 ;
        RECT 82.320 33.000 82.490 33.245 ;
        RECT 84.350 31.580 84.640 37.540 ;
        RECT 86.440 33.245 86.730 37.840 ;
        RECT 86.500 33.235 86.695 33.245 ;
        RECT 86.500 33.000 86.670 33.235 ;
        RECT 87.070 33.090 87.240 37.840 ;
        RECT 95.545 38.180 97.890 38.320 ;
        RECT 98.690 38.180 101.035 38.320 ;
        RECT 95.545 38.010 101.035 38.180 ;
        RECT 95.545 37.840 97.890 38.010 ;
        RECT 98.690 37.840 101.035 38.010 ;
        RECT 95.545 33.485 95.715 37.840 ;
        RECT 96.055 33.490 96.345 37.840 ;
        RECT 100.235 33.490 100.525 37.840 ;
        RECT 100.865 33.485 101.035 37.840 ;
        RECT 107.070 38.190 109.415 38.320 ;
        RECT 110.480 38.190 113.340 38.320 ;
        RECT 114.395 38.190 116.740 38.320 ;
        RECT 107.070 38.020 116.740 38.190 ;
        RECT 107.070 37.840 109.415 38.020 ;
        RECT 110.480 37.840 113.340 38.020 ;
        RECT 114.395 37.840 116.740 38.020 ;
        RECT 96.290 31.580 97.490 31.890 ;
        RECT 102.525 31.675 102.820 34.750 ;
        RECT 107.070 33.190 107.240 37.840 ;
        RECT 107.580 33.245 107.870 37.840 ;
        RECT 107.640 33.000 107.810 33.245 ;
        RECT 84.350 31.480 85.170 31.580 ;
        RECT 80.170 30.980 85.170 31.480 ;
        RECT 75.120 22.000 75.410 26.345 ;
        RECT 75.750 22.000 75.920 26.350 ;
        RECT 80.170 25.030 80.460 30.980 ;
        RECT 95.790 30.960 97.490 31.580 ;
        RECT 96.290 30.760 97.490 30.960 ;
        RECT 102.295 30.895 103.035 31.675 ;
        RECT 70.430 21.825 72.775 22.000 ;
        RECT 73.575 21.825 75.920 22.000 ;
        RECT 70.430 21.655 75.920 21.825 ;
        RECT 70.430 21.520 72.775 21.655 ;
        RECT 73.575 21.520 75.920 21.655 ;
        RECT 84.220 22.000 84.390 26.740 ;
        RECT 84.790 26.595 84.960 26.830 ;
        RECT 84.765 26.585 84.960 26.595 ;
        RECT 88.970 26.585 89.140 26.810 ;
        RECT 93.150 26.585 93.320 26.810 ;
        RECT 84.730 22.000 85.020 26.585 ;
        RECT 88.910 22.000 89.200 26.585 ;
        RECT 93.090 22.000 93.380 26.585 ;
        RECT 93.720 22.000 93.890 26.640 ;
        RECT 84.220 21.810 86.565 22.000 ;
        RECT 87.620 21.810 90.480 22.000 ;
        RECT 91.545 21.810 93.890 22.000 ;
        RECT 84.220 21.640 93.890 21.810 ;
        RECT 84.220 21.520 86.565 21.640 ;
        RECT 87.620 21.520 90.480 21.640 ;
        RECT 91.545 21.520 93.890 21.640 ;
        RECT 99.930 22.000 100.100 26.350 ;
        RECT 100.440 22.000 100.730 26.345 ;
        RECT 102.525 22.305 102.820 30.895 ;
        RECT 107.790 30.790 108.920 31.790 ;
        RECT 109.670 31.480 109.960 37.540 ;
        RECT 111.760 33.245 112.050 37.840 ;
        RECT 111.820 33.000 111.990 33.245 ;
        RECT 113.850 31.580 114.140 37.540 ;
        RECT 115.940 33.245 116.230 37.840 ;
        RECT 116.000 33.235 116.195 33.245 ;
        RECT 116.000 33.000 116.170 33.235 ;
        RECT 116.570 33.090 116.740 37.840 ;
        RECT 125.045 38.180 127.390 38.320 ;
        RECT 128.190 38.180 130.535 38.320 ;
        RECT 125.045 38.010 130.535 38.180 ;
        RECT 125.045 37.840 127.390 38.010 ;
        RECT 128.190 37.840 130.535 38.010 ;
        RECT 125.045 33.485 125.215 37.840 ;
        RECT 125.555 33.490 125.845 37.840 ;
        RECT 129.735 33.490 130.025 37.840 ;
        RECT 130.365 33.485 130.535 37.840 ;
        RECT 136.570 38.190 138.915 38.320 ;
        RECT 139.980 38.190 142.840 38.320 ;
        RECT 143.895 38.190 146.240 38.320 ;
        RECT 136.570 38.020 146.240 38.190 ;
        RECT 136.570 37.840 138.915 38.020 ;
        RECT 139.980 37.840 142.840 38.020 ;
        RECT 143.895 37.840 146.240 38.020 ;
        RECT 125.790 31.580 126.990 31.890 ;
        RECT 132.025 31.675 132.320 34.750 ;
        RECT 136.570 33.190 136.740 37.840 ;
        RECT 137.080 33.245 137.370 37.840 ;
        RECT 137.140 33.000 137.310 33.245 ;
        RECT 113.850 31.480 114.670 31.580 ;
        RECT 109.670 30.980 114.670 31.480 ;
        RECT 104.620 22.000 104.910 26.345 ;
        RECT 105.250 22.000 105.420 26.350 ;
        RECT 109.670 25.030 109.960 30.980 ;
        RECT 125.290 30.960 126.990 31.580 ;
        RECT 125.790 30.760 126.990 30.960 ;
        RECT 131.795 30.895 132.535 31.675 ;
        RECT 99.930 21.825 102.275 22.000 ;
        RECT 103.075 21.825 105.420 22.000 ;
        RECT 99.930 21.655 105.420 21.825 ;
        RECT 99.930 21.520 102.275 21.655 ;
        RECT 103.075 21.520 105.420 21.655 ;
        RECT 113.720 22.000 113.890 26.740 ;
        RECT 114.290 26.595 114.460 26.830 ;
        RECT 114.265 26.585 114.460 26.595 ;
        RECT 118.470 26.585 118.640 26.810 ;
        RECT 122.650 26.585 122.820 26.810 ;
        RECT 114.230 22.000 114.520 26.585 ;
        RECT 118.410 22.000 118.700 26.585 ;
        RECT 122.590 22.000 122.880 26.585 ;
        RECT 123.220 22.000 123.390 26.640 ;
        RECT 113.720 21.810 116.065 22.000 ;
        RECT 117.120 21.810 119.980 22.000 ;
        RECT 121.045 21.810 123.390 22.000 ;
        RECT 113.720 21.640 123.390 21.810 ;
        RECT 113.720 21.520 116.065 21.640 ;
        RECT 117.120 21.520 119.980 21.640 ;
        RECT 121.045 21.520 123.390 21.640 ;
        RECT 129.430 22.000 129.600 26.350 ;
        RECT 129.940 22.000 130.230 26.345 ;
        RECT 132.025 22.305 132.320 30.895 ;
        RECT 137.290 30.790 138.420 31.790 ;
        RECT 139.170 31.480 139.460 37.540 ;
        RECT 141.260 33.245 141.550 37.840 ;
        RECT 141.320 33.000 141.490 33.245 ;
        RECT 143.350 31.580 143.640 37.540 ;
        RECT 145.440 33.245 145.730 37.840 ;
        RECT 145.500 33.235 145.695 33.245 ;
        RECT 145.500 33.000 145.670 33.235 ;
        RECT 146.070 33.090 146.240 37.840 ;
        RECT 154.545 38.180 156.890 38.320 ;
        RECT 157.690 38.180 160.035 38.320 ;
        RECT 154.545 38.010 160.035 38.180 ;
        RECT 154.545 37.840 156.890 38.010 ;
        RECT 157.690 37.840 160.035 38.010 ;
        RECT 154.545 33.485 154.715 37.840 ;
        RECT 155.055 33.490 155.345 37.840 ;
        RECT 159.235 33.490 159.525 37.840 ;
        RECT 159.865 33.485 160.035 37.840 ;
        RECT 155.290 31.580 156.490 31.890 ;
        RECT 161.525 31.675 161.820 34.750 ;
        RECT 143.350 31.480 144.170 31.580 ;
        RECT 139.170 30.980 144.170 31.480 ;
        RECT 134.120 22.000 134.410 26.345 ;
        RECT 134.750 22.000 134.920 26.350 ;
        RECT 139.170 25.030 139.460 30.980 ;
        RECT 154.790 30.960 156.490 31.580 ;
        RECT 155.290 30.760 156.490 30.960 ;
        RECT 161.295 30.895 162.035 31.675 ;
        RECT 129.430 21.825 131.775 22.000 ;
        RECT 132.575 21.825 134.920 22.000 ;
        RECT 129.430 21.655 134.920 21.825 ;
        RECT 129.430 21.520 131.775 21.655 ;
        RECT 132.575 21.520 134.920 21.655 ;
        RECT 143.220 22.000 143.390 26.740 ;
        RECT 143.790 26.595 143.960 26.830 ;
        RECT 143.765 26.585 143.960 26.595 ;
        RECT 147.970 26.585 148.140 26.810 ;
        RECT 152.150 26.585 152.320 26.810 ;
        RECT 143.730 22.000 144.020 26.585 ;
        RECT 147.910 22.000 148.200 26.585 ;
        RECT 152.090 22.000 152.380 26.585 ;
        RECT 152.720 22.000 152.890 26.640 ;
        RECT 143.220 21.810 145.565 22.000 ;
        RECT 146.620 21.810 149.480 22.000 ;
        RECT 150.545 21.810 152.890 22.000 ;
        RECT 143.220 21.640 152.890 21.810 ;
        RECT 143.220 21.520 145.565 21.640 ;
        RECT 146.620 21.520 149.480 21.640 ;
        RECT 150.545 21.520 152.890 21.640 ;
        RECT 158.930 22.000 159.100 26.350 ;
        RECT 159.440 22.000 159.730 26.345 ;
        RECT 161.525 22.305 161.820 30.895 ;
        RECT 171.770 26.930 175.070 27.100 ;
        RECT 163.620 22.000 163.910 26.345 ;
        RECT 164.250 22.000 164.420 26.350 ;
        RECT 158.930 21.825 161.275 22.000 ;
        RECT 162.075 21.825 164.420 22.000 ;
        RECT 158.930 21.655 164.420 21.825 ;
        RECT 158.930 21.520 161.275 21.655 ;
        RECT 162.075 21.520 164.420 21.655 ;
        RECT 171.770 21.090 171.940 26.930 ;
        RECT 174.900 26.640 175.070 26.930 ;
        RECT 174.900 26.470 178.200 26.640 ;
        RECT 172.500 21.820 174.340 21.850 ;
        RECT 172.420 21.650 174.420 21.820 ;
        RECT 174.900 21.090 175.070 26.470 ;
        RECT 175.630 21.360 177.470 21.390 ;
        RECT 175.550 21.190 177.550 21.360 ;
        RECT 171.770 20.920 175.070 21.090 ;
        RECT 174.900 20.630 175.070 20.920 ;
        RECT 178.030 20.630 178.200 26.470 ;
        RECT 174.900 20.460 178.200 20.630 ;
        RECT 2.970 16.425 5.315 16.560 ;
        RECT 6.115 16.425 8.460 16.560 ;
        RECT 2.970 16.255 8.460 16.425 ;
        RECT 2.970 16.080 5.315 16.255 ;
        RECT 6.115 16.080 8.460 16.255 ;
        RECT 2.970 11.730 3.140 16.080 ;
        RECT 3.480 11.735 3.770 16.080 ;
        RECT 5.570 7.185 5.865 15.775 ;
        RECT 7.660 11.735 7.950 16.080 ;
        RECT 8.290 11.730 8.460 16.080 ;
        RECT 14.500 16.440 16.845 16.560 ;
        RECT 17.910 16.440 20.770 16.560 ;
        RECT 21.825 16.440 24.170 16.560 ;
        RECT 14.500 16.270 24.170 16.440 ;
        RECT 14.500 16.080 16.845 16.270 ;
        RECT 17.910 16.080 20.770 16.270 ;
        RECT 21.825 16.080 24.170 16.270 ;
        RECT 14.500 11.440 14.670 16.080 ;
        RECT 15.010 11.495 15.300 16.080 ;
        RECT 19.190 11.495 19.480 16.080 ;
        RECT 23.370 11.495 23.660 16.080 ;
        RECT 15.070 11.270 15.240 11.495 ;
        RECT 19.250 11.270 19.420 11.495 ;
        RECT 23.430 11.485 23.625 11.495 ;
        RECT 23.430 11.250 23.600 11.485 ;
        RECT 24.000 11.340 24.170 16.080 ;
        RECT 32.470 16.425 34.815 16.560 ;
        RECT 35.615 16.425 37.960 16.560 ;
        RECT 32.470 16.255 37.960 16.425 ;
        RECT 32.470 16.080 34.815 16.255 ;
        RECT 35.615 16.080 37.960 16.255 ;
        RECT 5.355 6.405 6.095 7.185 ;
        RECT 10.900 7.120 12.100 7.320 ;
        RECT 10.900 6.500 12.600 7.120 ;
        RECT 27.930 7.100 28.220 13.050 ;
        RECT 32.470 11.730 32.640 16.080 ;
        RECT 32.980 11.735 33.270 16.080 ;
        RECT 23.220 6.600 28.220 7.100 ;
        RECT 23.220 6.500 24.040 6.600 ;
        RECT 5.570 3.330 5.865 6.405 ;
        RECT 10.900 6.190 12.100 6.500 ;
        RECT 7.355 0.240 7.525 4.595 ;
        RECT 7.865 0.240 8.155 4.590 ;
        RECT 12.045 0.240 12.335 4.590 ;
        RECT 12.675 0.240 12.845 4.595 ;
        RECT 7.355 0.070 9.700 0.240 ;
        RECT 10.500 0.070 12.845 0.240 ;
        RECT 7.355 -0.100 12.845 0.070 ;
        RECT 7.355 -0.240 9.700 -0.100 ;
        RECT 10.500 -0.240 12.845 -0.100 ;
        RECT 21.150 0.240 21.320 4.990 ;
        RECT 21.720 4.845 21.890 5.080 ;
        RECT 21.695 4.835 21.890 4.845 ;
        RECT 21.660 0.240 21.950 4.835 ;
        RECT 23.750 0.540 24.040 6.500 ;
        RECT 25.900 4.835 26.070 5.080 ;
        RECT 25.840 0.240 26.130 4.835 ;
        RECT 27.930 0.540 28.220 6.600 ;
        RECT 28.970 6.290 30.100 7.290 ;
        RECT 35.070 7.185 35.365 15.775 ;
        RECT 37.160 11.735 37.450 16.080 ;
        RECT 37.790 11.730 37.960 16.080 ;
        RECT 44.000 16.440 46.345 16.560 ;
        RECT 47.410 16.440 50.270 16.560 ;
        RECT 51.325 16.440 53.670 16.560 ;
        RECT 44.000 16.270 53.670 16.440 ;
        RECT 44.000 16.080 46.345 16.270 ;
        RECT 47.410 16.080 50.270 16.270 ;
        RECT 51.325 16.080 53.670 16.270 ;
        RECT 44.000 11.440 44.170 16.080 ;
        RECT 44.510 11.495 44.800 16.080 ;
        RECT 48.690 11.495 48.980 16.080 ;
        RECT 52.870 11.495 53.160 16.080 ;
        RECT 44.570 11.270 44.740 11.495 ;
        RECT 48.750 11.270 48.920 11.495 ;
        RECT 52.930 11.485 53.125 11.495 ;
        RECT 52.930 11.250 53.100 11.485 ;
        RECT 53.500 11.340 53.670 16.080 ;
        RECT 61.970 16.425 64.315 16.560 ;
        RECT 65.115 16.425 67.460 16.560 ;
        RECT 61.970 16.255 67.460 16.425 ;
        RECT 61.970 16.080 64.315 16.255 ;
        RECT 65.115 16.080 67.460 16.255 ;
        RECT 34.855 6.405 35.595 7.185 ;
        RECT 40.400 7.120 41.600 7.320 ;
        RECT 40.400 6.500 42.100 7.120 ;
        RECT 57.430 7.100 57.720 13.050 ;
        RECT 61.970 11.730 62.140 16.080 ;
        RECT 62.480 11.735 62.770 16.080 ;
        RECT 52.720 6.600 57.720 7.100 ;
        RECT 52.720 6.500 53.540 6.600 ;
        RECT 30.080 4.835 30.250 5.080 ;
        RECT 30.020 0.240 30.310 4.835 ;
        RECT 30.650 0.240 30.820 4.890 ;
        RECT 35.070 3.330 35.365 6.405 ;
        RECT 40.400 6.190 41.600 6.500 ;
        RECT 21.150 0.060 23.495 0.240 ;
        RECT 24.550 0.060 27.410 0.240 ;
        RECT 28.475 0.060 30.820 0.240 ;
        RECT 21.150 -0.110 30.820 0.060 ;
        RECT 21.150 -0.240 23.495 -0.110 ;
        RECT 24.550 -0.240 27.410 -0.110 ;
        RECT 28.475 -0.240 30.820 -0.110 ;
        RECT 36.855 0.240 37.025 4.595 ;
        RECT 37.365 0.240 37.655 4.590 ;
        RECT 41.545 0.240 41.835 4.590 ;
        RECT 42.175 0.240 42.345 4.595 ;
        RECT 36.855 0.070 39.200 0.240 ;
        RECT 40.000 0.070 42.345 0.240 ;
        RECT 36.855 -0.100 42.345 0.070 ;
        RECT 36.855 -0.240 39.200 -0.100 ;
        RECT 40.000 -0.240 42.345 -0.100 ;
        RECT 50.650 0.240 50.820 4.990 ;
        RECT 51.220 4.845 51.390 5.080 ;
        RECT 51.195 4.835 51.390 4.845 ;
        RECT 51.160 0.240 51.450 4.835 ;
        RECT 53.250 0.540 53.540 6.500 ;
        RECT 55.400 4.835 55.570 5.080 ;
        RECT 55.340 0.240 55.630 4.835 ;
        RECT 57.430 0.540 57.720 6.600 ;
        RECT 58.470 6.290 59.600 7.290 ;
        RECT 64.570 7.185 64.865 15.775 ;
        RECT 66.660 11.735 66.950 16.080 ;
        RECT 67.290 11.730 67.460 16.080 ;
        RECT 73.500 16.440 75.845 16.560 ;
        RECT 76.910 16.440 79.770 16.560 ;
        RECT 80.825 16.440 83.170 16.560 ;
        RECT 73.500 16.270 83.170 16.440 ;
        RECT 73.500 16.080 75.845 16.270 ;
        RECT 76.910 16.080 79.770 16.270 ;
        RECT 80.825 16.080 83.170 16.270 ;
        RECT 73.500 11.440 73.670 16.080 ;
        RECT 74.010 11.495 74.300 16.080 ;
        RECT 78.190 11.495 78.480 16.080 ;
        RECT 82.370 11.495 82.660 16.080 ;
        RECT 74.070 11.270 74.240 11.495 ;
        RECT 78.250 11.270 78.420 11.495 ;
        RECT 82.430 11.485 82.625 11.495 ;
        RECT 82.430 11.250 82.600 11.485 ;
        RECT 83.000 11.340 83.170 16.080 ;
        RECT 91.470 16.425 93.815 16.560 ;
        RECT 94.615 16.425 96.960 16.560 ;
        RECT 91.470 16.255 96.960 16.425 ;
        RECT 91.470 16.080 93.815 16.255 ;
        RECT 94.615 16.080 96.960 16.255 ;
        RECT 64.355 6.405 65.095 7.185 ;
        RECT 69.900 7.120 71.100 7.320 ;
        RECT 69.900 6.500 71.600 7.120 ;
        RECT 86.930 7.100 87.220 13.050 ;
        RECT 91.470 11.730 91.640 16.080 ;
        RECT 91.980 11.735 92.270 16.080 ;
        RECT 82.220 6.600 87.220 7.100 ;
        RECT 82.220 6.500 83.040 6.600 ;
        RECT 59.580 4.835 59.750 5.080 ;
        RECT 59.520 0.240 59.810 4.835 ;
        RECT 60.150 0.240 60.320 4.890 ;
        RECT 64.570 3.330 64.865 6.405 ;
        RECT 69.900 6.190 71.100 6.500 ;
        RECT 50.650 0.060 52.995 0.240 ;
        RECT 54.050 0.060 56.910 0.240 ;
        RECT 57.975 0.060 60.320 0.240 ;
        RECT 50.650 -0.110 60.320 0.060 ;
        RECT 50.650 -0.240 52.995 -0.110 ;
        RECT 54.050 -0.240 56.910 -0.110 ;
        RECT 57.975 -0.240 60.320 -0.110 ;
        RECT 66.355 0.240 66.525 4.595 ;
        RECT 66.865 0.240 67.155 4.590 ;
        RECT 71.045 0.240 71.335 4.590 ;
        RECT 71.675 0.240 71.845 4.595 ;
        RECT 66.355 0.070 68.700 0.240 ;
        RECT 69.500 0.070 71.845 0.240 ;
        RECT 66.355 -0.100 71.845 0.070 ;
        RECT 66.355 -0.240 68.700 -0.100 ;
        RECT 69.500 -0.240 71.845 -0.100 ;
        RECT 80.150 0.240 80.320 4.990 ;
        RECT 80.720 4.845 80.890 5.080 ;
        RECT 80.695 4.835 80.890 4.845 ;
        RECT 80.660 0.240 80.950 4.835 ;
        RECT 82.750 0.540 83.040 6.500 ;
        RECT 84.900 4.835 85.070 5.080 ;
        RECT 84.840 0.240 85.130 4.835 ;
        RECT 86.930 0.540 87.220 6.600 ;
        RECT 87.970 6.290 89.100 7.290 ;
        RECT 94.070 7.185 94.365 15.775 ;
        RECT 96.160 11.735 96.450 16.080 ;
        RECT 96.790 11.730 96.960 16.080 ;
        RECT 103.000 16.440 105.345 16.560 ;
        RECT 106.410 16.440 109.270 16.560 ;
        RECT 110.325 16.440 112.670 16.560 ;
        RECT 103.000 16.270 112.670 16.440 ;
        RECT 103.000 16.080 105.345 16.270 ;
        RECT 106.410 16.080 109.270 16.270 ;
        RECT 110.325 16.080 112.670 16.270 ;
        RECT 103.000 11.440 103.170 16.080 ;
        RECT 103.510 11.495 103.800 16.080 ;
        RECT 107.690 11.495 107.980 16.080 ;
        RECT 111.870 11.495 112.160 16.080 ;
        RECT 103.570 11.270 103.740 11.495 ;
        RECT 107.750 11.270 107.920 11.495 ;
        RECT 111.930 11.485 112.125 11.495 ;
        RECT 111.930 11.250 112.100 11.485 ;
        RECT 112.500 11.340 112.670 16.080 ;
        RECT 120.970 16.425 123.315 16.560 ;
        RECT 124.115 16.425 126.460 16.560 ;
        RECT 120.970 16.255 126.460 16.425 ;
        RECT 120.970 16.080 123.315 16.255 ;
        RECT 124.115 16.080 126.460 16.255 ;
        RECT 93.855 6.405 94.595 7.185 ;
        RECT 99.400 7.120 100.600 7.320 ;
        RECT 99.400 6.500 101.100 7.120 ;
        RECT 116.430 7.100 116.720 13.050 ;
        RECT 120.970 11.730 121.140 16.080 ;
        RECT 121.480 11.735 121.770 16.080 ;
        RECT 111.720 6.600 116.720 7.100 ;
        RECT 111.720 6.500 112.540 6.600 ;
        RECT 89.080 4.835 89.250 5.080 ;
        RECT 89.020 0.240 89.310 4.835 ;
        RECT 89.650 0.240 89.820 4.890 ;
        RECT 94.070 3.330 94.365 6.405 ;
        RECT 99.400 6.190 100.600 6.500 ;
        RECT 80.150 0.060 82.495 0.240 ;
        RECT 83.550 0.060 86.410 0.240 ;
        RECT 87.475 0.060 89.820 0.240 ;
        RECT 80.150 -0.110 89.820 0.060 ;
        RECT 80.150 -0.240 82.495 -0.110 ;
        RECT 83.550 -0.240 86.410 -0.110 ;
        RECT 87.475 -0.240 89.820 -0.110 ;
        RECT 95.855 0.240 96.025 4.595 ;
        RECT 96.365 0.240 96.655 4.590 ;
        RECT 100.545 0.240 100.835 4.590 ;
        RECT 101.175 0.240 101.345 4.595 ;
        RECT 95.855 0.070 98.200 0.240 ;
        RECT 99.000 0.070 101.345 0.240 ;
        RECT 95.855 -0.100 101.345 0.070 ;
        RECT 95.855 -0.240 98.200 -0.100 ;
        RECT 99.000 -0.240 101.345 -0.100 ;
        RECT 109.650 0.240 109.820 4.990 ;
        RECT 110.220 4.845 110.390 5.080 ;
        RECT 110.195 4.835 110.390 4.845 ;
        RECT 110.160 0.240 110.450 4.835 ;
        RECT 112.250 0.540 112.540 6.500 ;
        RECT 114.400 4.835 114.570 5.080 ;
        RECT 114.340 0.240 114.630 4.835 ;
        RECT 116.430 0.540 116.720 6.600 ;
        RECT 117.470 6.290 118.600 7.290 ;
        RECT 123.570 7.185 123.865 15.775 ;
        RECT 125.660 11.735 125.950 16.080 ;
        RECT 126.290 11.730 126.460 16.080 ;
        RECT 132.500 16.440 134.845 16.560 ;
        RECT 135.910 16.440 138.770 16.560 ;
        RECT 139.825 16.440 142.170 16.560 ;
        RECT 132.500 16.270 142.170 16.440 ;
        RECT 132.500 16.080 134.845 16.270 ;
        RECT 135.910 16.080 138.770 16.270 ;
        RECT 139.825 16.080 142.170 16.270 ;
        RECT 132.500 11.440 132.670 16.080 ;
        RECT 133.010 11.495 133.300 16.080 ;
        RECT 137.190 11.495 137.480 16.080 ;
        RECT 141.370 11.495 141.660 16.080 ;
        RECT 133.070 11.270 133.240 11.495 ;
        RECT 137.250 11.270 137.420 11.495 ;
        RECT 141.430 11.485 141.625 11.495 ;
        RECT 141.430 11.250 141.600 11.485 ;
        RECT 142.000 11.340 142.170 16.080 ;
        RECT 150.470 16.425 152.815 16.560 ;
        RECT 153.615 16.425 155.960 16.560 ;
        RECT 150.470 16.255 155.960 16.425 ;
        RECT 150.470 16.080 152.815 16.255 ;
        RECT 153.615 16.080 155.960 16.255 ;
        RECT 123.355 6.405 124.095 7.185 ;
        RECT 128.900 7.120 130.100 7.320 ;
        RECT 128.900 6.500 130.600 7.120 ;
        RECT 145.930 7.100 146.220 13.050 ;
        RECT 150.470 11.730 150.640 16.080 ;
        RECT 150.980 11.735 151.270 16.080 ;
        RECT 141.220 6.600 146.220 7.100 ;
        RECT 141.220 6.500 142.040 6.600 ;
        RECT 118.580 4.835 118.750 5.080 ;
        RECT 118.520 0.240 118.810 4.835 ;
        RECT 119.150 0.240 119.320 4.890 ;
        RECT 123.570 3.330 123.865 6.405 ;
        RECT 128.900 6.190 130.100 6.500 ;
        RECT 109.650 0.060 111.995 0.240 ;
        RECT 113.050 0.060 115.910 0.240 ;
        RECT 116.975 0.060 119.320 0.240 ;
        RECT 109.650 -0.110 119.320 0.060 ;
        RECT 109.650 -0.240 111.995 -0.110 ;
        RECT 113.050 -0.240 115.910 -0.110 ;
        RECT 116.975 -0.240 119.320 -0.110 ;
        RECT 125.355 0.240 125.525 4.595 ;
        RECT 125.865 0.240 126.155 4.590 ;
        RECT 130.045 0.240 130.335 4.590 ;
        RECT 130.675 0.240 130.845 4.595 ;
        RECT 125.355 0.070 127.700 0.240 ;
        RECT 128.500 0.070 130.845 0.240 ;
        RECT 125.355 -0.100 130.845 0.070 ;
        RECT 125.355 -0.240 127.700 -0.100 ;
        RECT 128.500 -0.240 130.845 -0.100 ;
        RECT 139.150 0.240 139.320 4.990 ;
        RECT 139.720 4.845 139.890 5.080 ;
        RECT 139.695 4.835 139.890 4.845 ;
        RECT 139.660 0.240 139.950 4.835 ;
        RECT 141.750 0.540 142.040 6.500 ;
        RECT 143.900 4.835 144.070 5.080 ;
        RECT 143.840 0.240 144.130 4.835 ;
        RECT 145.930 0.540 146.220 6.600 ;
        RECT 146.970 6.290 148.100 7.290 ;
        RECT 153.070 7.185 153.365 15.775 ;
        RECT 155.160 11.735 155.450 16.080 ;
        RECT 155.790 11.730 155.960 16.080 ;
        RECT 162.000 16.440 164.345 16.560 ;
        RECT 165.410 16.440 168.270 16.560 ;
        RECT 169.325 16.440 171.670 16.560 ;
        RECT 162.000 16.270 171.670 16.440 ;
        RECT 162.000 16.080 164.345 16.270 ;
        RECT 165.410 16.080 168.270 16.270 ;
        RECT 169.325 16.080 171.670 16.270 ;
        RECT 162.000 11.440 162.170 16.080 ;
        RECT 162.510 11.495 162.800 16.080 ;
        RECT 166.690 11.495 166.980 16.080 ;
        RECT 170.870 11.495 171.160 16.080 ;
        RECT 162.570 11.270 162.740 11.495 ;
        RECT 166.750 11.270 166.920 11.495 ;
        RECT 170.930 11.485 171.125 11.495 ;
        RECT 170.930 11.250 171.100 11.485 ;
        RECT 171.500 11.340 171.670 16.080 ;
        RECT 152.855 6.405 153.595 7.185 ;
        RECT 158.400 7.120 159.600 7.320 ;
        RECT 158.400 6.500 160.100 7.120 ;
        RECT 175.430 7.100 175.720 13.050 ;
        RECT 170.720 6.600 175.720 7.100 ;
        RECT 170.720 6.500 171.540 6.600 ;
        RECT 148.080 4.835 148.250 5.080 ;
        RECT 148.020 0.240 148.310 4.835 ;
        RECT 148.650 0.240 148.820 4.890 ;
        RECT 153.070 3.330 153.365 6.405 ;
        RECT 158.400 6.190 159.600 6.500 ;
        RECT 139.150 0.060 141.495 0.240 ;
        RECT 142.550 0.060 145.410 0.240 ;
        RECT 146.475 0.060 148.820 0.240 ;
        RECT 139.150 -0.110 148.820 0.060 ;
        RECT 139.150 -0.240 141.495 -0.110 ;
        RECT 142.550 -0.240 145.410 -0.110 ;
        RECT 146.475 -0.240 148.820 -0.110 ;
        RECT 154.855 0.240 155.025 4.595 ;
        RECT 155.365 0.240 155.655 4.590 ;
        RECT 159.545 0.240 159.835 4.590 ;
        RECT 160.175 0.240 160.345 4.595 ;
        RECT 154.855 0.070 157.200 0.240 ;
        RECT 158.000 0.070 160.345 0.240 ;
        RECT 154.855 -0.100 160.345 0.070 ;
        RECT 154.855 -0.240 157.200 -0.100 ;
        RECT 158.000 -0.240 160.345 -0.100 ;
        RECT 168.650 0.240 168.820 4.990 ;
        RECT 169.220 4.845 169.390 5.080 ;
        RECT 169.195 4.835 169.390 4.845 ;
        RECT 169.160 0.240 169.450 4.835 ;
        RECT 171.250 0.540 171.540 6.500 ;
        RECT 173.400 4.835 173.570 5.080 ;
        RECT 173.340 0.240 173.630 4.835 ;
        RECT 175.430 0.540 175.720 6.600 ;
        RECT 176.470 6.290 177.600 7.290 ;
        RECT 177.580 4.835 177.750 5.080 ;
        RECT 177.520 0.240 177.810 4.835 ;
        RECT 178.150 0.240 178.320 4.890 ;
        RECT 168.650 0.060 170.995 0.240 ;
        RECT 172.050 0.060 174.910 0.240 ;
        RECT 175.975 0.060 178.320 0.240 ;
        RECT 168.650 -0.110 178.320 0.060 ;
        RECT 168.650 -0.240 170.995 -0.110 ;
        RECT 172.050 -0.240 174.910 -0.110 ;
        RECT 175.975 -0.240 178.320 -0.110 ;
      LAYER mcon ;
        RECT 18.570 37.870 19.085 38.290 ;
        RECT 19.275 37.870 19.695 38.290 ;
        RECT 19.885 37.870 20.305 38.290 ;
        RECT 20.495 37.870 20.915 38.290 ;
        RECT 21.980 37.870 22.400 38.290 ;
        RECT 22.590 37.870 23.010 38.290 ;
        RECT 23.200 37.870 23.620 38.290 ;
        RECT 23.810 37.870 24.230 38.290 ;
        RECT 24.420 37.870 24.840 38.290 ;
        RECT 25.895 37.870 26.315 38.290 ;
        RECT 26.505 37.870 26.925 38.290 ;
        RECT 27.115 37.870 27.535 38.290 ;
        RECT 27.725 37.870 28.240 38.290 ;
        RECT 19.320 30.820 20.330 31.760 ;
        RECT 36.545 37.870 36.965 38.290 ;
        RECT 37.155 37.870 37.575 38.290 ;
        RECT 37.765 37.870 38.185 38.290 ;
        RECT 38.375 37.870 38.890 38.290 ;
        RECT 39.690 37.870 40.205 38.290 ;
        RECT 40.395 37.870 40.815 38.290 ;
        RECT 41.005 37.870 41.425 38.290 ;
        RECT 41.615 37.870 42.035 38.290 ;
        RECT 48.070 37.870 48.585 38.290 ;
        RECT 48.775 37.870 49.195 38.290 ;
        RECT 49.385 37.870 49.805 38.290 ;
        RECT 49.995 37.870 50.415 38.290 ;
        RECT 51.480 37.870 51.900 38.290 ;
        RECT 52.090 37.870 52.510 38.290 ;
        RECT 52.700 37.870 53.120 38.290 ;
        RECT 53.310 37.870 53.730 38.290 ;
        RECT 53.920 37.870 54.340 38.290 ;
        RECT 55.395 37.870 55.815 38.290 ;
        RECT 56.005 37.870 56.425 38.290 ;
        RECT 56.615 37.870 57.035 38.290 ;
        RECT 57.225 37.870 57.740 38.290 ;
        RECT 25.350 30.980 26.170 31.580 ;
        RECT 36.820 30.990 37.270 31.580 ;
        RECT 37.460 30.990 38.490 31.580 ;
        RECT 43.355 30.925 43.975 31.645 ;
        RECT 25.220 21.550 25.735 21.970 ;
        RECT 25.925 21.550 26.345 21.970 ;
        RECT 26.535 21.550 26.955 21.970 ;
        RECT 27.145 21.550 27.565 21.970 ;
        RECT 28.620 21.550 29.040 21.970 ;
        RECT 29.230 21.550 29.650 21.970 ;
        RECT 29.840 21.550 30.260 21.970 ;
        RECT 30.450 21.550 30.870 21.970 ;
        RECT 31.060 21.550 31.480 21.970 ;
        RECT 32.545 21.550 32.965 21.970 ;
        RECT 33.155 21.550 33.575 21.970 ;
        RECT 33.765 21.550 34.185 21.970 ;
        RECT 34.375 21.550 34.890 21.970 ;
        RECT 48.820 30.820 49.830 31.760 ;
        RECT 66.045 37.870 66.465 38.290 ;
        RECT 66.655 37.870 67.075 38.290 ;
        RECT 67.265 37.870 67.685 38.290 ;
        RECT 67.875 37.870 68.390 38.290 ;
        RECT 69.190 37.870 69.705 38.290 ;
        RECT 69.895 37.870 70.315 38.290 ;
        RECT 70.505 37.870 70.925 38.290 ;
        RECT 71.115 37.870 71.535 38.290 ;
        RECT 77.570 37.870 78.085 38.290 ;
        RECT 78.275 37.870 78.695 38.290 ;
        RECT 78.885 37.870 79.305 38.290 ;
        RECT 79.495 37.870 79.915 38.290 ;
        RECT 80.980 37.870 81.400 38.290 ;
        RECT 81.590 37.870 82.010 38.290 ;
        RECT 82.200 37.870 82.620 38.290 ;
        RECT 82.810 37.870 83.230 38.290 ;
        RECT 83.420 37.870 83.840 38.290 ;
        RECT 84.895 37.870 85.315 38.290 ;
        RECT 85.505 37.870 85.925 38.290 ;
        RECT 86.115 37.870 86.535 38.290 ;
        RECT 86.725 37.870 87.240 38.290 ;
        RECT 54.850 30.980 55.670 31.580 ;
        RECT 66.320 30.990 66.770 31.580 ;
        RECT 66.960 30.990 67.990 31.580 ;
        RECT 72.855 30.925 73.475 31.645 ;
        RECT 40.930 21.550 41.445 21.970 ;
        RECT 41.635 21.550 42.055 21.970 ;
        RECT 42.245 21.550 42.665 21.970 ;
        RECT 42.855 21.550 43.275 21.970 ;
        RECT 44.075 21.550 44.495 21.970 ;
        RECT 44.685 21.550 45.105 21.970 ;
        RECT 45.295 21.550 45.715 21.970 ;
        RECT 45.905 21.550 46.420 21.970 ;
        RECT 54.720 21.550 55.235 21.970 ;
        RECT 55.425 21.550 55.845 21.970 ;
        RECT 56.035 21.550 56.455 21.970 ;
        RECT 56.645 21.550 57.065 21.970 ;
        RECT 58.120 21.550 58.540 21.970 ;
        RECT 58.730 21.550 59.150 21.970 ;
        RECT 59.340 21.550 59.760 21.970 ;
        RECT 59.950 21.550 60.370 21.970 ;
        RECT 60.560 21.550 60.980 21.970 ;
        RECT 62.045 21.550 62.465 21.970 ;
        RECT 62.655 21.550 63.075 21.970 ;
        RECT 63.265 21.550 63.685 21.970 ;
        RECT 63.875 21.550 64.390 21.970 ;
        RECT 78.320 30.820 79.330 31.760 ;
        RECT 95.545 37.870 95.965 38.290 ;
        RECT 96.155 37.870 96.575 38.290 ;
        RECT 96.765 37.870 97.185 38.290 ;
        RECT 97.375 37.870 97.890 38.290 ;
        RECT 98.690 37.870 99.205 38.290 ;
        RECT 99.395 37.870 99.815 38.290 ;
        RECT 100.005 37.870 100.425 38.290 ;
        RECT 100.615 37.870 101.035 38.290 ;
        RECT 107.070 37.870 107.585 38.290 ;
        RECT 107.775 37.870 108.195 38.290 ;
        RECT 108.385 37.870 108.805 38.290 ;
        RECT 108.995 37.870 109.415 38.290 ;
        RECT 110.480 37.870 110.900 38.290 ;
        RECT 111.090 37.870 111.510 38.290 ;
        RECT 111.700 37.870 112.120 38.290 ;
        RECT 112.310 37.870 112.730 38.290 ;
        RECT 112.920 37.870 113.340 38.290 ;
        RECT 114.395 37.870 114.815 38.290 ;
        RECT 115.005 37.870 115.425 38.290 ;
        RECT 115.615 37.870 116.035 38.290 ;
        RECT 116.225 37.870 116.740 38.290 ;
        RECT 84.350 30.980 85.170 31.580 ;
        RECT 95.820 30.990 96.270 31.580 ;
        RECT 96.460 30.990 97.490 31.580 ;
        RECT 102.355 30.925 102.975 31.645 ;
        RECT 70.430 21.550 70.945 21.970 ;
        RECT 71.135 21.550 71.555 21.970 ;
        RECT 71.745 21.550 72.165 21.970 ;
        RECT 72.355 21.550 72.775 21.970 ;
        RECT 73.575 21.550 73.995 21.970 ;
        RECT 74.185 21.550 74.605 21.970 ;
        RECT 74.795 21.550 75.215 21.970 ;
        RECT 75.405 21.550 75.920 21.970 ;
        RECT 84.220 21.550 84.735 21.970 ;
        RECT 84.925 21.550 85.345 21.970 ;
        RECT 85.535 21.550 85.955 21.970 ;
        RECT 86.145 21.550 86.565 21.970 ;
        RECT 87.620 21.550 88.040 21.970 ;
        RECT 88.230 21.550 88.650 21.970 ;
        RECT 88.840 21.550 89.260 21.970 ;
        RECT 89.450 21.550 89.870 21.970 ;
        RECT 90.060 21.550 90.480 21.970 ;
        RECT 91.545 21.550 91.965 21.970 ;
        RECT 92.155 21.550 92.575 21.970 ;
        RECT 92.765 21.550 93.185 21.970 ;
        RECT 93.375 21.550 93.890 21.970 ;
        RECT 107.820 30.820 108.830 31.760 ;
        RECT 125.045 37.870 125.465 38.290 ;
        RECT 125.655 37.870 126.075 38.290 ;
        RECT 126.265 37.870 126.685 38.290 ;
        RECT 126.875 37.870 127.390 38.290 ;
        RECT 128.190 37.870 128.705 38.290 ;
        RECT 128.895 37.870 129.315 38.290 ;
        RECT 129.505 37.870 129.925 38.290 ;
        RECT 130.115 37.870 130.535 38.290 ;
        RECT 136.570 37.870 137.085 38.290 ;
        RECT 137.275 37.870 137.695 38.290 ;
        RECT 137.885 37.870 138.305 38.290 ;
        RECT 138.495 37.870 138.915 38.290 ;
        RECT 139.980 37.870 140.400 38.290 ;
        RECT 140.590 37.870 141.010 38.290 ;
        RECT 141.200 37.870 141.620 38.290 ;
        RECT 141.810 37.870 142.230 38.290 ;
        RECT 142.420 37.870 142.840 38.290 ;
        RECT 143.895 37.870 144.315 38.290 ;
        RECT 144.505 37.870 144.925 38.290 ;
        RECT 145.115 37.870 145.535 38.290 ;
        RECT 145.725 37.870 146.240 38.290 ;
        RECT 113.850 30.980 114.670 31.580 ;
        RECT 125.320 30.990 125.770 31.580 ;
        RECT 125.960 30.990 126.990 31.580 ;
        RECT 131.855 30.925 132.475 31.645 ;
        RECT 99.930 21.550 100.445 21.970 ;
        RECT 100.635 21.550 101.055 21.970 ;
        RECT 101.245 21.550 101.665 21.970 ;
        RECT 101.855 21.550 102.275 21.970 ;
        RECT 103.075 21.550 103.495 21.970 ;
        RECT 103.685 21.550 104.105 21.970 ;
        RECT 104.295 21.550 104.715 21.970 ;
        RECT 104.905 21.550 105.420 21.970 ;
        RECT 113.720 21.550 114.235 21.970 ;
        RECT 114.425 21.550 114.845 21.970 ;
        RECT 115.035 21.550 115.455 21.970 ;
        RECT 115.645 21.550 116.065 21.970 ;
        RECT 117.120 21.550 117.540 21.970 ;
        RECT 117.730 21.550 118.150 21.970 ;
        RECT 118.340 21.550 118.760 21.970 ;
        RECT 118.950 21.550 119.370 21.970 ;
        RECT 119.560 21.550 119.980 21.970 ;
        RECT 121.045 21.550 121.465 21.970 ;
        RECT 121.655 21.550 122.075 21.970 ;
        RECT 122.265 21.550 122.685 21.970 ;
        RECT 122.875 21.550 123.390 21.970 ;
        RECT 137.320 30.820 138.330 31.760 ;
        RECT 154.545 37.870 154.965 38.290 ;
        RECT 155.155 37.870 155.575 38.290 ;
        RECT 155.765 37.870 156.185 38.290 ;
        RECT 156.375 37.870 156.890 38.290 ;
        RECT 157.690 37.870 158.205 38.290 ;
        RECT 158.395 37.870 158.815 38.290 ;
        RECT 159.005 37.870 159.425 38.290 ;
        RECT 159.615 37.870 160.035 38.290 ;
        RECT 143.350 30.980 144.170 31.580 ;
        RECT 154.820 30.990 155.270 31.580 ;
        RECT 155.460 30.990 156.490 31.580 ;
        RECT 161.355 30.925 161.975 31.645 ;
        RECT 129.430 21.550 129.945 21.970 ;
        RECT 130.135 21.550 130.555 21.970 ;
        RECT 130.745 21.550 131.165 21.970 ;
        RECT 131.355 21.550 131.775 21.970 ;
        RECT 132.575 21.550 132.995 21.970 ;
        RECT 133.185 21.550 133.605 21.970 ;
        RECT 133.795 21.550 134.215 21.970 ;
        RECT 134.405 21.550 134.920 21.970 ;
        RECT 143.220 21.550 143.735 21.970 ;
        RECT 143.925 21.550 144.345 21.970 ;
        RECT 144.535 21.550 144.955 21.970 ;
        RECT 145.145 21.550 145.565 21.970 ;
        RECT 146.620 21.550 147.040 21.970 ;
        RECT 147.230 21.550 147.650 21.970 ;
        RECT 147.840 21.550 148.260 21.970 ;
        RECT 148.450 21.550 148.870 21.970 ;
        RECT 149.060 21.550 149.480 21.970 ;
        RECT 150.545 21.550 150.965 21.970 ;
        RECT 151.155 21.550 151.575 21.970 ;
        RECT 151.765 21.550 152.185 21.970 ;
        RECT 152.375 21.550 152.890 21.970 ;
        RECT 158.930 21.550 159.445 21.970 ;
        RECT 159.635 21.550 160.055 21.970 ;
        RECT 160.245 21.550 160.665 21.970 ;
        RECT 160.855 21.550 161.275 21.970 ;
        RECT 162.075 21.550 162.495 21.970 ;
        RECT 162.685 21.550 163.105 21.970 ;
        RECT 163.295 21.550 163.715 21.970 ;
        RECT 163.905 21.550 164.420 21.970 ;
        RECT 172.500 21.650 174.340 21.850 ;
        RECT 175.630 21.190 177.470 21.390 ;
        RECT 2.970 16.110 3.485 16.530 ;
        RECT 3.675 16.110 4.095 16.530 ;
        RECT 4.285 16.110 4.705 16.530 ;
        RECT 4.895 16.110 5.315 16.530 ;
        RECT 6.115 16.110 6.535 16.530 ;
        RECT 6.725 16.110 7.145 16.530 ;
        RECT 7.335 16.110 7.755 16.530 ;
        RECT 7.945 16.110 8.460 16.530 ;
        RECT 14.500 16.110 15.015 16.530 ;
        RECT 15.205 16.110 15.625 16.530 ;
        RECT 15.815 16.110 16.235 16.530 ;
        RECT 16.425 16.110 16.845 16.530 ;
        RECT 17.910 16.110 18.330 16.530 ;
        RECT 18.520 16.110 18.940 16.530 ;
        RECT 19.130 16.110 19.550 16.530 ;
        RECT 19.740 16.110 20.160 16.530 ;
        RECT 20.350 16.110 20.770 16.530 ;
        RECT 21.825 16.110 22.245 16.530 ;
        RECT 22.435 16.110 22.855 16.530 ;
        RECT 23.045 16.110 23.465 16.530 ;
        RECT 23.655 16.110 24.170 16.530 ;
        RECT 32.470 16.110 32.985 16.530 ;
        RECT 33.175 16.110 33.595 16.530 ;
        RECT 33.785 16.110 34.205 16.530 ;
        RECT 34.395 16.110 34.815 16.530 ;
        RECT 35.615 16.110 36.035 16.530 ;
        RECT 36.225 16.110 36.645 16.530 ;
        RECT 36.835 16.110 37.255 16.530 ;
        RECT 37.445 16.110 37.960 16.530 ;
        RECT 5.415 6.435 6.035 7.155 ;
        RECT 10.900 6.500 11.930 7.090 ;
        RECT 12.120 6.500 12.570 7.090 ;
        RECT 7.355 -0.210 7.775 0.210 ;
        RECT 7.965 -0.210 8.385 0.210 ;
        RECT 8.575 -0.210 8.995 0.210 ;
        RECT 9.185 -0.210 9.700 0.210 ;
        RECT 10.500 -0.210 11.015 0.210 ;
        RECT 11.205 -0.210 11.625 0.210 ;
        RECT 11.815 -0.210 12.235 0.210 ;
        RECT 12.425 -0.210 12.845 0.210 ;
        RECT 29.060 6.320 30.070 7.260 ;
        RECT 44.000 16.110 44.515 16.530 ;
        RECT 44.705 16.110 45.125 16.530 ;
        RECT 45.315 16.110 45.735 16.530 ;
        RECT 45.925 16.110 46.345 16.530 ;
        RECT 47.410 16.110 47.830 16.530 ;
        RECT 48.020 16.110 48.440 16.530 ;
        RECT 48.630 16.110 49.050 16.530 ;
        RECT 49.240 16.110 49.660 16.530 ;
        RECT 49.850 16.110 50.270 16.530 ;
        RECT 51.325 16.110 51.745 16.530 ;
        RECT 51.935 16.110 52.355 16.530 ;
        RECT 52.545 16.110 52.965 16.530 ;
        RECT 53.155 16.110 53.670 16.530 ;
        RECT 61.970 16.110 62.485 16.530 ;
        RECT 62.675 16.110 63.095 16.530 ;
        RECT 63.285 16.110 63.705 16.530 ;
        RECT 63.895 16.110 64.315 16.530 ;
        RECT 65.115 16.110 65.535 16.530 ;
        RECT 65.725 16.110 66.145 16.530 ;
        RECT 66.335 16.110 66.755 16.530 ;
        RECT 66.945 16.110 67.460 16.530 ;
        RECT 34.915 6.435 35.535 7.155 ;
        RECT 40.400 6.500 41.430 7.090 ;
        RECT 41.620 6.500 42.070 7.090 ;
        RECT 21.150 -0.210 21.665 0.210 ;
        RECT 21.855 -0.210 22.275 0.210 ;
        RECT 22.465 -0.210 22.885 0.210 ;
        RECT 23.075 -0.210 23.495 0.210 ;
        RECT 24.550 -0.210 24.970 0.210 ;
        RECT 25.160 -0.210 25.580 0.210 ;
        RECT 25.770 -0.210 26.190 0.210 ;
        RECT 26.380 -0.210 26.800 0.210 ;
        RECT 26.990 -0.210 27.410 0.210 ;
        RECT 28.475 -0.210 28.895 0.210 ;
        RECT 29.085 -0.210 29.505 0.210 ;
        RECT 29.695 -0.210 30.115 0.210 ;
        RECT 30.305 -0.210 30.820 0.210 ;
        RECT 36.855 -0.210 37.275 0.210 ;
        RECT 37.465 -0.210 37.885 0.210 ;
        RECT 38.075 -0.210 38.495 0.210 ;
        RECT 38.685 -0.210 39.200 0.210 ;
        RECT 40.000 -0.210 40.515 0.210 ;
        RECT 40.705 -0.210 41.125 0.210 ;
        RECT 41.315 -0.210 41.735 0.210 ;
        RECT 41.925 -0.210 42.345 0.210 ;
        RECT 58.560 6.320 59.570 7.260 ;
        RECT 73.500 16.110 74.015 16.530 ;
        RECT 74.205 16.110 74.625 16.530 ;
        RECT 74.815 16.110 75.235 16.530 ;
        RECT 75.425 16.110 75.845 16.530 ;
        RECT 76.910 16.110 77.330 16.530 ;
        RECT 77.520 16.110 77.940 16.530 ;
        RECT 78.130 16.110 78.550 16.530 ;
        RECT 78.740 16.110 79.160 16.530 ;
        RECT 79.350 16.110 79.770 16.530 ;
        RECT 80.825 16.110 81.245 16.530 ;
        RECT 81.435 16.110 81.855 16.530 ;
        RECT 82.045 16.110 82.465 16.530 ;
        RECT 82.655 16.110 83.170 16.530 ;
        RECT 91.470 16.110 91.985 16.530 ;
        RECT 92.175 16.110 92.595 16.530 ;
        RECT 92.785 16.110 93.205 16.530 ;
        RECT 93.395 16.110 93.815 16.530 ;
        RECT 94.615 16.110 95.035 16.530 ;
        RECT 95.225 16.110 95.645 16.530 ;
        RECT 95.835 16.110 96.255 16.530 ;
        RECT 96.445 16.110 96.960 16.530 ;
        RECT 64.415 6.435 65.035 7.155 ;
        RECT 69.900 6.500 70.930 7.090 ;
        RECT 71.120 6.500 71.570 7.090 ;
        RECT 50.650 -0.210 51.165 0.210 ;
        RECT 51.355 -0.210 51.775 0.210 ;
        RECT 51.965 -0.210 52.385 0.210 ;
        RECT 52.575 -0.210 52.995 0.210 ;
        RECT 54.050 -0.210 54.470 0.210 ;
        RECT 54.660 -0.210 55.080 0.210 ;
        RECT 55.270 -0.210 55.690 0.210 ;
        RECT 55.880 -0.210 56.300 0.210 ;
        RECT 56.490 -0.210 56.910 0.210 ;
        RECT 57.975 -0.210 58.395 0.210 ;
        RECT 58.585 -0.210 59.005 0.210 ;
        RECT 59.195 -0.210 59.615 0.210 ;
        RECT 59.805 -0.210 60.320 0.210 ;
        RECT 66.355 -0.210 66.775 0.210 ;
        RECT 66.965 -0.210 67.385 0.210 ;
        RECT 67.575 -0.210 67.995 0.210 ;
        RECT 68.185 -0.210 68.700 0.210 ;
        RECT 69.500 -0.210 70.015 0.210 ;
        RECT 70.205 -0.210 70.625 0.210 ;
        RECT 70.815 -0.210 71.235 0.210 ;
        RECT 71.425 -0.210 71.845 0.210 ;
        RECT 88.060 6.320 89.070 7.260 ;
        RECT 103.000 16.110 103.515 16.530 ;
        RECT 103.705 16.110 104.125 16.530 ;
        RECT 104.315 16.110 104.735 16.530 ;
        RECT 104.925 16.110 105.345 16.530 ;
        RECT 106.410 16.110 106.830 16.530 ;
        RECT 107.020 16.110 107.440 16.530 ;
        RECT 107.630 16.110 108.050 16.530 ;
        RECT 108.240 16.110 108.660 16.530 ;
        RECT 108.850 16.110 109.270 16.530 ;
        RECT 110.325 16.110 110.745 16.530 ;
        RECT 110.935 16.110 111.355 16.530 ;
        RECT 111.545 16.110 111.965 16.530 ;
        RECT 112.155 16.110 112.670 16.530 ;
        RECT 120.970 16.110 121.485 16.530 ;
        RECT 121.675 16.110 122.095 16.530 ;
        RECT 122.285 16.110 122.705 16.530 ;
        RECT 122.895 16.110 123.315 16.530 ;
        RECT 124.115 16.110 124.535 16.530 ;
        RECT 124.725 16.110 125.145 16.530 ;
        RECT 125.335 16.110 125.755 16.530 ;
        RECT 125.945 16.110 126.460 16.530 ;
        RECT 93.915 6.435 94.535 7.155 ;
        RECT 99.400 6.500 100.430 7.090 ;
        RECT 100.620 6.500 101.070 7.090 ;
        RECT 80.150 -0.210 80.665 0.210 ;
        RECT 80.855 -0.210 81.275 0.210 ;
        RECT 81.465 -0.210 81.885 0.210 ;
        RECT 82.075 -0.210 82.495 0.210 ;
        RECT 83.550 -0.210 83.970 0.210 ;
        RECT 84.160 -0.210 84.580 0.210 ;
        RECT 84.770 -0.210 85.190 0.210 ;
        RECT 85.380 -0.210 85.800 0.210 ;
        RECT 85.990 -0.210 86.410 0.210 ;
        RECT 87.475 -0.210 87.895 0.210 ;
        RECT 88.085 -0.210 88.505 0.210 ;
        RECT 88.695 -0.210 89.115 0.210 ;
        RECT 89.305 -0.210 89.820 0.210 ;
        RECT 95.855 -0.210 96.275 0.210 ;
        RECT 96.465 -0.210 96.885 0.210 ;
        RECT 97.075 -0.210 97.495 0.210 ;
        RECT 97.685 -0.210 98.200 0.210 ;
        RECT 99.000 -0.210 99.515 0.210 ;
        RECT 99.705 -0.210 100.125 0.210 ;
        RECT 100.315 -0.210 100.735 0.210 ;
        RECT 100.925 -0.210 101.345 0.210 ;
        RECT 117.560 6.320 118.570 7.260 ;
        RECT 132.500 16.110 133.015 16.530 ;
        RECT 133.205 16.110 133.625 16.530 ;
        RECT 133.815 16.110 134.235 16.530 ;
        RECT 134.425 16.110 134.845 16.530 ;
        RECT 135.910 16.110 136.330 16.530 ;
        RECT 136.520 16.110 136.940 16.530 ;
        RECT 137.130 16.110 137.550 16.530 ;
        RECT 137.740 16.110 138.160 16.530 ;
        RECT 138.350 16.110 138.770 16.530 ;
        RECT 139.825 16.110 140.245 16.530 ;
        RECT 140.435 16.110 140.855 16.530 ;
        RECT 141.045 16.110 141.465 16.530 ;
        RECT 141.655 16.110 142.170 16.530 ;
        RECT 150.470 16.110 150.985 16.530 ;
        RECT 151.175 16.110 151.595 16.530 ;
        RECT 151.785 16.110 152.205 16.530 ;
        RECT 152.395 16.110 152.815 16.530 ;
        RECT 153.615 16.110 154.035 16.530 ;
        RECT 154.225 16.110 154.645 16.530 ;
        RECT 154.835 16.110 155.255 16.530 ;
        RECT 155.445 16.110 155.960 16.530 ;
        RECT 123.415 6.435 124.035 7.155 ;
        RECT 128.900 6.500 129.930 7.090 ;
        RECT 130.120 6.500 130.570 7.090 ;
        RECT 109.650 -0.210 110.165 0.210 ;
        RECT 110.355 -0.210 110.775 0.210 ;
        RECT 110.965 -0.210 111.385 0.210 ;
        RECT 111.575 -0.210 111.995 0.210 ;
        RECT 113.050 -0.210 113.470 0.210 ;
        RECT 113.660 -0.210 114.080 0.210 ;
        RECT 114.270 -0.210 114.690 0.210 ;
        RECT 114.880 -0.210 115.300 0.210 ;
        RECT 115.490 -0.210 115.910 0.210 ;
        RECT 116.975 -0.210 117.395 0.210 ;
        RECT 117.585 -0.210 118.005 0.210 ;
        RECT 118.195 -0.210 118.615 0.210 ;
        RECT 118.805 -0.210 119.320 0.210 ;
        RECT 125.355 -0.210 125.775 0.210 ;
        RECT 125.965 -0.210 126.385 0.210 ;
        RECT 126.575 -0.210 126.995 0.210 ;
        RECT 127.185 -0.210 127.700 0.210 ;
        RECT 128.500 -0.210 129.015 0.210 ;
        RECT 129.205 -0.210 129.625 0.210 ;
        RECT 129.815 -0.210 130.235 0.210 ;
        RECT 130.425 -0.210 130.845 0.210 ;
        RECT 147.060 6.320 148.070 7.260 ;
        RECT 162.000 16.110 162.515 16.530 ;
        RECT 162.705 16.110 163.125 16.530 ;
        RECT 163.315 16.110 163.735 16.530 ;
        RECT 163.925 16.110 164.345 16.530 ;
        RECT 165.410 16.110 165.830 16.530 ;
        RECT 166.020 16.110 166.440 16.530 ;
        RECT 166.630 16.110 167.050 16.530 ;
        RECT 167.240 16.110 167.660 16.530 ;
        RECT 167.850 16.110 168.270 16.530 ;
        RECT 169.325 16.110 169.745 16.530 ;
        RECT 169.935 16.110 170.355 16.530 ;
        RECT 170.545 16.110 170.965 16.530 ;
        RECT 171.155 16.110 171.670 16.530 ;
        RECT 152.915 6.435 153.535 7.155 ;
        RECT 158.400 6.500 159.430 7.090 ;
        RECT 159.620 6.500 160.070 7.090 ;
        RECT 139.150 -0.210 139.665 0.210 ;
        RECT 139.855 -0.210 140.275 0.210 ;
        RECT 140.465 -0.210 140.885 0.210 ;
        RECT 141.075 -0.210 141.495 0.210 ;
        RECT 142.550 -0.210 142.970 0.210 ;
        RECT 143.160 -0.210 143.580 0.210 ;
        RECT 143.770 -0.210 144.190 0.210 ;
        RECT 144.380 -0.210 144.800 0.210 ;
        RECT 144.990 -0.210 145.410 0.210 ;
        RECT 146.475 -0.210 146.895 0.210 ;
        RECT 147.085 -0.210 147.505 0.210 ;
        RECT 147.695 -0.210 148.115 0.210 ;
        RECT 148.305 -0.210 148.820 0.210 ;
        RECT 154.855 -0.210 155.275 0.210 ;
        RECT 155.465 -0.210 155.885 0.210 ;
        RECT 156.075 -0.210 156.495 0.210 ;
        RECT 156.685 -0.210 157.200 0.210 ;
        RECT 158.000 -0.210 158.515 0.210 ;
        RECT 158.705 -0.210 159.125 0.210 ;
        RECT 159.315 -0.210 159.735 0.210 ;
        RECT 159.925 -0.210 160.345 0.210 ;
        RECT 176.560 6.320 177.570 7.260 ;
        RECT 168.650 -0.210 169.165 0.210 ;
        RECT 169.355 -0.210 169.775 0.210 ;
        RECT 169.965 -0.210 170.385 0.210 ;
        RECT 170.575 -0.210 170.995 0.210 ;
        RECT 172.050 -0.210 172.470 0.210 ;
        RECT 172.660 -0.210 173.080 0.210 ;
        RECT 173.270 -0.210 173.690 0.210 ;
        RECT 173.880 -0.210 174.300 0.210 ;
        RECT 174.490 -0.210 174.910 0.210 ;
        RECT 175.975 -0.210 176.395 0.210 ;
        RECT 176.585 -0.210 177.005 0.210 ;
        RECT 177.195 -0.210 177.615 0.210 ;
        RECT 177.805 -0.210 178.320 0.210 ;
      LAYER met1 ;
        RECT 2.000 37.840 173.490 38.320 ;
        RECT 19.290 31.615 20.420 31.840 ;
        RECT 43.295 31.615 44.035 31.675 ;
        RECT 48.790 31.615 49.920 31.840 ;
        RECT 72.795 31.615 73.535 31.675 ;
        RECT 78.290 31.615 79.420 31.840 ;
        RECT 102.295 31.615 103.035 31.675 ;
        RECT 107.790 31.615 108.920 31.840 ;
        RECT 131.795 31.615 132.535 31.675 ;
        RECT 137.290 31.615 138.420 31.840 ;
        RECT 161.295 31.615 162.035 31.675 ;
        RECT 17.840 30.955 20.420 31.615 ;
        RECT 35.060 31.610 49.920 31.615 ;
        RECT 64.560 31.610 79.420 31.615 ;
        RECT 94.060 31.610 108.920 31.615 ;
        RECT 123.560 31.610 138.420 31.615 ;
        RECT 153.060 31.610 165.440 31.615 ;
        RECT 19.290 30.740 20.420 30.955 ;
        RECT 25.290 30.955 49.920 31.610 ;
        RECT 25.290 30.950 38.550 30.955 ;
        RECT 43.295 30.895 44.035 30.955 ;
        RECT 48.790 30.740 49.920 30.955 ;
        RECT 54.790 30.955 79.420 31.610 ;
        RECT 54.790 30.950 68.050 30.955 ;
        RECT 72.795 30.895 73.535 30.955 ;
        RECT 78.290 30.740 79.420 30.955 ;
        RECT 84.290 30.955 108.920 31.610 ;
        RECT 84.290 30.950 97.550 30.955 ;
        RECT 102.295 30.895 103.035 30.955 ;
        RECT 107.790 30.740 108.920 30.955 ;
        RECT 113.790 30.955 138.420 31.610 ;
        RECT 113.790 30.950 127.050 30.955 ;
        RECT 131.795 30.895 132.535 30.955 ;
        RECT 137.290 30.740 138.420 30.955 ;
        RECT 143.290 30.955 165.440 31.610 ;
        RECT 143.290 30.950 156.550 30.955 ;
        RECT 161.295 30.895 162.035 30.955 ;
        RECT 17.890 21.990 165.390 22.000 ;
        RECT 2.000 21.510 177.530 21.990 ;
        RECT 175.570 21.160 177.530 21.510 ;
        RECT 2.000 16.080 180.440 16.560 ;
        RECT 5.355 7.125 6.095 7.185 ;
        RECT 10.840 7.125 24.100 7.130 ;
        RECT 2.000 6.470 24.100 7.125 ;
        RECT 28.970 7.125 30.100 7.340 ;
        RECT 34.855 7.125 35.595 7.185 ;
        RECT 40.340 7.125 53.600 7.130 ;
        RECT 28.970 6.470 53.600 7.125 ;
        RECT 58.470 7.125 59.600 7.340 ;
        RECT 64.355 7.125 65.095 7.185 ;
        RECT 69.840 7.125 83.100 7.130 ;
        RECT 58.470 6.470 83.100 7.125 ;
        RECT 87.970 7.125 89.100 7.340 ;
        RECT 93.855 7.125 94.595 7.185 ;
        RECT 99.340 7.125 112.600 7.130 ;
        RECT 87.970 6.470 112.600 7.125 ;
        RECT 117.470 7.125 118.600 7.340 ;
        RECT 123.355 7.125 124.095 7.185 ;
        RECT 128.840 7.125 142.100 7.130 ;
        RECT 117.470 6.470 142.100 7.125 ;
        RECT 146.970 7.125 148.100 7.340 ;
        RECT 152.855 7.125 153.595 7.185 ;
        RECT 158.340 7.125 171.600 7.130 ;
        RECT 146.970 6.470 171.600 7.125 ;
        RECT 176.470 7.125 177.600 7.340 ;
        RECT 176.470 7.095 179.000 7.125 ;
        RECT 172.640 6.495 179.000 7.095 ;
        RECT 2.000 6.465 14.330 6.470 ;
        RECT 28.970 6.465 43.830 6.470 ;
        RECT 58.470 6.465 73.330 6.470 ;
        RECT 87.970 6.465 102.830 6.470 ;
        RECT 117.470 6.465 132.330 6.470 ;
        RECT 146.970 6.465 161.830 6.470 ;
        RECT 176.470 6.465 179.000 6.495 ;
        RECT 5.355 6.405 6.095 6.465 ;
        RECT 28.970 6.240 30.100 6.465 ;
        RECT 34.855 6.405 35.595 6.465 ;
        RECT 58.470 6.240 59.600 6.465 ;
        RECT 64.355 6.405 65.095 6.465 ;
        RECT 87.970 6.240 89.100 6.465 ;
        RECT 93.855 6.405 94.595 6.465 ;
        RECT 117.470 6.240 118.600 6.465 ;
        RECT 123.355 6.405 124.095 6.465 ;
        RECT 146.970 6.240 148.100 6.465 ;
        RECT 152.855 6.405 153.595 6.465 ;
        RECT 176.470 6.240 177.600 6.465 ;
        RECT 2.000 -0.240 180.440 0.240 ;
      LAYER via ;
        RECT 172.440 37.840 173.440 38.320 ;
        RECT 17.890 30.955 18.785 31.615 ;
        RECT 164.470 30.955 165.390 31.615 ;
        RECT 172.440 21.510 174.440 21.990 ;
        RECT 179.440 16.080 180.390 16.560 ;
        RECT 3.995 6.465 4.695 7.125 ;
        RECT 172.700 6.495 173.400 7.095 ;
        RECT 179.440 -0.240 180.410 0.240 ;
      LAYER met2 ;
        RECT 17.890 31.635 18.785 31.665 ;
        RECT 14.420 30.935 18.785 31.635 ;
        RECT 14.420 20.050 15.120 30.935 ;
        RECT 17.890 30.905 18.785 30.935 ;
        RECT 164.470 31.635 165.390 31.665 ;
        RECT 164.470 30.935 169.490 31.635 ;
        RECT 164.470 30.905 165.390 30.935 ;
        RECT 4.000 19.350 15.120 20.050 ;
        RECT 4.000 18.535 4.700 19.350 ;
        RECT 3.995 12.965 4.700 18.535 ;
        RECT 168.790 17.635 169.490 30.935 ;
        RECT 172.440 22.240 173.440 38.370 ;
        RECT 172.440 21.240 180.440 22.240 ;
        RECT 179.440 20.700 180.435 21.240 ;
        RECT 168.790 16.935 173.400 17.635 ;
        RECT 3.995 6.415 4.695 12.965 ;
        RECT 172.700 6.445 173.400 16.935 ;
        RECT 179.440 -0.290 180.440 20.700 ;
  END
END ring_osc_3-1
MACRO power_ring
  CLASS BLOCK ;
  FOREIGN power_ring ;
  ORIGIN -63.000 24.000 ;
  SIZE 291.000 BY 133.000 ;
  OBS
      LAYER met4 ;
        RECT 63.000 -24.000 65.000 109.000 ;
        RECT 69.000 -19.000 71.000 104.000 ;
        RECT 79.000 -24.000 81.000 109.000 ;
        RECT 99.000 -19.000 101.000 104.000 ;
        RECT 117.000 -24.000 119.000 109.000 ;
        RECT 135.000 -19.000 137.000 104.000 ;
        RECT 153.000 -24.000 155.000 109.000 ;
        RECT 171.000 -19.000 173.000 104.000 ;
        RECT 189.000 -24.000 191.000 109.000 ;
        RECT 207.000 -19.000 209.000 104.000 ;
        RECT 225.000 -24.000 227.000 109.000 ;
        RECT 243.000 -19.000 245.000 104.000 ;
        RECT 261.000 -24.000 263.000 109.000 ;
        RECT 279.000 -19.000 281.000 104.000 ;
        RECT 297.000 -24.000 299.000 109.000 ;
        RECT 315.000 -19.000 317.000 104.000 ;
        RECT 336.000 -24.000 338.000 109.000 ;
        RECT 346.000 -19.000 348.000 104.000 ;
        RECT 352.000 -24.000 354.000 109.000 ;
      LAYER via4 ;
        RECT 63.250 107.250 64.750 108.750 ;
        RECT 79.250 107.250 80.750 108.750 ;
        RECT 69.250 102.250 70.750 103.750 ;
        RECT 69.250 -18.750 70.750 -17.250 ;
        RECT 63.250 -23.750 64.750 -22.250 ;
        RECT 117.250 107.250 118.750 108.750 ;
        RECT 99.250 102.250 100.750 103.750 ;
        RECT 99.250 -18.750 100.750 -17.250 ;
        RECT 79.250 -23.750 80.750 -22.250 ;
        RECT 153.250 107.250 154.750 108.750 ;
        RECT 135.250 102.250 136.750 103.750 ;
        RECT 135.250 -18.750 136.750 -17.250 ;
        RECT 117.250 -23.750 118.750 -22.250 ;
        RECT 189.250 107.250 190.750 108.750 ;
        RECT 171.250 102.250 172.750 103.750 ;
        RECT 171.250 -18.750 172.750 -17.250 ;
        RECT 153.250 -23.750 154.750 -22.250 ;
        RECT 225.250 107.250 226.750 108.750 ;
        RECT 207.250 102.250 208.750 103.750 ;
        RECT 207.250 -18.750 208.750 -17.250 ;
        RECT 189.250 -23.750 190.750 -22.250 ;
        RECT 261.250 107.250 262.750 108.750 ;
        RECT 243.250 102.250 244.750 103.750 ;
        RECT 243.250 -18.750 244.750 -17.250 ;
        RECT 225.250 -23.750 226.750 -22.250 ;
        RECT 297.250 107.250 298.750 108.750 ;
        RECT 279.250 102.250 280.750 103.750 ;
        RECT 279.250 -18.750 280.750 -17.250 ;
        RECT 261.250 -23.750 262.750 -22.250 ;
        RECT 336.250 107.250 337.750 108.750 ;
        RECT 315.250 102.250 316.750 103.750 ;
        RECT 315.250 -18.750 316.750 -17.250 ;
        RECT 297.250 -23.750 298.750 -22.250 ;
        RECT 352.250 107.250 353.750 108.750 ;
        RECT 346.250 102.250 347.750 103.750 ;
        RECT 346.250 -18.750 347.750 -17.250 ;
        RECT 336.250 -23.750 337.750 -22.250 ;
        RECT 352.250 -23.750 353.750 -22.250 ;
      LAYER met5 ;
        RECT 63.000 107.000 354.000 109.000 ;
        RECT 69.000 102.000 348.000 104.000 ;
        RECT 69.000 -19.000 348.000 -17.000 ;
        RECT 63.000 -24.000 354.000 -22.000 ;
  END
END power_ring
MACRO vco
  CLASS BLOCK ;
  FOREIGN vco ;
  ORIGIN 0.000 0.000 ;
  SIZE 291.000 BY 133.000 ;
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 204.810 56.170 206.010 56.750 ;
        RECT 204.010 56.050 206.010 56.170 ;
        RECT 222.780 56.110 223.960 56.390 ;
        RECT 204.010 55.450 208.010 56.050 ;
        RECT 222.280 55.510 223.960 56.110 ;
        RECT 222.780 55.310 223.960 55.510 ;
        RECT 226.445 55.020 226.945 56.170 ;
        RECT 228.960 55.020 229.255 59.285 ;
        RECT 236.110 56.750 236.400 62.080 ;
        RECT 240.290 56.750 240.580 62.080 ;
        RECT 236.110 56.460 240.580 56.750 ;
        RECT 238.540 55.020 239.040 56.460 ;
        RECT 226.445 54.520 239.040 55.020 ;
        RECT 228.965 46.840 229.260 54.520 ;
        RECT 236.110 49.520 236.400 54.520 ;
      LAYER mcon ;
        RECT 204.070 55.510 204.710 56.140 ;
        RECT 204.910 55.450 205.610 56.140 ;
        RECT 205.810 55.450 206.410 56.050 ;
        RECT 206.610 55.450 207.210 56.050 ;
        RECT 207.410 55.450 208.010 56.050 ;
        RECT 222.330 55.560 222.730 56.060 ;
        RECT 222.930 55.560 223.880 56.060 ;
        RECT 226.445 55.510 226.945 56.110 ;
      LAYER met1 ;
        RECT 204.010 56.110 208.110 56.170 ;
        RECT 226.415 56.110 226.975 56.170 ;
        RECT 204.010 55.510 226.975 56.110 ;
        RECT 204.010 55.450 208.110 55.510 ;
        RECT 226.415 55.450 226.975 55.510 ;
        RECT 204.810 55.420 208.110 55.450 ;
      LAYER via ;
        RECT 220.510 55.510 221.110 56.110 ;
        RECT 221.250 55.510 221.850 56.110 ;
      LAYER met2 ;
        RECT 220.510 55.480 221.850 56.160 ;
        RECT 220.780 45.000 221.580 55.480 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 175.310 56.170 176.510 56.750 ;
        RECT 174.510 56.050 176.510 56.170 ;
        RECT 193.280 56.110 194.460 56.390 ;
        RECT 174.510 55.450 178.510 56.050 ;
        RECT 192.780 55.510 194.460 56.110 ;
        RECT 193.280 55.310 194.460 55.510 ;
        RECT 196.945 55.020 197.445 56.170 ;
        RECT 199.460 55.020 199.755 59.285 ;
        RECT 206.610 56.750 206.900 62.080 ;
        RECT 210.790 56.750 211.080 62.080 ;
        RECT 206.610 56.460 211.080 56.750 ;
        RECT 209.040 55.020 209.540 56.460 ;
        RECT 196.945 54.520 209.540 55.020 ;
        RECT 199.465 46.840 199.760 54.520 ;
        RECT 206.610 49.520 206.900 54.520 ;
      LAYER mcon ;
        RECT 174.570 55.510 175.210 56.140 ;
        RECT 175.410 55.450 176.110 56.140 ;
        RECT 176.310 55.450 176.910 56.050 ;
        RECT 177.110 55.450 177.710 56.050 ;
        RECT 177.910 55.450 178.510 56.050 ;
        RECT 192.830 55.560 193.230 56.060 ;
        RECT 193.430 55.560 194.380 56.060 ;
        RECT 196.945 55.510 197.445 56.110 ;
      LAYER met1 ;
        RECT 174.510 56.110 178.610 56.170 ;
        RECT 196.915 56.110 197.475 56.170 ;
        RECT 174.510 55.510 197.475 56.110 ;
        RECT 174.510 55.450 178.610 55.510 ;
        RECT 196.915 55.450 197.475 55.510 ;
        RECT 175.310 55.420 178.610 55.450 ;
      LAYER via ;
        RECT 191.010 55.510 191.610 56.110 ;
        RECT 191.750 55.510 192.350 56.110 ;
      LAYER met2 ;
        RECT 191.010 55.480 192.350 56.160 ;
        RECT 191.280 45.000 192.080 55.480 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 145.810 56.170 147.010 56.750 ;
        RECT 145.010 56.050 147.010 56.170 ;
        RECT 163.780 56.110 164.960 56.390 ;
        RECT 145.010 55.450 149.010 56.050 ;
        RECT 163.280 55.510 164.960 56.110 ;
        RECT 163.780 55.310 164.960 55.510 ;
        RECT 167.445 55.020 167.945 56.170 ;
        RECT 169.960 55.020 170.255 59.285 ;
        RECT 177.110 56.750 177.400 62.080 ;
        RECT 181.290 56.750 181.580 62.080 ;
        RECT 177.110 56.460 181.580 56.750 ;
        RECT 179.540 55.020 180.040 56.460 ;
        RECT 167.445 54.520 180.040 55.020 ;
        RECT 169.965 46.840 170.260 54.520 ;
        RECT 177.110 49.520 177.400 54.520 ;
      LAYER mcon ;
        RECT 145.070 55.510 145.710 56.140 ;
        RECT 145.910 55.450 146.610 56.140 ;
        RECT 146.810 55.450 147.410 56.050 ;
        RECT 147.610 55.450 148.210 56.050 ;
        RECT 148.410 55.450 149.010 56.050 ;
        RECT 163.330 55.560 163.730 56.060 ;
        RECT 163.930 55.560 164.880 56.060 ;
        RECT 167.445 55.510 167.945 56.110 ;
      LAYER met1 ;
        RECT 145.010 56.110 149.110 56.170 ;
        RECT 167.415 56.110 167.975 56.170 ;
        RECT 145.010 55.510 167.975 56.110 ;
        RECT 145.010 55.450 149.110 55.510 ;
        RECT 167.415 55.450 167.975 55.510 ;
        RECT 145.810 55.420 149.110 55.450 ;
      LAYER via ;
        RECT 161.510 55.510 162.110 56.110 ;
        RECT 162.250 55.510 162.850 56.110 ;
      LAYER met2 ;
        RECT 161.510 55.480 162.850 56.160 ;
        RECT 161.780 45.000 162.580 55.480 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 116.310 56.170 117.510 56.750 ;
        RECT 115.510 56.050 117.510 56.170 ;
        RECT 134.280 56.110 135.460 56.390 ;
        RECT 115.510 55.450 119.510 56.050 ;
        RECT 133.780 55.510 135.460 56.110 ;
        RECT 134.280 55.310 135.460 55.510 ;
        RECT 137.945 55.020 138.445 56.170 ;
        RECT 140.460 55.020 140.755 59.285 ;
        RECT 147.610 56.750 147.900 62.080 ;
        RECT 151.790 56.750 152.080 62.080 ;
        RECT 147.610 56.460 152.080 56.750 ;
        RECT 150.040 55.020 150.540 56.460 ;
        RECT 137.945 54.520 150.540 55.020 ;
        RECT 140.465 46.840 140.760 54.520 ;
        RECT 147.610 49.520 147.900 54.520 ;
      LAYER mcon ;
        RECT 115.570 55.510 116.210 56.140 ;
        RECT 116.410 55.450 117.110 56.140 ;
        RECT 117.310 55.450 117.910 56.050 ;
        RECT 118.110 55.450 118.710 56.050 ;
        RECT 118.910 55.450 119.510 56.050 ;
        RECT 133.830 55.560 134.230 56.060 ;
        RECT 134.430 55.560 135.380 56.060 ;
        RECT 137.945 55.510 138.445 56.110 ;
      LAYER met1 ;
        RECT 115.510 56.110 119.610 56.170 ;
        RECT 137.915 56.110 138.475 56.170 ;
        RECT 115.510 55.510 138.475 56.110 ;
        RECT 115.510 55.450 119.610 55.510 ;
        RECT 137.915 55.450 138.475 55.510 ;
        RECT 116.310 55.420 119.610 55.450 ;
      LAYER via ;
        RECT 132.010 55.510 132.610 56.110 ;
        RECT 132.750 55.510 133.350 56.110 ;
      LAYER met2 ;
        RECT 132.010 55.480 133.350 56.160 ;
        RECT 132.280 45.000 133.080 55.480 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 86.810 56.170 88.010 56.750 ;
        RECT 86.010 56.050 88.010 56.170 ;
        RECT 104.780 56.110 105.960 56.390 ;
        RECT 86.010 55.450 90.010 56.050 ;
        RECT 104.280 55.510 105.960 56.110 ;
        RECT 104.780 55.310 105.960 55.510 ;
        RECT 108.445 55.020 108.945 56.170 ;
        RECT 110.960 55.020 111.255 59.285 ;
        RECT 118.110 56.750 118.400 62.080 ;
        RECT 122.290 56.750 122.580 62.080 ;
        RECT 118.110 56.460 122.580 56.750 ;
        RECT 120.540 55.020 121.040 56.460 ;
        RECT 108.445 54.520 121.040 55.020 ;
        RECT 110.965 46.840 111.260 54.520 ;
        RECT 118.110 49.520 118.400 54.520 ;
      LAYER mcon ;
        RECT 86.070 55.510 86.710 56.140 ;
        RECT 86.910 55.450 87.610 56.140 ;
        RECT 87.810 55.450 88.410 56.050 ;
        RECT 88.610 55.450 89.210 56.050 ;
        RECT 89.410 55.450 90.010 56.050 ;
        RECT 104.330 55.560 104.730 56.060 ;
        RECT 104.930 55.560 105.880 56.060 ;
        RECT 108.445 55.510 108.945 56.110 ;
      LAYER met1 ;
        RECT 86.010 56.110 90.110 56.170 ;
        RECT 108.415 56.110 108.975 56.170 ;
        RECT 86.010 55.510 108.975 56.110 ;
        RECT 86.010 55.450 90.110 55.510 ;
        RECT 108.415 55.450 108.975 55.510 ;
        RECT 86.810 55.420 90.110 55.450 ;
      LAYER via ;
        RECT 102.510 55.510 103.110 56.110 ;
        RECT 103.250 55.510 103.850 56.110 ;
      LAYER met2 ;
        RECT 102.510 55.480 103.850 56.160 ;
        RECT 102.780 45.000 103.580 55.480 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 102.400 74.610 106.400 75.210 ;
        RECT 104.400 74.490 106.400 74.610 ;
        RECT 104.400 73.910 105.600 74.490 ;
        RECT 75.280 56.110 76.460 56.390 ;
        RECT 74.780 55.510 76.460 56.110 ;
        RECT 75.280 55.310 76.460 55.510 ;
        RECT 78.945 55.020 79.445 56.170 ;
        RECT 81.460 55.020 81.755 59.285 ;
        RECT 88.610 56.750 88.900 62.080 ;
        RECT 92.790 56.750 93.080 62.080 ;
        RECT 88.610 56.460 93.080 56.750 ;
        RECT 91.040 55.020 91.540 56.460 ;
        RECT 78.945 54.520 91.540 55.020 ;
        RECT 81.465 46.840 81.760 54.520 ;
        RECT 88.610 49.520 88.900 54.520 ;
      LAYER mcon ;
        RECT 102.400 74.610 103.000 75.210 ;
        RECT 103.200 74.610 103.800 75.210 ;
        RECT 104.000 74.610 104.600 75.210 ;
        RECT 104.800 74.520 105.500 75.210 ;
        RECT 105.700 74.520 106.340 75.150 ;
        RECT 74.830 55.560 75.230 56.060 ;
        RECT 75.430 55.560 76.380 56.060 ;
        RECT 78.945 55.510 79.445 56.110 ;
      LAYER met1 ;
        RECT 102.300 75.210 105.600 75.240 ;
        RECT 102.300 75.150 106.400 75.210 ;
        RECT 89.350 74.550 106.400 75.150 ;
        RECT 102.300 74.490 106.400 74.550 ;
        RECT 78.915 56.110 79.475 56.170 ;
        RECT 73.510 55.510 79.475 56.110 ;
        RECT 78.915 55.450 79.475 55.510 ;
      LAYER via ;
        RECT 89.400 74.550 90.375 75.150 ;
        RECT 78.215 55.510 78.915 56.110 ;
      LAYER met2 ;
        RECT 88.630 74.500 90.375 75.200 ;
        RECT 88.630 63.640 89.330 74.500 ;
        RECT 78.215 62.940 89.330 63.640 ;
        RECT 78.215 55.460 78.915 62.940 ;
        RECT 84.780 45.000 85.580 62.940 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 103.510 76.140 103.800 81.140 ;
        RECT 110.650 76.140 110.945 83.820 ;
        RECT 100.870 75.640 113.465 76.140 ;
        RECT 100.870 74.200 101.370 75.640 ;
        RECT 99.330 73.910 103.800 74.200 ;
        RECT 99.330 68.580 99.620 73.910 ;
        RECT 103.510 68.580 103.800 73.910 ;
        RECT 110.655 71.375 110.950 75.640 ;
        RECT 112.965 74.490 113.465 75.640 ;
        RECT 115.950 75.150 117.130 75.350 ;
        RECT 115.950 74.550 117.630 75.150 ;
        RECT 131.900 74.610 135.900 75.210 ;
        RECT 115.950 74.270 117.130 74.550 ;
        RECT 133.900 74.490 135.900 74.610 ;
        RECT 133.900 73.910 135.100 74.490 ;
      LAYER mcon ;
        RECT 112.965 74.550 113.465 75.150 ;
        RECT 116.030 74.600 116.980 75.100 ;
        RECT 117.180 74.600 117.580 75.100 ;
        RECT 131.900 74.610 132.500 75.210 ;
        RECT 132.700 74.610 133.300 75.210 ;
        RECT 133.500 74.610 134.100 75.210 ;
        RECT 134.300 74.520 135.000 75.210 ;
        RECT 135.200 74.520 135.840 75.150 ;
      LAYER met1 ;
        RECT 131.800 75.210 135.100 75.240 ;
        RECT 112.935 75.150 113.495 75.210 ;
        RECT 131.800 75.150 135.900 75.210 ;
        RECT 112.935 74.550 135.900 75.150 ;
        RECT 112.935 74.490 113.495 74.550 ;
        RECT 131.800 74.490 135.900 74.550 ;
      LAYER via ;
        RECT 118.060 74.550 118.660 75.150 ;
        RECT 118.800 74.550 119.400 75.150 ;
      LAYER met2 ;
        RECT 118.330 75.210 119.130 85.660 ;
        RECT 118.060 74.500 119.400 75.210 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 133.010 76.140 133.300 81.140 ;
        RECT 140.150 76.140 140.445 83.820 ;
        RECT 130.370 75.640 142.965 76.140 ;
        RECT 130.370 74.200 130.870 75.640 ;
        RECT 128.830 73.910 133.300 74.200 ;
        RECT 128.830 68.580 129.120 73.910 ;
        RECT 133.010 68.580 133.300 73.910 ;
        RECT 140.155 71.375 140.450 75.640 ;
        RECT 142.465 74.490 142.965 75.640 ;
        RECT 145.450 75.150 146.630 75.350 ;
        RECT 145.450 74.550 147.130 75.150 ;
        RECT 161.400 74.610 165.400 75.210 ;
        RECT 145.450 74.270 146.630 74.550 ;
        RECT 163.400 74.490 165.400 74.610 ;
        RECT 163.400 73.910 164.600 74.490 ;
      LAYER mcon ;
        RECT 142.465 74.550 142.965 75.150 ;
        RECT 145.530 74.600 146.480 75.100 ;
        RECT 146.680 74.600 147.080 75.100 ;
        RECT 161.400 74.610 162.000 75.210 ;
        RECT 162.200 74.610 162.800 75.210 ;
        RECT 163.000 74.610 163.600 75.210 ;
        RECT 163.800 74.520 164.500 75.210 ;
        RECT 164.700 74.520 165.340 75.150 ;
      LAYER met1 ;
        RECT 161.300 75.210 164.600 75.240 ;
        RECT 142.435 75.150 142.995 75.210 ;
        RECT 161.300 75.150 165.400 75.210 ;
        RECT 142.435 74.550 165.400 75.150 ;
        RECT 142.435 74.490 142.995 74.550 ;
        RECT 161.300 74.490 165.400 74.550 ;
      LAYER via ;
        RECT 147.560 74.550 148.160 75.150 ;
        RECT 148.300 74.550 148.900 75.150 ;
      LAYER met2 ;
        RECT 147.830 75.210 148.630 85.660 ;
        RECT 147.560 74.500 148.900 75.210 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 162.510 76.140 162.800 81.140 ;
        RECT 169.650 76.140 169.945 83.820 ;
        RECT 159.870 75.640 172.465 76.140 ;
        RECT 159.870 74.200 160.370 75.640 ;
        RECT 158.330 73.910 162.800 74.200 ;
        RECT 158.330 68.580 158.620 73.910 ;
        RECT 162.510 68.580 162.800 73.910 ;
        RECT 169.655 71.375 169.950 75.640 ;
        RECT 171.965 74.490 172.465 75.640 ;
        RECT 174.950 75.150 176.130 75.350 ;
        RECT 174.950 74.550 176.630 75.150 ;
        RECT 190.900 74.610 194.900 75.210 ;
        RECT 174.950 74.270 176.130 74.550 ;
        RECT 192.900 74.490 194.900 74.610 ;
        RECT 192.900 73.910 194.100 74.490 ;
      LAYER mcon ;
        RECT 171.965 74.550 172.465 75.150 ;
        RECT 175.030 74.600 175.980 75.100 ;
        RECT 176.180 74.600 176.580 75.100 ;
        RECT 190.900 74.610 191.500 75.210 ;
        RECT 191.700 74.610 192.300 75.210 ;
        RECT 192.500 74.610 193.100 75.210 ;
        RECT 193.300 74.520 194.000 75.210 ;
        RECT 194.200 74.520 194.840 75.150 ;
      LAYER met1 ;
        RECT 190.800 75.210 194.100 75.240 ;
        RECT 171.935 75.150 172.495 75.210 ;
        RECT 190.800 75.150 194.900 75.210 ;
        RECT 171.935 74.550 194.900 75.150 ;
        RECT 171.935 74.490 172.495 74.550 ;
        RECT 190.800 74.490 194.900 74.550 ;
      LAYER via ;
        RECT 177.060 74.550 177.660 75.150 ;
        RECT 177.800 74.550 178.400 75.150 ;
      LAYER met2 ;
        RECT 177.330 75.210 178.130 85.660 ;
        RECT 177.060 74.500 178.400 75.210 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 192.010 76.140 192.300 81.140 ;
        RECT 199.150 76.140 199.445 83.820 ;
        RECT 189.370 75.640 201.965 76.140 ;
        RECT 189.370 74.200 189.870 75.640 ;
        RECT 187.830 73.910 192.300 74.200 ;
        RECT 187.830 68.580 188.120 73.910 ;
        RECT 192.010 68.580 192.300 73.910 ;
        RECT 199.155 71.375 199.450 75.640 ;
        RECT 201.465 74.490 201.965 75.640 ;
        RECT 204.450 75.150 205.630 75.350 ;
        RECT 204.450 74.550 206.130 75.150 ;
        RECT 220.400 74.610 224.400 75.210 ;
        RECT 204.450 74.270 205.630 74.550 ;
        RECT 222.400 74.490 224.400 74.610 ;
        RECT 222.400 73.910 223.600 74.490 ;
      LAYER mcon ;
        RECT 201.465 74.550 201.965 75.150 ;
        RECT 204.530 74.600 205.480 75.100 ;
        RECT 205.680 74.600 206.080 75.100 ;
        RECT 220.400 74.610 221.000 75.210 ;
        RECT 221.200 74.610 221.800 75.210 ;
        RECT 222.000 74.610 222.600 75.210 ;
        RECT 222.800 74.520 223.500 75.210 ;
        RECT 223.700 74.520 224.340 75.150 ;
      LAYER met1 ;
        RECT 220.300 75.210 223.600 75.240 ;
        RECT 201.435 75.150 201.995 75.210 ;
        RECT 220.300 75.150 224.400 75.210 ;
        RECT 201.435 74.550 224.400 75.150 ;
        RECT 201.435 74.490 201.995 74.550 ;
        RECT 220.300 74.490 224.400 74.550 ;
      LAYER via ;
        RECT 206.560 74.550 207.160 75.150 ;
        RECT 207.300 74.550 207.900 75.150 ;
      LAYER met2 ;
        RECT 206.830 75.210 207.630 85.660 ;
        RECT 206.560 74.500 207.900 75.210 ;
    END
  END p[9]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER li1 ;
        RECT 221.510 76.140 221.800 81.140 ;
        RECT 228.650 76.140 228.945 83.820 ;
        RECT 218.870 75.640 231.465 76.140 ;
        RECT 218.870 74.200 219.370 75.640 ;
        RECT 217.330 73.910 221.800 74.200 ;
        RECT 217.330 68.580 217.620 73.910 ;
        RECT 221.510 68.580 221.800 73.910 ;
        RECT 228.655 71.375 228.950 75.640 ;
        RECT 230.965 74.490 231.465 75.640 ;
        RECT 233.950 75.150 235.130 75.350 ;
        RECT 233.950 74.550 235.630 75.150 ;
        RECT 233.950 74.270 235.130 74.550 ;
        RECT 234.310 56.170 235.510 56.750 ;
        RECT 233.510 56.050 235.510 56.170 ;
        RECT 233.510 55.450 237.510 56.050 ;
      LAYER mcon ;
        RECT 230.965 74.550 231.465 75.150 ;
        RECT 234.030 74.600 234.980 75.100 ;
        RECT 235.180 74.600 235.580 75.100 ;
        RECT 233.570 55.510 234.210 56.140 ;
        RECT 234.410 55.450 235.110 56.140 ;
        RECT 235.310 55.450 235.910 56.050 ;
        RECT 236.110 55.450 236.710 56.050 ;
        RECT 236.910 55.450 237.510 56.050 ;
      LAYER met1 ;
        RECT 230.935 75.150 231.495 75.210 ;
        RECT 230.935 74.550 236.950 75.150 ;
        RECT 230.935 74.490 231.495 74.550 ;
        RECT 233.510 56.110 237.610 56.170 ;
        RECT 233.510 55.510 250.510 56.110 ;
        RECT 233.510 55.450 237.610 55.510 ;
        RECT 234.310 55.420 237.610 55.450 ;
      LAYER via ;
        RECT 235.960 74.550 236.900 75.150 ;
        RECT 237.600 55.510 238.300 56.110 ;
        RECT 238.370 55.510 238.970 56.110 ;
      LAYER met2 ;
        RECT 235.960 74.500 238.300 75.200 ;
        RECT 237.600 56.160 238.300 74.500 ;
        RECT 237.600 55.430 238.970 56.160 ;
        RECT 237.870 45.000 238.670 55.430 ;
    END
  END p[10]
  PIN input_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 247.060 72.030 249.060 72.200 ;
        RECT 247.140 72.000 248.980 72.030 ;
      LAYER met1 ;
        RECT 247.030 71.970 249.090 72.230 ;
      LAYER via ;
        RECT 247.080 71.970 249.040 72.230 ;
      LAYER met2 ;
        RECT 247.080 71.680 253.010 72.480 ;
        RECT 247.660 71.490 249.040 71.680 ;
    END
  END input_analog
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
        RECT 198.000 84.130 200.000 84.610 ;
        RECT 90.000 81.410 92.000 81.890 ;
        RECT 126.000 81.410 128.000 81.890 ;
        RECT 162.000 81.410 164.000 81.890 ;
        RECT 234.000 81.410 236.000 81.890 ;
        RECT 90.000 70.530 92.000 71.010 ;
        RECT 126.000 70.530 128.000 71.010 ;
        RECT 198.000 70.530 200.000 71.010 ;
        RECT 234.000 67.800 236.000 68.280 ;
        RECT 234.000 62.370 236.000 62.850 ;
        RECT 90.000 59.650 92.000 60.130 ;
        RECT 126.000 59.650 128.000 60.130 ;
        RECT 162.000 59.650 164.000 60.130 ;
        RECT 198.000 59.650 200.000 60.130 ;
        RECT 90.000 48.770 92.000 49.250 ;
        RECT 126.000 48.770 128.000 49.250 ;
        RECT 198.000 48.770 200.000 49.250 ;
        RECT 234.000 48.770 236.000 49.250 ;
      LAYER via3 ;
        RECT 198.160 84.190 198.520 84.550 ;
        RECT 198.600 84.190 198.960 84.550 ;
        RECT 199.040 84.190 199.400 84.550 ;
        RECT 199.480 84.190 199.840 84.550 ;
        RECT 90.160 81.470 90.520 81.830 ;
        RECT 90.600 81.470 90.960 81.830 ;
        RECT 91.040 81.470 91.400 81.830 ;
        RECT 91.480 81.470 91.840 81.830 ;
        RECT 126.160 81.470 126.520 81.830 ;
        RECT 126.600 81.470 126.960 81.830 ;
        RECT 127.040 81.470 127.400 81.830 ;
        RECT 127.480 81.470 127.840 81.830 ;
        RECT 162.160 81.470 162.520 81.830 ;
        RECT 162.600 81.470 162.960 81.830 ;
        RECT 163.040 81.470 163.400 81.830 ;
        RECT 163.480 81.470 163.840 81.830 ;
        RECT 234.160 81.470 234.520 81.830 ;
        RECT 234.600 81.470 234.960 81.830 ;
        RECT 235.040 81.470 235.400 81.830 ;
        RECT 235.480 81.470 235.840 81.830 ;
        RECT 90.160 70.590 90.520 70.950 ;
        RECT 90.600 70.590 90.960 70.950 ;
        RECT 91.040 70.590 91.400 70.950 ;
        RECT 91.480 70.590 91.840 70.950 ;
        RECT 126.160 70.590 126.520 70.950 ;
        RECT 126.600 70.590 126.960 70.950 ;
        RECT 127.040 70.590 127.400 70.950 ;
        RECT 127.480 70.590 127.840 70.950 ;
        RECT 198.160 70.590 198.520 70.950 ;
        RECT 198.600 70.590 198.960 70.950 ;
        RECT 199.040 70.590 199.400 70.950 ;
        RECT 199.480 70.590 199.840 70.950 ;
        RECT 234.160 67.860 234.520 68.220 ;
        RECT 234.600 67.860 234.960 68.220 ;
        RECT 235.040 67.860 235.400 68.220 ;
        RECT 235.480 67.860 235.840 68.220 ;
        RECT 234.160 62.430 234.520 62.790 ;
        RECT 234.600 62.430 234.960 62.790 ;
        RECT 235.040 62.430 235.400 62.790 ;
        RECT 235.480 62.430 235.840 62.790 ;
        RECT 90.160 59.710 90.520 60.070 ;
        RECT 90.600 59.710 90.960 60.070 ;
        RECT 91.040 59.710 91.400 60.070 ;
        RECT 91.480 59.710 91.840 60.070 ;
        RECT 126.160 59.710 126.520 60.070 ;
        RECT 126.600 59.710 126.960 60.070 ;
        RECT 127.040 59.710 127.400 60.070 ;
        RECT 127.480 59.710 127.840 60.070 ;
        RECT 162.160 59.710 162.520 60.070 ;
        RECT 162.600 59.710 162.960 60.070 ;
        RECT 163.040 59.710 163.400 60.070 ;
        RECT 163.480 59.710 163.840 60.070 ;
        RECT 198.160 59.710 198.520 60.070 ;
        RECT 198.600 59.710 198.960 60.070 ;
        RECT 199.040 59.710 199.400 60.070 ;
        RECT 199.480 59.710 199.840 60.070 ;
        RECT 90.160 48.830 90.520 49.190 ;
        RECT 90.600 48.830 90.960 49.190 ;
        RECT 91.040 48.830 91.400 49.190 ;
        RECT 91.480 48.830 91.840 49.190 ;
        RECT 126.160 48.830 126.520 49.190 ;
        RECT 126.600 48.830 126.960 49.190 ;
        RECT 127.040 48.830 127.400 49.190 ;
        RECT 127.480 48.830 127.840 49.190 ;
        RECT 198.160 48.830 198.520 49.190 ;
        RECT 198.600 48.830 198.960 49.190 ;
        RECT 199.040 48.830 199.400 49.190 ;
        RECT 199.480 48.830 199.840 49.190 ;
        RECT 234.160 48.830 234.520 49.190 ;
        RECT 234.600 48.830 234.960 49.190 ;
        RECT 235.040 48.830 235.400 49.190 ;
        RECT 235.480 48.830 235.840 49.190 ;
      LAYER met4 ;
        RECT 0.000 0.000 2.000 133.000 ;
        RECT 16.000 0.000 18.000 133.000 ;
        RECT 54.000 0.000 56.000 133.000 ;
        RECT 90.000 0.000 92.000 133.000 ;
        RECT 126.000 0.000 128.000 133.000 ;
        RECT 162.000 0.000 164.000 133.000 ;
        RECT 198.000 0.000 200.000 133.000 ;
        RECT 234.000 0.000 236.000 133.000 ;
        RECT 273.000 0.000 275.000 133.000 ;
        RECT 289.000 0.000 291.000 133.000 ;
      LAYER via4 ;
        RECT 0.250 131.250 1.750 132.750 ;
        RECT 0.250 0.250 1.750 1.750 ;
        RECT 16.250 131.250 17.750 132.750 ;
        RECT 16.250 0.250 17.750 1.750 ;
        RECT 54.250 131.250 55.750 132.750 ;
        RECT 54.250 0.250 55.750 1.750 ;
        RECT 90.250 131.250 91.750 132.750 ;
        RECT 90.250 0.250 91.750 1.750 ;
        RECT 126.250 131.250 127.750 132.750 ;
        RECT 126.250 0.250 127.750 1.750 ;
        RECT 162.250 131.250 163.750 132.750 ;
        RECT 162.250 0.250 163.750 1.750 ;
        RECT 198.250 131.250 199.750 132.750 ;
        RECT 198.250 0.250 199.750 1.750 ;
        RECT 234.250 131.250 235.750 132.750 ;
        RECT 234.250 0.250 235.750 1.750 ;
        RECT 273.250 131.250 274.750 132.750 ;
        RECT 273.250 0.250 274.750 1.750 ;
        RECT 289.250 131.250 290.750 132.750 ;
        RECT 289.250 0.250 290.750 1.750 ;
      LAYER met5 ;
        RECT 0.000 131.000 291.000 133.000 ;
        RECT 0.000 0.000 291.000 2.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met3 ;
        RECT 108.000 81.410 110.000 81.890 ;
        RECT 252.000 73.250 254.000 73.730 ;
        RECT 108.000 70.530 110.000 71.010 ;
        RECT 108.000 59.650 110.000 60.130 ;
        RECT 108.000 48.770 110.000 49.250 ;
      LAYER via3 ;
        RECT 108.160 81.470 108.520 81.830 ;
        RECT 108.600 81.470 108.960 81.830 ;
        RECT 109.040 81.470 109.400 81.830 ;
        RECT 109.480 81.470 109.840 81.830 ;
        RECT 252.160 73.310 252.520 73.670 ;
        RECT 252.600 73.310 252.960 73.670 ;
        RECT 253.040 73.310 253.400 73.670 ;
        RECT 253.480 73.310 253.840 73.670 ;
        RECT 108.160 70.590 108.520 70.950 ;
        RECT 108.600 70.590 108.960 70.950 ;
        RECT 109.040 70.590 109.400 70.950 ;
        RECT 109.480 70.590 109.840 70.950 ;
        RECT 108.160 59.710 108.520 60.070 ;
        RECT 108.600 59.710 108.960 60.070 ;
        RECT 109.040 59.710 109.400 60.070 ;
        RECT 109.480 59.710 109.840 60.070 ;
        RECT 108.160 48.830 108.520 49.190 ;
        RECT 108.600 48.830 108.960 49.190 ;
        RECT 109.040 48.830 109.400 49.190 ;
        RECT 109.480 48.830 109.840 49.190 ;
      LAYER met4 ;
        RECT 6.000 5.000 8.000 128.000 ;
        RECT 36.000 5.000 38.000 128.000 ;
        RECT 72.000 5.000 74.000 128.000 ;
        RECT 108.000 5.000 110.000 128.000 ;
        RECT 144.000 5.000 146.000 128.000 ;
        RECT 180.000 5.000 182.000 128.000 ;
        RECT 216.000 5.000 218.000 128.000 ;
        RECT 252.000 5.000 254.000 128.000 ;
        RECT 283.000 5.000 285.000 128.000 ;
      LAYER via4 ;
        RECT 6.250 126.250 7.750 127.750 ;
        RECT 6.250 5.250 7.750 6.750 ;
        RECT 36.250 126.250 37.750 127.750 ;
        RECT 36.250 5.250 37.750 6.750 ;
        RECT 72.250 126.250 73.750 127.750 ;
        RECT 72.250 5.250 73.750 6.750 ;
        RECT 108.250 126.250 109.750 127.750 ;
        RECT 108.250 5.250 109.750 6.750 ;
        RECT 144.250 126.250 145.750 127.750 ;
        RECT 144.250 5.250 145.750 6.750 ;
        RECT 180.250 126.250 181.750 127.750 ;
        RECT 180.250 5.250 181.750 6.750 ;
        RECT 216.250 126.250 217.750 127.750 ;
        RECT 216.250 5.250 217.750 6.750 ;
        RECT 252.250 126.250 253.750 127.750 ;
        RECT 252.250 5.250 253.750 6.750 ;
        RECT 283.250 126.250 284.750 127.750 ;
        RECT 283.250 5.250 284.750 6.750 ;
      LAYER met5 ;
        RECT 6.000 126.000 285.000 128.000 ;
        RECT 6.000 5.000 285.000 7.000 ;
    END
  END vssd1
  OBS
      LAYER pwell ;
        RECT 89.900 78.600 99.930 84.660 ;
      LAYER nwell ;
        RECT 89.900 70.535 95.750 76.410 ;
        RECT 100.730 76.070 106.580 81.925 ;
      LAYER pwell ;
        RECT 107.875 78.560 113.725 84.660 ;
      LAYER nwell ;
        RECT 114.350 76.600 118.110 81.875 ;
      LAYER pwell ;
        RECT 119.400 78.600 129.430 84.660 ;
        RECT 96.550 67.750 106.580 74.150 ;
      LAYER nwell ;
        RECT 107.875 70.540 111.635 75.850 ;
      LAYER pwell ;
        RECT 112.255 72.915 118.105 73.855 ;
        RECT 112.255 72.865 118.110 72.915 ;
        RECT 112.260 67.755 118.110 72.865 ;
      LAYER nwell ;
        RECT 119.400 70.535 125.250 76.410 ;
        RECT 130.230 76.070 136.080 81.925 ;
      LAYER pwell ;
        RECT 137.375 78.560 143.225 84.660 ;
      LAYER nwell ;
        RECT 143.850 76.600 147.610 81.875 ;
      LAYER pwell ;
        RECT 148.900 78.600 158.930 84.660 ;
        RECT 126.050 67.750 136.080 74.150 ;
      LAYER nwell ;
        RECT 137.375 70.540 141.135 75.850 ;
      LAYER pwell ;
        RECT 141.755 72.915 147.605 73.855 ;
        RECT 141.755 72.865 147.610 72.915 ;
        RECT 141.760 67.755 147.610 72.865 ;
      LAYER nwell ;
        RECT 148.900 70.535 154.750 76.410 ;
        RECT 159.730 76.070 165.580 81.925 ;
      LAYER pwell ;
        RECT 166.875 78.560 172.725 84.660 ;
      LAYER nwell ;
        RECT 173.350 76.600 177.110 81.875 ;
      LAYER pwell ;
        RECT 178.400 78.600 188.430 84.660 ;
        RECT 155.550 67.750 165.580 74.150 ;
      LAYER nwell ;
        RECT 166.875 70.540 170.635 75.850 ;
      LAYER pwell ;
        RECT 171.255 72.915 177.105 73.855 ;
        RECT 171.255 72.865 177.110 72.915 ;
        RECT 171.260 67.755 177.110 72.865 ;
      LAYER nwell ;
        RECT 178.400 70.535 184.250 76.410 ;
        RECT 189.230 76.070 195.080 81.925 ;
      LAYER pwell ;
        RECT 196.375 78.560 202.225 84.660 ;
      LAYER nwell ;
        RECT 202.850 76.600 206.610 81.875 ;
      LAYER pwell ;
        RECT 207.900 78.600 217.930 84.660 ;
        RECT 185.050 67.750 195.080 74.150 ;
      LAYER nwell ;
        RECT 196.375 70.540 200.135 75.850 ;
      LAYER pwell ;
        RECT 200.755 72.915 206.605 73.855 ;
        RECT 200.755 72.865 206.610 72.915 ;
        RECT 200.760 67.755 206.610 72.865 ;
      LAYER nwell ;
        RECT 207.900 70.535 213.750 76.410 ;
        RECT 218.730 76.070 224.580 81.925 ;
      LAYER pwell ;
        RECT 225.875 78.560 231.725 84.660 ;
      LAYER nwell ;
        RECT 232.350 76.600 236.110 81.875 ;
      LAYER pwell ;
        RECT 214.550 67.750 224.580 74.150 ;
      LAYER nwell ;
        RECT 225.875 70.540 229.635 75.850 ;
      LAYER pwell ;
        RECT 230.255 72.915 236.105 73.855 ;
        RECT 230.255 72.865 236.110 72.915 ;
        RECT 230.260 67.755 236.110 72.865 ;
      LAYER nwell ;
        RECT 243.100 66.570 249.890 73.570 ;
      LAYER pwell ;
        RECT 74.300 57.795 80.150 62.905 ;
        RECT 74.300 57.745 80.155 57.795 ;
        RECT 74.305 56.805 80.155 57.745 ;
      LAYER nwell ;
        RECT 80.775 54.810 84.535 60.120 ;
      LAYER pwell ;
        RECT 85.830 56.510 95.860 62.910 ;
      LAYER nwell ;
        RECT 74.300 48.785 78.060 54.060 ;
      LAYER pwell ;
        RECT 78.685 46.000 84.535 52.100 ;
      LAYER nwell ;
        RECT 85.830 48.735 91.680 54.590 ;
        RECT 96.660 54.250 102.510 60.125 ;
      LAYER pwell ;
        RECT 103.800 57.795 109.650 62.905 ;
        RECT 103.800 57.745 109.655 57.795 ;
        RECT 103.805 56.805 109.655 57.745 ;
      LAYER nwell ;
        RECT 110.275 54.810 114.035 60.120 ;
      LAYER pwell ;
        RECT 115.330 56.510 125.360 62.910 ;
        RECT 92.480 46.000 102.510 52.060 ;
      LAYER nwell ;
        RECT 103.800 48.785 107.560 54.060 ;
      LAYER pwell ;
        RECT 108.185 46.000 114.035 52.100 ;
      LAYER nwell ;
        RECT 115.330 48.735 121.180 54.590 ;
        RECT 126.160 54.250 132.010 60.125 ;
      LAYER pwell ;
        RECT 133.300 57.795 139.150 62.905 ;
        RECT 133.300 57.745 139.155 57.795 ;
        RECT 133.305 56.805 139.155 57.745 ;
      LAYER nwell ;
        RECT 139.775 54.810 143.535 60.120 ;
      LAYER pwell ;
        RECT 144.830 56.510 154.860 62.910 ;
        RECT 121.980 46.000 132.010 52.060 ;
      LAYER nwell ;
        RECT 133.300 48.785 137.060 54.060 ;
      LAYER pwell ;
        RECT 137.685 46.000 143.535 52.100 ;
      LAYER nwell ;
        RECT 144.830 48.735 150.680 54.590 ;
        RECT 155.660 54.250 161.510 60.125 ;
      LAYER pwell ;
        RECT 162.800 57.795 168.650 62.905 ;
        RECT 162.800 57.745 168.655 57.795 ;
        RECT 162.805 56.805 168.655 57.745 ;
      LAYER nwell ;
        RECT 169.275 54.810 173.035 60.120 ;
      LAYER pwell ;
        RECT 174.330 56.510 184.360 62.910 ;
        RECT 151.480 46.000 161.510 52.060 ;
      LAYER nwell ;
        RECT 162.800 48.785 166.560 54.060 ;
      LAYER pwell ;
        RECT 167.185 46.000 173.035 52.100 ;
      LAYER nwell ;
        RECT 174.330 48.735 180.180 54.590 ;
        RECT 185.160 54.250 191.010 60.125 ;
      LAYER pwell ;
        RECT 192.300 57.795 198.150 62.905 ;
        RECT 192.300 57.745 198.155 57.795 ;
        RECT 192.305 56.805 198.155 57.745 ;
      LAYER nwell ;
        RECT 198.775 54.810 202.535 60.120 ;
      LAYER pwell ;
        RECT 203.830 56.510 213.860 62.910 ;
        RECT 180.980 46.000 191.010 52.060 ;
      LAYER nwell ;
        RECT 192.300 48.785 196.060 54.060 ;
      LAYER pwell ;
        RECT 196.685 46.000 202.535 52.100 ;
      LAYER nwell ;
        RECT 203.830 48.735 209.680 54.590 ;
        RECT 214.660 54.250 220.510 60.125 ;
      LAYER pwell ;
        RECT 221.800 57.795 227.650 62.905 ;
        RECT 221.800 57.745 227.655 57.795 ;
        RECT 221.805 56.805 227.655 57.745 ;
      LAYER nwell ;
        RECT 228.275 54.810 232.035 60.120 ;
      LAYER pwell ;
        RECT 233.330 56.510 243.360 62.910 ;
        RECT 210.480 46.000 220.510 52.060 ;
      LAYER nwell ;
        RECT 221.800 48.785 225.560 54.060 ;
      LAYER pwell ;
        RECT 226.185 46.000 232.035 52.100 ;
      LAYER nwell ;
        RECT 233.330 48.735 239.180 54.590 ;
        RECT 244.160 54.250 250.010 60.125 ;
      LAYER pwell ;
        RECT 239.980 46.000 250.010 52.060 ;
      LAYER li1 ;
        RECT 90.080 84.480 92.425 84.610 ;
        RECT 93.490 84.480 96.350 84.610 ;
        RECT 97.405 84.480 99.750 84.610 ;
        RECT 90.080 84.310 99.750 84.480 ;
        RECT 90.080 84.130 92.425 84.310 ;
        RECT 93.490 84.130 96.350 84.310 ;
        RECT 97.405 84.130 99.750 84.310 ;
        RECT 90.080 79.480 90.250 84.130 ;
        RECT 90.590 79.535 90.880 84.130 ;
        RECT 90.650 79.290 90.820 79.535 ;
        RECT 90.800 77.080 91.930 78.080 ;
        RECT 92.680 77.770 92.970 83.830 ;
        RECT 94.770 79.535 95.060 84.130 ;
        RECT 94.830 79.290 95.000 79.535 ;
        RECT 96.860 77.870 97.150 83.830 ;
        RECT 98.950 79.535 99.240 84.130 ;
        RECT 99.010 79.525 99.205 79.535 ;
        RECT 99.010 79.290 99.180 79.525 ;
        RECT 99.580 79.380 99.750 84.130 ;
        RECT 108.055 84.470 110.400 84.610 ;
        RECT 111.200 84.470 113.545 84.610 ;
        RECT 108.055 84.300 113.545 84.470 ;
        RECT 108.055 84.130 110.400 84.300 ;
        RECT 111.200 84.130 113.545 84.300 ;
        RECT 100.910 81.745 103.255 81.890 ;
        RECT 104.055 81.745 106.400 81.890 ;
        RECT 100.910 81.575 106.400 81.745 ;
        RECT 100.910 81.410 103.255 81.575 ;
        RECT 104.055 81.410 106.400 81.575 ;
        RECT 96.860 77.770 97.680 77.870 ;
        RECT 92.680 77.270 97.680 77.770 ;
        RECT 90.080 71.010 90.250 75.865 ;
        RECT 90.590 71.010 90.880 75.860 ;
        RECT 92.680 71.320 92.970 77.270 ;
        RECT 100.910 76.750 101.080 81.410 ;
        RECT 101.420 76.580 101.710 81.410 ;
        RECT 105.600 76.580 105.890 81.410 ;
        RECT 106.230 76.810 106.400 81.410 ;
        RECT 108.055 79.775 108.225 84.130 ;
        RECT 108.565 79.780 108.855 84.130 ;
        RECT 112.745 79.780 113.035 84.130 ;
        RECT 113.375 79.775 113.545 84.130 ;
        RECT 119.580 84.480 121.925 84.610 ;
        RECT 122.990 84.480 125.850 84.610 ;
        RECT 126.905 84.480 129.250 84.610 ;
        RECT 119.580 84.310 129.250 84.480 ;
        RECT 119.580 84.130 121.925 84.310 ;
        RECT 122.990 84.130 125.850 84.310 ;
        RECT 126.905 84.130 129.250 84.310 ;
        RECT 115.835 81.860 117.930 81.890 ;
        RECT 115.680 81.695 117.930 81.860 ;
        RECT 114.530 81.525 117.930 81.695 ;
        RECT 114.530 78.550 114.700 81.525 ;
        RECT 115.680 81.440 117.930 81.525 ;
        RECT 115.835 81.410 117.930 81.440 ;
        RECT 108.800 77.870 110.000 78.180 ;
        RECT 115.035 77.965 115.330 81.040 ;
        RECT 108.300 77.250 110.000 77.870 ;
        RECT 108.800 77.050 110.000 77.250 ;
        RECT 114.805 77.185 115.545 77.965 ;
        RECT 94.770 71.010 95.060 75.860 ;
        RECT 95.400 71.010 95.570 75.865 ;
        RECT 90.080 70.885 92.425 71.010 ;
        RECT 93.225 70.980 95.570 71.010 ;
        RECT 93.225 70.885 95.750 70.980 ;
        RECT 90.080 70.715 95.750 70.885 ;
        RECT 90.080 70.530 92.425 70.715 ;
        RECT 93.225 70.560 95.750 70.715 ;
        RECT 93.225 70.530 95.570 70.560 ;
        RECT 96.730 68.290 96.900 73.030 ;
        RECT 97.300 72.885 97.470 73.120 ;
        RECT 97.275 72.875 97.470 72.885 ;
        RECT 101.480 72.875 101.650 73.100 ;
        RECT 105.660 72.875 105.830 73.100 ;
        RECT 97.240 68.290 97.530 72.875 ;
        RECT 101.420 68.290 101.710 72.875 ;
        RECT 105.600 68.290 105.890 72.875 ;
        RECT 106.230 68.290 106.400 72.930 ;
        RECT 108.055 71.010 108.225 74.935 ;
        RECT 108.565 71.010 108.855 75.080 ;
        RECT 108.055 70.980 110.150 71.010 ;
        RECT 108.055 70.890 110.305 70.980 ;
        RECT 111.285 70.890 111.455 74.925 ;
        RECT 108.055 70.720 111.455 70.890 ;
        RECT 108.055 70.560 110.305 70.720 ;
        RECT 108.055 70.530 110.150 70.560 ;
        RECT 96.730 68.100 99.075 68.290 ;
        RECT 100.130 68.100 102.990 68.290 ;
        RECT 104.055 68.100 106.400 68.290 ;
        RECT 96.730 67.930 106.400 68.100 ;
        RECT 96.730 67.810 99.075 67.930 ;
        RECT 100.130 67.810 102.990 67.930 ;
        RECT 104.055 67.810 106.400 67.930 ;
        RECT 112.440 68.290 112.610 72.640 ;
        RECT 112.950 68.290 113.240 72.635 ;
        RECT 115.035 68.595 115.330 77.185 ;
        RECT 117.130 77.000 117.420 81.410 ;
        RECT 117.760 76.995 117.930 81.410 ;
        RECT 119.580 79.480 119.750 84.130 ;
        RECT 120.090 79.535 120.380 84.130 ;
        RECT 120.150 79.290 120.320 79.535 ;
        RECT 120.300 77.080 121.430 78.080 ;
        RECT 122.180 77.770 122.470 83.830 ;
        RECT 124.270 79.535 124.560 84.130 ;
        RECT 124.330 79.290 124.500 79.535 ;
        RECT 126.360 77.870 126.650 83.830 ;
        RECT 128.450 79.535 128.740 84.130 ;
        RECT 128.510 79.525 128.705 79.535 ;
        RECT 128.510 79.290 128.680 79.525 ;
        RECT 129.080 79.380 129.250 84.130 ;
        RECT 137.555 84.470 139.900 84.610 ;
        RECT 140.700 84.470 143.045 84.610 ;
        RECT 137.555 84.300 143.045 84.470 ;
        RECT 137.555 84.130 139.900 84.300 ;
        RECT 140.700 84.130 143.045 84.300 ;
        RECT 130.410 81.745 132.755 81.890 ;
        RECT 133.555 81.745 135.900 81.890 ;
        RECT 130.410 81.575 135.900 81.745 ;
        RECT 130.410 81.410 132.755 81.575 ;
        RECT 133.555 81.410 135.900 81.575 ;
        RECT 126.360 77.770 127.180 77.870 ;
        RECT 122.180 77.270 127.180 77.770 ;
        RECT 117.130 68.290 117.420 72.635 ;
        RECT 117.760 68.290 117.930 72.640 ;
        RECT 119.580 71.010 119.750 75.865 ;
        RECT 120.090 71.010 120.380 75.860 ;
        RECT 122.180 71.320 122.470 77.270 ;
        RECT 130.410 76.750 130.580 81.410 ;
        RECT 130.920 76.580 131.210 81.410 ;
        RECT 135.100 76.580 135.390 81.410 ;
        RECT 135.730 76.810 135.900 81.410 ;
        RECT 137.555 79.775 137.725 84.130 ;
        RECT 138.065 79.780 138.355 84.130 ;
        RECT 142.245 79.780 142.535 84.130 ;
        RECT 142.875 79.775 143.045 84.130 ;
        RECT 149.080 84.480 151.425 84.610 ;
        RECT 152.490 84.480 155.350 84.610 ;
        RECT 156.405 84.480 158.750 84.610 ;
        RECT 149.080 84.310 158.750 84.480 ;
        RECT 149.080 84.130 151.425 84.310 ;
        RECT 152.490 84.130 155.350 84.310 ;
        RECT 156.405 84.130 158.750 84.310 ;
        RECT 145.335 81.860 147.430 81.890 ;
        RECT 145.180 81.695 147.430 81.860 ;
        RECT 144.030 81.525 147.430 81.695 ;
        RECT 144.030 78.550 144.200 81.525 ;
        RECT 145.180 81.440 147.430 81.525 ;
        RECT 145.335 81.410 147.430 81.440 ;
        RECT 138.300 77.870 139.500 78.180 ;
        RECT 144.535 77.965 144.830 81.040 ;
        RECT 137.800 77.250 139.500 77.870 ;
        RECT 138.300 77.050 139.500 77.250 ;
        RECT 144.305 77.185 145.045 77.965 ;
        RECT 124.270 71.010 124.560 75.860 ;
        RECT 124.900 71.010 125.070 75.865 ;
        RECT 119.580 70.885 121.925 71.010 ;
        RECT 122.725 70.980 125.070 71.010 ;
        RECT 122.725 70.885 125.250 70.980 ;
        RECT 119.580 70.715 125.250 70.885 ;
        RECT 119.580 70.530 121.925 70.715 ;
        RECT 122.725 70.560 125.250 70.715 ;
        RECT 122.725 70.530 125.070 70.560 ;
        RECT 112.440 68.115 114.785 68.290 ;
        RECT 115.585 68.115 117.930 68.290 ;
        RECT 112.440 67.945 117.930 68.115 ;
        RECT 112.440 67.810 114.785 67.945 ;
        RECT 115.585 67.810 117.930 67.945 ;
        RECT 126.230 68.290 126.400 73.030 ;
        RECT 126.800 72.885 126.970 73.120 ;
        RECT 126.775 72.875 126.970 72.885 ;
        RECT 130.980 72.875 131.150 73.100 ;
        RECT 135.160 72.875 135.330 73.100 ;
        RECT 126.740 68.290 127.030 72.875 ;
        RECT 130.920 68.290 131.210 72.875 ;
        RECT 135.100 68.290 135.390 72.875 ;
        RECT 135.730 68.290 135.900 72.930 ;
        RECT 137.555 71.010 137.725 74.935 ;
        RECT 138.065 71.010 138.355 75.080 ;
        RECT 137.555 70.980 139.650 71.010 ;
        RECT 137.555 70.890 139.805 70.980 ;
        RECT 140.785 70.890 140.955 74.925 ;
        RECT 137.555 70.720 140.955 70.890 ;
        RECT 137.555 70.560 139.805 70.720 ;
        RECT 137.555 70.530 139.650 70.560 ;
        RECT 126.230 68.100 128.575 68.290 ;
        RECT 129.630 68.100 132.490 68.290 ;
        RECT 133.555 68.100 135.900 68.290 ;
        RECT 126.230 67.930 135.900 68.100 ;
        RECT 126.230 67.810 128.575 67.930 ;
        RECT 129.630 67.810 132.490 67.930 ;
        RECT 133.555 67.810 135.900 67.930 ;
        RECT 141.940 68.290 142.110 72.640 ;
        RECT 142.450 68.290 142.740 72.635 ;
        RECT 144.535 68.595 144.830 77.185 ;
        RECT 146.630 77.000 146.920 81.410 ;
        RECT 147.260 76.995 147.430 81.410 ;
        RECT 149.080 79.480 149.250 84.130 ;
        RECT 149.590 79.535 149.880 84.130 ;
        RECT 149.650 79.290 149.820 79.535 ;
        RECT 149.800 77.080 150.930 78.080 ;
        RECT 151.680 77.770 151.970 83.830 ;
        RECT 153.770 79.535 154.060 84.130 ;
        RECT 153.830 79.290 154.000 79.535 ;
        RECT 155.860 77.870 156.150 83.830 ;
        RECT 157.950 79.535 158.240 84.130 ;
        RECT 158.010 79.525 158.205 79.535 ;
        RECT 158.010 79.290 158.180 79.525 ;
        RECT 158.580 79.380 158.750 84.130 ;
        RECT 167.055 84.470 169.400 84.610 ;
        RECT 170.200 84.470 172.545 84.610 ;
        RECT 167.055 84.300 172.545 84.470 ;
        RECT 167.055 84.130 169.400 84.300 ;
        RECT 170.200 84.130 172.545 84.300 ;
        RECT 159.910 81.745 162.255 81.890 ;
        RECT 163.055 81.745 165.400 81.890 ;
        RECT 159.910 81.575 165.400 81.745 ;
        RECT 159.910 81.410 162.255 81.575 ;
        RECT 163.055 81.410 165.400 81.575 ;
        RECT 155.860 77.770 156.680 77.870 ;
        RECT 151.680 77.270 156.680 77.770 ;
        RECT 146.630 68.290 146.920 72.635 ;
        RECT 147.260 68.290 147.430 72.640 ;
        RECT 149.080 71.010 149.250 75.865 ;
        RECT 149.590 71.010 149.880 75.860 ;
        RECT 151.680 71.320 151.970 77.270 ;
        RECT 159.910 76.750 160.080 81.410 ;
        RECT 160.420 76.580 160.710 81.410 ;
        RECT 164.600 76.580 164.890 81.410 ;
        RECT 165.230 76.810 165.400 81.410 ;
        RECT 167.055 79.775 167.225 84.130 ;
        RECT 167.565 79.780 167.855 84.130 ;
        RECT 171.745 79.780 172.035 84.130 ;
        RECT 172.375 79.775 172.545 84.130 ;
        RECT 178.580 84.480 180.925 84.610 ;
        RECT 181.990 84.480 184.850 84.610 ;
        RECT 185.905 84.480 188.250 84.610 ;
        RECT 178.580 84.310 188.250 84.480 ;
        RECT 178.580 84.130 180.925 84.310 ;
        RECT 181.990 84.130 184.850 84.310 ;
        RECT 185.905 84.130 188.250 84.310 ;
        RECT 174.835 81.860 176.930 81.890 ;
        RECT 174.680 81.695 176.930 81.860 ;
        RECT 173.530 81.525 176.930 81.695 ;
        RECT 173.530 78.550 173.700 81.525 ;
        RECT 174.680 81.440 176.930 81.525 ;
        RECT 174.835 81.410 176.930 81.440 ;
        RECT 167.800 77.870 169.000 78.180 ;
        RECT 174.035 77.965 174.330 81.040 ;
        RECT 167.300 77.250 169.000 77.870 ;
        RECT 167.800 77.050 169.000 77.250 ;
        RECT 173.805 77.185 174.545 77.965 ;
        RECT 153.770 71.010 154.060 75.860 ;
        RECT 154.400 71.010 154.570 75.865 ;
        RECT 149.080 70.885 151.425 71.010 ;
        RECT 152.225 70.980 154.570 71.010 ;
        RECT 152.225 70.885 154.750 70.980 ;
        RECT 149.080 70.715 154.750 70.885 ;
        RECT 149.080 70.530 151.425 70.715 ;
        RECT 152.225 70.560 154.750 70.715 ;
        RECT 152.225 70.530 154.570 70.560 ;
        RECT 141.940 68.115 144.285 68.290 ;
        RECT 145.085 68.115 147.430 68.290 ;
        RECT 141.940 67.945 147.430 68.115 ;
        RECT 141.940 67.810 144.285 67.945 ;
        RECT 145.085 67.810 147.430 67.945 ;
        RECT 155.730 68.290 155.900 73.030 ;
        RECT 156.300 72.885 156.470 73.120 ;
        RECT 156.275 72.875 156.470 72.885 ;
        RECT 160.480 72.875 160.650 73.100 ;
        RECT 164.660 72.875 164.830 73.100 ;
        RECT 156.240 68.290 156.530 72.875 ;
        RECT 160.420 68.290 160.710 72.875 ;
        RECT 164.600 68.290 164.890 72.875 ;
        RECT 165.230 68.290 165.400 72.930 ;
        RECT 167.055 71.010 167.225 74.935 ;
        RECT 167.565 71.010 167.855 75.080 ;
        RECT 167.055 70.980 169.150 71.010 ;
        RECT 167.055 70.890 169.305 70.980 ;
        RECT 170.285 70.890 170.455 74.925 ;
        RECT 167.055 70.720 170.455 70.890 ;
        RECT 167.055 70.560 169.305 70.720 ;
        RECT 167.055 70.530 169.150 70.560 ;
        RECT 155.730 68.100 158.075 68.290 ;
        RECT 159.130 68.100 161.990 68.290 ;
        RECT 163.055 68.100 165.400 68.290 ;
        RECT 155.730 67.930 165.400 68.100 ;
        RECT 155.730 67.810 158.075 67.930 ;
        RECT 159.130 67.810 161.990 67.930 ;
        RECT 163.055 67.810 165.400 67.930 ;
        RECT 171.440 68.290 171.610 72.640 ;
        RECT 171.950 68.290 172.240 72.635 ;
        RECT 174.035 68.595 174.330 77.185 ;
        RECT 176.130 77.000 176.420 81.410 ;
        RECT 176.760 76.995 176.930 81.410 ;
        RECT 178.580 79.480 178.750 84.130 ;
        RECT 179.090 79.535 179.380 84.130 ;
        RECT 179.150 79.290 179.320 79.535 ;
        RECT 179.300 77.080 180.430 78.080 ;
        RECT 181.180 77.770 181.470 83.830 ;
        RECT 183.270 79.535 183.560 84.130 ;
        RECT 183.330 79.290 183.500 79.535 ;
        RECT 185.360 77.870 185.650 83.830 ;
        RECT 187.450 79.535 187.740 84.130 ;
        RECT 187.510 79.525 187.705 79.535 ;
        RECT 187.510 79.290 187.680 79.525 ;
        RECT 188.080 79.380 188.250 84.130 ;
        RECT 196.555 84.470 198.900 84.610 ;
        RECT 199.700 84.470 202.045 84.610 ;
        RECT 196.555 84.300 202.045 84.470 ;
        RECT 196.555 84.130 198.900 84.300 ;
        RECT 199.700 84.130 202.045 84.300 ;
        RECT 189.410 81.745 191.755 81.890 ;
        RECT 192.555 81.745 194.900 81.890 ;
        RECT 189.410 81.575 194.900 81.745 ;
        RECT 189.410 81.410 191.755 81.575 ;
        RECT 192.555 81.410 194.900 81.575 ;
        RECT 185.360 77.770 186.180 77.870 ;
        RECT 181.180 77.270 186.180 77.770 ;
        RECT 176.130 68.290 176.420 72.635 ;
        RECT 176.760 68.290 176.930 72.640 ;
        RECT 178.580 71.010 178.750 75.865 ;
        RECT 179.090 71.010 179.380 75.860 ;
        RECT 181.180 71.320 181.470 77.270 ;
        RECT 189.410 76.750 189.580 81.410 ;
        RECT 189.920 76.580 190.210 81.410 ;
        RECT 194.100 76.580 194.390 81.410 ;
        RECT 194.730 76.810 194.900 81.410 ;
        RECT 196.555 79.775 196.725 84.130 ;
        RECT 197.065 79.780 197.355 84.130 ;
        RECT 201.245 79.780 201.535 84.130 ;
        RECT 201.875 79.775 202.045 84.130 ;
        RECT 208.080 84.480 210.425 84.610 ;
        RECT 211.490 84.480 214.350 84.610 ;
        RECT 215.405 84.480 217.750 84.610 ;
        RECT 208.080 84.310 217.750 84.480 ;
        RECT 208.080 84.130 210.425 84.310 ;
        RECT 211.490 84.130 214.350 84.310 ;
        RECT 215.405 84.130 217.750 84.310 ;
        RECT 204.335 81.860 206.430 81.890 ;
        RECT 204.180 81.695 206.430 81.860 ;
        RECT 203.030 81.525 206.430 81.695 ;
        RECT 203.030 78.550 203.200 81.525 ;
        RECT 204.180 81.440 206.430 81.525 ;
        RECT 204.335 81.410 206.430 81.440 ;
        RECT 197.300 77.870 198.500 78.180 ;
        RECT 203.535 77.965 203.830 81.040 ;
        RECT 196.800 77.250 198.500 77.870 ;
        RECT 197.300 77.050 198.500 77.250 ;
        RECT 203.305 77.185 204.045 77.965 ;
        RECT 183.270 71.010 183.560 75.860 ;
        RECT 183.900 71.010 184.070 75.865 ;
        RECT 178.580 70.885 180.925 71.010 ;
        RECT 181.725 70.980 184.070 71.010 ;
        RECT 181.725 70.885 184.250 70.980 ;
        RECT 178.580 70.715 184.250 70.885 ;
        RECT 178.580 70.530 180.925 70.715 ;
        RECT 181.725 70.560 184.250 70.715 ;
        RECT 181.725 70.530 184.070 70.560 ;
        RECT 171.440 68.115 173.785 68.290 ;
        RECT 174.585 68.115 176.930 68.290 ;
        RECT 171.440 67.945 176.930 68.115 ;
        RECT 171.440 67.810 173.785 67.945 ;
        RECT 174.585 67.810 176.930 67.945 ;
        RECT 185.230 68.290 185.400 73.030 ;
        RECT 185.800 72.885 185.970 73.120 ;
        RECT 185.775 72.875 185.970 72.885 ;
        RECT 189.980 72.875 190.150 73.100 ;
        RECT 194.160 72.875 194.330 73.100 ;
        RECT 185.740 68.290 186.030 72.875 ;
        RECT 189.920 68.290 190.210 72.875 ;
        RECT 194.100 68.290 194.390 72.875 ;
        RECT 194.730 68.290 194.900 72.930 ;
        RECT 196.555 71.010 196.725 74.935 ;
        RECT 197.065 71.010 197.355 75.080 ;
        RECT 196.555 70.980 198.650 71.010 ;
        RECT 196.555 70.890 198.805 70.980 ;
        RECT 199.785 70.890 199.955 74.925 ;
        RECT 196.555 70.720 199.955 70.890 ;
        RECT 196.555 70.560 198.805 70.720 ;
        RECT 196.555 70.530 198.650 70.560 ;
        RECT 185.230 68.100 187.575 68.290 ;
        RECT 188.630 68.100 191.490 68.290 ;
        RECT 192.555 68.100 194.900 68.290 ;
        RECT 185.230 67.930 194.900 68.100 ;
        RECT 185.230 67.810 187.575 67.930 ;
        RECT 188.630 67.810 191.490 67.930 ;
        RECT 192.555 67.810 194.900 67.930 ;
        RECT 200.940 68.290 201.110 72.640 ;
        RECT 201.450 68.290 201.740 72.635 ;
        RECT 203.535 68.595 203.830 77.185 ;
        RECT 205.630 77.000 205.920 81.410 ;
        RECT 206.260 76.995 206.430 81.410 ;
        RECT 208.080 79.480 208.250 84.130 ;
        RECT 208.590 79.535 208.880 84.130 ;
        RECT 208.650 79.290 208.820 79.535 ;
        RECT 208.800 77.080 209.930 78.080 ;
        RECT 210.680 77.770 210.970 83.830 ;
        RECT 212.770 79.535 213.060 84.130 ;
        RECT 212.830 79.290 213.000 79.535 ;
        RECT 214.860 77.870 215.150 83.830 ;
        RECT 216.950 79.535 217.240 84.130 ;
        RECT 217.010 79.525 217.205 79.535 ;
        RECT 217.010 79.290 217.180 79.525 ;
        RECT 217.580 79.380 217.750 84.130 ;
        RECT 226.055 84.470 228.400 84.610 ;
        RECT 229.200 84.470 231.545 84.610 ;
        RECT 226.055 84.300 231.545 84.470 ;
        RECT 226.055 84.130 228.400 84.300 ;
        RECT 229.200 84.130 231.545 84.300 ;
        RECT 218.910 81.745 221.255 81.890 ;
        RECT 222.055 81.745 224.400 81.890 ;
        RECT 218.910 81.575 224.400 81.745 ;
        RECT 218.910 81.410 221.255 81.575 ;
        RECT 222.055 81.410 224.400 81.575 ;
        RECT 214.860 77.770 215.680 77.870 ;
        RECT 210.680 77.270 215.680 77.770 ;
        RECT 205.630 68.290 205.920 72.635 ;
        RECT 206.260 68.290 206.430 72.640 ;
        RECT 208.080 71.010 208.250 75.865 ;
        RECT 208.590 71.010 208.880 75.860 ;
        RECT 210.680 71.320 210.970 77.270 ;
        RECT 218.910 76.750 219.080 81.410 ;
        RECT 219.420 76.580 219.710 81.410 ;
        RECT 223.600 76.580 223.890 81.410 ;
        RECT 224.230 76.810 224.400 81.410 ;
        RECT 226.055 79.775 226.225 84.130 ;
        RECT 226.565 79.780 226.855 84.130 ;
        RECT 230.745 79.780 231.035 84.130 ;
        RECT 231.375 79.775 231.545 84.130 ;
        RECT 233.835 81.860 235.930 81.890 ;
        RECT 233.680 81.695 235.930 81.860 ;
        RECT 232.530 81.525 235.930 81.695 ;
        RECT 232.530 78.550 232.700 81.525 ;
        RECT 233.680 81.440 235.930 81.525 ;
        RECT 233.835 81.410 235.930 81.440 ;
        RECT 226.800 77.870 228.000 78.180 ;
        RECT 233.035 77.965 233.330 81.040 ;
        RECT 226.300 77.250 228.000 77.870 ;
        RECT 226.800 77.050 228.000 77.250 ;
        RECT 232.805 77.185 233.545 77.965 ;
        RECT 212.770 71.010 213.060 75.860 ;
        RECT 213.400 71.010 213.570 75.865 ;
        RECT 208.080 70.885 210.425 71.010 ;
        RECT 211.225 70.980 213.570 71.010 ;
        RECT 211.225 70.885 213.750 70.980 ;
        RECT 208.080 70.715 213.750 70.885 ;
        RECT 208.080 70.530 210.425 70.715 ;
        RECT 211.225 70.560 213.750 70.715 ;
        RECT 211.225 70.530 213.570 70.560 ;
        RECT 200.940 68.115 203.285 68.290 ;
        RECT 204.085 68.115 206.430 68.290 ;
        RECT 200.940 67.945 206.430 68.115 ;
        RECT 200.940 67.810 203.285 67.945 ;
        RECT 204.085 67.810 206.430 67.945 ;
        RECT 214.730 68.290 214.900 73.030 ;
        RECT 215.300 72.885 215.470 73.120 ;
        RECT 215.275 72.875 215.470 72.885 ;
        RECT 219.480 72.875 219.650 73.100 ;
        RECT 223.660 72.875 223.830 73.100 ;
        RECT 215.240 68.290 215.530 72.875 ;
        RECT 219.420 68.290 219.710 72.875 ;
        RECT 223.600 68.290 223.890 72.875 ;
        RECT 224.230 68.290 224.400 72.930 ;
        RECT 226.055 71.010 226.225 74.935 ;
        RECT 226.565 71.010 226.855 75.080 ;
        RECT 226.055 70.980 228.150 71.010 ;
        RECT 226.055 70.890 228.305 70.980 ;
        RECT 229.285 70.890 229.455 74.925 ;
        RECT 226.055 70.720 229.455 70.890 ;
        RECT 226.055 70.560 228.305 70.720 ;
        RECT 226.055 70.530 228.150 70.560 ;
        RECT 214.730 68.100 217.075 68.290 ;
        RECT 218.130 68.100 220.990 68.290 ;
        RECT 222.055 68.100 224.400 68.290 ;
        RECT 214.730 67.930 224.400 68.100 ;
        RECT 214.730 67.810 217.075 67.930 ;
        RECT 218.130 67.810 220.990 67.930 ;
        RECT 222.055 67.810 224.400 67.930 ;
        RECT 230.440 68.290 230.610 72.640 ;
        RECT 230.950 68.290 231.240 72.635 ;
        RECT 233.035 68.595 233.330 77.185 ;
        RECT 235.130 77.000 235.420 81.410 ;
        RECT 235.760 76.995 235.930 81.410 ;
        RECT 243.280 73.220 246.580 73.390 ;
        RECT 235.130 68.290 235.420 72.635 ;
        RECT 235.760 68.290 235.930 72.640 ;
        RECT 230.440 68.115 232.785 68.290 ;
        RECT 233.585 68.115 235.930 68.290 ;
        RECT 230.440 67.945 235.930 68.115 ;
        RECT 230.440 67.810 232.785 67.945 ;
        RECT 233.585 67.810 235.930 67.945 ;
        RECT 243.280 67.380 243.450 73.220 ;
        RECT 246.410 72.930 246.580 73.220 ;
        RECT 246.410 72.760 249.710 72.930 ;
        RECT 243.930 72.490 245.930 72.660 ;
        RECT 244.010 72.460 245.850 72.490 ;
        RECT 244.010 68.110 245.850 68.140 ;
        RECT 243.930 67.940 245.930 68.110 ;
        RECT 246.410 67.380 246.580 72.760 ;
        RECT 247.140 67.650 248.980 67.680 ;
        RECT 247.060 67.480 249.060 67.650 ;
        RECT 243.280 67.210 246.580 67.380 ;
        RECT 246.410 66.920 246.580 67.210 ;
        RECT 249.540 66.920 249.710 72.760 ;
        RECT 246.410 66.750 249.710 66.920 ;
        RECT 74.480 62.715 76.825 62.850 ;
        RECT 77.625 62.715 79.970 62.850 ;
        RECT 74.480 62.545 79.970 62.715 ;
        RECT 74.480 62.370 76.825 62.545 ;
        RECT 77.625 62.370 79.970 62.545 ;
        RECT 74.480 58.020 74.650 62.370 ;
        RECT 74.990 58.025 75.280 62.370 ;
        RECT 74.480 49.250 74.650 53.665 ;
        RECT 74.990 49.250 75.280 53.660 ;
        RECT 77.080 53.475 77.375 62.065 ;
        RECT 79.170 58.025 79.460 62.370 ;
        RECT 79.800 58.020 79.970 62.370 ;
        RECT 86.010 62.730 88.355 62.850 ;
        RECT 89.420 62.730 92.280 62.850 ;
        RECT 93.335 62.730 95.680 62.850 ;
        RECT 86.010 62.560 95.680 62.730 ;
        RECT 86.010 62.370 88.355 62.560 ;
        RECT 89.420 62.370 92.280 62.560 ;
        RECT 93.335 62.370 95.680 62.560 ;
        RECT 82.260 60.100 84.355 60.130 ;
        RECT 82.105 59.940 84.355 60.100 ;
        RECT 80.955 59.770 84.355 59.940 ;
        RECT 80.955 55.735 81.125 59.770 ;
        RECT 82.105 59.680 84.355 59.770 ;
        RECT 82.260 59.650 84.355 59.680 ;
        RECT 83.555 55.580 83.845 59.650 ;
        RECT 84.185 55.725 84.355 59.650 ;
        RECT 86.010 57.730 86.180 62.370 ;
        RECT 86.520 57.785 86.810 62.370 ;
        RECT 90.700 57.785 90.990 62.370 ;
        RECT 94.880 57.785 95.170 62.370 ;
        RECT 86.580 57.560 86.750 57.785 ;
        RECT 90.760 57.560 90.930 57.785 ;
        RECT 94.940 57.775 95.135 57.785 ;
        RECT 94.940 57.540 95.110 57.775 ;
        RECT 95.510 57.630 95.680 62.370 ;
        RECT 103.980 62.715 106.325 62.850 ;
        RECT 107.125 62.715 109.470 62.850 ;
        RECT 103.980 62.545 109.470 62.715 ;
        RECT 103.980 62.370 106.325 62.545 ;
        RECT 107.125 62.370 109.470 62.545 ;
        RECT 96.840 60.100 99.185 60.130 ;
        RECT 96.660 59.945 99.185 60.100 ;
        RECT 99.985 59.945 102.330 60.130 ;
        RECT 96.660 59.775 102.330 59.945 ;
        RECT 96.660 59.680 99.185 59.775 ;
        RECT 96.840 59.650 99.185 59.680 ;
        RECT 99.985 59.650 102.330 59.775 ;
        RECT 96.840 54.795 97.010 59.650 ;
        RECT 97.350 54.800 97.640 59.650 ;
        RECT 76.865 52.695 77.605 53.475 ;
        RECT 82.410 53.410 83.610 53.610 ;
        RECT 82.410 52.790 84.110 53.410 ;
        RECT 77.080 49.620 77.375 52.695 ;
        RECT 82.410 52.480 83.610 52.790 ;
        RECT 74.480 49.220 76.575 49.250 ;
        RECT 74.480 49.135 76.730 49.220 ;
        RECT 77.710 49.135 77.880 52.110 ;
        RECT 74.480 48.965 77.880 49.135 ;
        RECT 74.480 48.800 76.730 48.965 ;
        RECT 74.480 48.770 76.575 48.800 ;
        RECT 78.865 46.530 79.035 50.885 ;
        RECT 79.375 46.530 79.665 50.880 ;
        RECT 83.555 46.530 83.845 50.880 ;
        RECT 84.185 46.530 84.355 50.885 ;
        RECT 86.010 49.250 86.180 53.850 ;
        RECT 86.520 49.250 86.810 54.080 ;
        RECT 90.700 49.250 90.990 54.080 ;
        RECT 91.330 49.250 91.500 53.910 ;
        RECT 99.440 53.390 99.730 59.340 ;
        RECT 101.530 54.800 101.820 59.650 ;
        RECT 102.160 54.795 102.330 59.650 ;
        RECT 103.980 58.020 104.150 62.370 ;
        RECT 104.490 58.025 104.780 62.370 ;
        RECT 94.730 52.890 99.730 53.390 ;
        RECT 94.730 52.790 95.550 52.890 ;
        RECT 86.010 49.085 88.355 49.250 ;
        RECT 89.155 49.085 91.500 49.250 ;
        RECT 86.010 48.915 91.500 49.085 ;
        RECT 86.010 48.770 88.355 48.915 ;
        RECT 89.155 48.770 91.500 48.915 ;
        RECT 78.865 46.360 81.210 46.530 ;
        RECT 82.010 46.360 84.355 46.530 ;
        RECT 78.865 46.190 84.355 46.360 ;
        RECT 78.865 46.050 81.210 46.190 ;
        RECT 82.010 46.050 84.355 46.190 ;
        RECT 92.660 46.530 92.830 51.280 ;
        RECT 93.230 51.135 93.400 51.370 ;
        RECT 93.205 51.125 93.400 51.135 ;
        RECT 93.170 46.530 93.460 51.125 ;
        RECT 95.260 46.830 95.550 52.790 ;
        RECT 97.410 51.125 97.580 51.370 ;
        RECT 97.350 46.530 97.640 51.125 ;
        RECT 99.440 46.830 99.730 52.890 ;
        RECT 100.480 52.580 101.610 53.580 ;
        RECT 101.590 51.125 101.760 51.370 ;
        RECT 101.530 46.530 101.820 51.125 ;
        RECT 102.160 46.530 102.330 51.180 ;
        RECT 103.980 49.250 104.150 53.665 ;
        RECT 104.490 49.250 104.780 53.660 ;
        RECT 106.580 53.475 106.875 62.065 ;
        RECT 108.670 58.025 108.960 62.370 ;
        RECT 109.300 58.020 109.470 62.370 ;
        RECT 115.510 62.730 117.855 62.850 ;
        RECT 118.920 62.730 121.780 62.850 ;
        RECT 122.835 62.730 125.180 62.850 ;
        RECT 115.510 62.560 125.180 62.730 ;
        RECT 115.510 62.370 117.855 62.560 ;
        RECT 118.920 62.370 121.780 62.560 ;
        RECT 122.835 62.370 125.180 62.560 ;
        RECT 111.760 60.100 113.855 60.130 ;
        RECT 111.605 59.940 113.855 60.100 ;
        RECT 110.455 59.770 113.855 59.940 ;
        RECT 110.455 55.735 110.625 59.770 ;
        RECT 111.605 59.680 113.855 59.770 ;
        RECT 111.760 59.650 113.855 59.680 ;
        RECT 113.055 55.580 113.345 59.650 ;
        RECT 113.685 55.725 113.855 59.650 ;
        RECT 115.510 57.730 115.680 62.370 ;
        RECT 116.020 57.785 116.310 62.370 ;
        RECT 120.200 57.785 120.490 62.370 ;
        RECT 124.380 57.785 124.670 62.370 ;
        RECT 116.080 57.560 116.250 57.785 ;
        RECT 120.260 57.560 120.430 57.785 ;
        RECT 124.440 57.775 124.635 57.785 ;
        RECT 124.440 57.540 124.610 57.775 ;
        RECT 125.010 57.630 125.180 62.370 ;
        RECT 133.480 62.715 135.825 62.850 ;
        RECT 136.625 62.715 138.970 62.850 ;
        RECT 133.480 62.545 138.970 62.715 ;
        RECT 133.480 62.370 135.825 62.545 ;
        RECT 136.625 62.370 138.970 62.545 ;
        RECT 126.340 60.100 128.685 60.130 ;
        RECT 126.160 59.945 128.685 60.100 ;
        RECT 129.485 59.945 131.830 60.130 ;
        RECT 126.160 59.775 131.830 59.945 ;
        RECT 126.160 59.680 128.685 59.775 ;
        RECT 126.340 59.650 128.685 59.680 ;
        RECT 129.485 59.650 131.830 59.775 ;
        RECT 126.340 54.795 126.510 59.650 ;
        RECT 126.850 54.800 127.140 59.650 ;
        RECT 106.365 52.695 107.105 53.475 ;
        RECT 111.910 53.410 113.110 53.610 ;
        RECT 111.910 52.790 113.610 53.410 ;
        RECT 106.580 49.620 106.875 52.695 ;
        RECT 111.910 52.480 113.110 52.790 ;
        RECT 103.980 49.220 106.075 49.250 ;
        RECT 103.980 49.135 106.230 49.220 ;
        RECT 107.210 49.135 107.380 52.110 ;
        RECT 103.980 48.965 107.380 49.135 ;
        RECT 103.980 48.800 106.230 48.965 ;
        RECT 103.980 48.770 106.075 48.800 ;
        RECT 92.660 46.350 95.005 46.530 ;
        RECT 96.060 46.350 98.920 46.530 ;
        RECT 99.985 46.350 102.330 46.530 ;
        RECT 92.660 46.180 102.330 46.350 ;
        RECT 92.660 46.050 95.005 46.180 ;
        RECT 96.060 46.050 98.920 46.180 ;
        RECT 99.985 46.050 102.330 46.180 ;
        RECT 108.365 46.530 108.535 50.885 ;
        RECT 108.875 46.530 109.165 50.880 ;
        RECT 113.055 46.530 113.345 50.880 ;
        RECT 113.685 46.530 113.855 50.885 ;
        RECT 115.510 49.250 115.680 53.850 ;
        RECT 116.020 49.250 116.310 54.080 ;
        RECT 120.200 49.250 120.490 54.080 ;
        RECT 120.830 49.250 121.000 53.910 ;
        RECT 128.940 53.390 129.230 59.340 ;
        RECT 131.030 54.800 131.320 59.650 ;
        RECT 131.660 54.795 131.830 59.650 ;
        RECT 133.480 58.020 133.650 62.370 ;
        RECT 133.990 58.025 134.280 62.370 ;
        RECT 124.230 52.890 129.230 53.390 ;
        RECT 124.230 52.790 125.050 52.890 ;
        RECT 115.510 49.085 117.855 49.250 ;
        RECT 118.655 49.085 121.000 49.250 ;
        RECT 115.510 48.915 121.000 49.085 ;
        RECT 115.510 48.770 117.855 48.915 ;
        RECT 118.655 48.770 121.000 48.915 ;
        RECT 108.365 46.360 110.710 46.530 ;
        RECT 111.510 46.360 113.855 46.530 ;
        RECT 108.365 46.190 113.855 46.360 ;
        RECT 108.365 46.050 110.710 46.190 ;
        RECT 111.510 46.050 113.855 46.190 ;
        RECT 122.160 46.530 122.330 51.280 ;
        RECT 122.730 51.135 122.900 51.370 ;
        RECT 122.705 51.125 122.900 51.135 ;
        RECT 122.670 46.530 122.960 51.125 ;
        RECT 124.760 46.830 125.050 52.790 ;
        RECT 126.910 51.125 127.080 51.370 ;
        RECT 126.850 46.530 127.140 51.125 ;
        RECT 128.940 46.830 129.230 52.890 ;
        RECT 129.980 52.580 131.110 53.580 ;
        RECT 131.090 51.125 131.260 51.370 ;
        RECT 131.030 46.530 131.320 51.125 ;
        RECT 131.660 46.530 131.830 51.180 ;
        RECT 133.480 49.250 133.650 53.665 ;
        RECT 133.990 49.250 134.280 53.660 ;
        RECT 136.080 53.475 136.375 62.065 ;
        RECT 138.170 58.025 138.460 62.370 ;
        RECT 138.800 58.020 138.970 62.370 ;
        RECT 145.010 62.730 147.355 62.850 ;
        RECT 148.420 62.730 151.280 62.850 ;
        RECT 152.335 62.730 154.680 62.850 ;
        RECT 145.010 62.560 154.680 62.730 ;
        RECT 145.010 62.370 147.355 62.560 ;
        RECT 148.420 62.370 151.280 62.560 ;
        RECT 152.335 62.370 154.680 62.560 ;
        RECT 141.260 60.100 143.355 60.130 ;
        RECT 141.105 59.940 143.355 60.100 ;
        RECT 139.955 59.770 143.355 59.940 ;
        RECT 139.955 55.735 140.125 59.770 ;
        RECT 141.105 59.680 143.355 59.770 ;
        RECT 141.260 59.650 143.355 59.680 ;
        RECT 142.555 55.580 142.845 59.650 ;
        RECT 143.185 55.725 143.355 59.650 ;
        RECT 145.010 57.730 145.180 62.370 ;
        RECT 145.520 57.785 145.810 62.370 ;
        RECT 149.700 57.785 149.990 62.370 ;
        RECT 153.880 57.785 154.170 62.370 ;
        RECT 145.580 57.560 145.750 57.785 ;
        RECT 149.760 57.560 149.930 57.785 ;
        RECT 153.940 57.775 154.135 57.785 ;
        RECT 153.940 57.540 154.110 57.775 ;
        RECT 154.510 57.630 154.680 62.370 ;
        RECT 162.980 62.715 165.325 62.850 ;
        RECT 166.125 62.715 168.470 62.850 ;
        RECT 162.980 62.545 168.470 62.715 ;
        RECT 162.980 62.370 165.325 62.545 ;
        RECT 166.125 62.370 168.470 62.545 ;
        RECT 155.840 60.100 158.185 60.130 ;
        RECT 155.660 59.945 158.185 60.100 ;
        RECT 158.985 59.945 161.330 60.130 ;
        RECT 155.660 59.775 161.330 59.945 ;
        RECT 155.660 59.680 158.185 59.775 ;
        RECT 155.840 59.650 158.185 59.680 ;
        RECT 158.985 59.650 161.330 59.775 ;
        RECT 155.840 54.795 156.010 59.650 ;
        RECT 156.350 54.800 156.640 59.650 ;
        RECT 135.865 52.695 136.605 53.475 ;
        RECT 141.410 53.410 142.610 53.610 ;
        RECT 141.410 52.790 143.110 53.410 ;
        RECT 136.080 49.620 136.375 52.695 ;
        RECT 141.410 52.480 142.610 52.790 ;
        RECT 133.480 49.220 135.575 49.250 ;
        RECT 133.480 49.135 135.730 49.220 ;
        RECT 136.710 49.135 136.880 52.110 ;
        RECT 133.480 48.965 136.880 49.135 ;
        RECT 133.480 48.800 135.730 48.965 ;
        RECT 133.480 48.770 135.575 48.800 ;
        RECT 122.160 46.350 124.505 46.530 ;
        RECT 125.560 46.350 128.420 46.530 ;
        RECT 129.485 46.350 131.830 46.530 ;
        RECT 122.160 46.180 131.830 46.350 ;
        RECT 122.160 46.050 124.505 46.180 ;
        RECT 125.560 46.050 128.420 46.180 ;
        RECT 129.485 46.050 131.830 46.180 ;
        RECT 137.865 46.530 138.035 50.885 ;
        RECT 138.375 46.530 138.665 50.880 ;
        RECT 142.555 46.530 142.845 50.880 ;
        RECT 143.185 46.530 143.355 50.885 ;
        RECT 145.010 49.250 145.180 53.850 ;
        RECT 145.520 49.250 145.810 54.080 ;
        RECT 149.700 49.250 149.990 54.080 ;
        RECT 150.330 49.250 150.500 53.910 ;
        RECT 158.440 53.390 158.730 59.340 ;
        RECT 160.530 54.800 160.820 59.650 ;
        RECT 161.160 54.795 161.330 59.650 ;
        RECT 162.980 58.020 163.150 62.370 ;
        RECT 163.490 58.025 163.780 62.370 ;
        RECT 153.730 52.890 158.730 53.390 ;
        RECT 153.730 52.790 154.550 52.890 ;
        RECT 145.010 49.085 147.355 49.250 ;
        RECT 148.155 49.085 150.500 49.250 ;
        RECT 145.010 48.915 150.500 49.085 ;
        RECT 145.010 48.770 147.355 48.915 ;
        RECT 148.155 48.770 150.500 48.915 ;
        RECT 137.865 46.360 140.210 46.530 ;
        RECT 141.010 46.360 143.355 46.530 ;
        RECT 137.865 46.190 143.355 46.360 ;
        RECT 137.865 46.050 140.210 46.190 ;
        RECT 141.010 46.050 143.355 46.190 ;
        RECT 151.660 46.530 151.830 51.280 ;
        RECT 152.230 51.135 152.400 51.370 ;
        RECT 152.205 51.125 152.400 51.135 ;
        RECT 152.170 46.530 152.460 51.125 ;
        RECT 154.260 46.830 154.550 52.790 ;
        RECT 156.410 51.125 156.580 51.370 ;
        RECT 156.350 46.530 156.640 51.125 ;
        RECT 158.440 46.830 158.730 52.890 ;
        RECT 159.480 52.580 160.610 53.580 ;
        RECT 160.590 51.125 160.760 51.370 ;
        RECT 160.530 46.530 160.820 51.125 ;
        RECT 161.160 46.530 161.330 51.180 ;
        RECT 162.980 49.250 163.150 53.665 ;
        RECT 163.490 49.250 163.780 53.660 ;
        RECT 165.580 53.475 165.875 62.065 ;
        RECT 167.670 58.025 167.960 62.370 ;
        RECT 168.300 58.020 168.470 62.370 ;
        RECT 174.510 62.730 176.855 62.850 ;
        RECT 177.920 62.730 180.780 62.850 ;
        RECT 181.835 62.730 184.180 62.850 ;
        RECT 174.510 62.560 184.180 62.730 ;
        RECT 174.510 62.370 176.855 62.560 ;
        RECT 177.920 62.370 180.780 62.560 ;
        RECT 181.835 62.370 184.180 62.560 ;
        RECT 170.760 60.100 172.855 60.130 ;
        RECT 170.605 59.940 172.855 60.100 ;
        RECT 169.455 59.770 172.855 59.940 ;
        RECT 169.455 55.735 169.625 59.770 ;
        RECT 170.605 59.680 172.855 59.770 ;
        RECT 170.760 59.650 172.855 59.680 ;
        RECT 172.055 55.580 172.345 59.650 ;
        RECT 172.685 55.725 172.855 59.650 ;
        RECT 174.510 57.730 174.680 62.370 ;
        RECT 175.020 57.785 175.310 62.370 ;
        RECT 179.200 57.785 179.490 62.370 ;
        RECT 183.380 57.785 183.670 62.370 ;
        RECT 175.080 57.560 175.250 57.785 ;
        RECT 179.260 57.560 179.430 57.785 ;
        RECT 183.440 57.775 183.635 57.785 ;
        RECT 183.440 57.540 183.610 57.775 ;
        RECT 184.010 57.630 184.180 62.370 ;
        RECT 192.480 62.715 194.825 62.850 ;
        RECT 195.625 62.715 197.970 62.850 ;
        RECT 192.480 62.545 197.970 62.715 ;
        RECT 192.480 62.370 194.825 62.545 ;
        RECT 195.625 62.370 197.970 62.545 ;
        RECT 185.340 60.100 187.685 60.130 ;
        RECT 185.160 59.945 187.685 60.100 ;
        RECT 188.485 59.945 190.830 60.130 ;
        RECT 185.160 59.775 190.830 59.945 ;
        RECT 185.160 59.680 187.685 59.775 ;
        RECT 185.340 59.650 187.685 59.680 ;
        RECT 188.485 59.650 190.830 59.775 ;
        RECT 185.340 54.795 185.510 59.650 ;
        RECT 185.850 54.800 186.140 59.650 ;
        RECT 165.365 52.695 166.105 53.475 ;
        RECT 170.910 53.410 172.110 53.610 ;
        RECT 170.910 52.790 172.610 53.410 ;
        RECT 165.580 49.620 165.875 52.695 ;
        RECT 170.910 52.480 172.110 52.790 ;
        RECT 162.980 49.220 165.075 49.250 ;
        RECT 162.980 49.135 165.230 49.220 ;
        RECT 166.210 49.135 166.380 52.110 ;
        RECT 162.980 48.965 166.380 49.135 ;
        RECT 162.980 48.800 165.230 48.965 ;
        RECT 162.980 48.770 165.075 48.800 ;
        RECT 151.660 46.350 154.005 46.530 ;
        RECT 155.060 46.350 157.920 46.530 ;
        RECT 158.985 46.350 161.330 46.530 ;
        RECT 151.660 46.180 161.330 46.350 ;
        RECT 151.660 46.050 154.005 46.180 ;
        RECT 155.060 46.050 157.920 46.180 ;
        RECT 158.985 46.050 161.330 46.180 ;
        RECT 167.365 46.530 167.535 50.885 ;
        RECT 167.875 46.530 168.165 50.880 ;
        RECT 172.055 46.530 172.345 50.880 ;
        RECT 172.685 46.530 172.855 50.885 ;
        RECT 174.510 49.250 174.680 53.850 ;
        RECT 175.020 49.250 175.310 54.080 ;
        RECT 179.200 49.250 179.490 54.080 ;
        RECT 179.830 49.250 180.000 53.910 ;
        RECT 187.940 53.390 188.230 59.340 ;
        RECT 190.030 54.800 190.320 59.650 ;
        RECT 190.660 54.795 190.830 59.650 ;
        RECT 192.480 58.020 192.650 62.370 ;
        RECT 192.990 58.025 193.280 62.370 ;
        RECT 183.230 52.890 188.230 53.390 ;
        RECT 183.230 52.790 184.050 52.890 ;
        RECT 174.510 49.085 176.855 49.250 ;
        RECT 177.655 49.085 180.000 49.250 ;
        RECT 174.510 48.915 180.000 49.085 ;
        RECT 174.510 48.770 176.855 48.915 ;
        RECT 177.655 48.770 180.000 48.915 ;
        RECT 167.365 46.360 169.710 46.530 ;
        RECT 170.510 46.360 172.855 46.530 ;
        RECT 167.365 46.190 172.855 46.360 ;
        RECT 167.365 46.050 169.710 46.190 ;
        RECT 170.510 46.050 172.855 46.190 ;
        RECT 181.160 46.530 181.330 51.280 ;
        RECT 181.730 51.135 181.900 51.370 ;
        RECT 181.705 51.125 181.900 51.135 ;
        RECT 181.670 46.530 181.960 51.125 ;
        RECT 183.760 46.830 184.050 52.790 ;
        RECT 185.910 51.125 186.080 51.370 ;
        RECT 185.850 46.530 186.140 51.125 ;
        RECT 187.940 46.830 188.230 52.890 ;
        RECT 188.980 52.580 190.110 53.580 ;
        RECT 190.090 51.125 190.260 51.370 ;
        RECT 190.030 46.530 190.320 51.125 ;
        RECT 190.660 46.530 190.830 51.180 ;
        RECT 192.480 49.250 192.650 53.665 ;
        RECT 192.990 49.250 193.280 53.660 ;
        RECT 195.080 53.475 195.375 62.065 ;
        RECT 197.170 58.025 197.460 62.370 ;
        RECT 197.800 58.020 197.970 62.370 ;
        RECT 204.010 62.730 206.355 62.850 ;
        RECT 207.420 62.730 210.280 62.850 ;
        RECT 211.335 62.730 213.680 62.850 ;
        RECT 204.010 62.560 213.680 62.730 ;
        RECT 204.010 62.370 206.355 62.560 ;
        RECT 207.420 62.370 210.280 62.560 ;
        RECT 211.335 62.370 213.680 62.560 ;
        RECT 200.260 60.100 202.355 60.130 ;
        RECT 200.105 59.940 202.355 60.100 ;
        RECT 198.955 59.770 202.355 59.940 ;
        RECT 198.955 55.735 199.125 59.770 ;
        RECT 200.105 59.680 202.355 59.770 ;
        RECT 200.260 59.650 202.355 59.680 ;
        RECT 201.555 55.580 201.845 59.650 ;
        RECT 202.185 55.725 202.355 59.650 ;
        RECT 204.010 57.730 204.180 62.370 ;
        RECT 204.520 57.785 204.810 62.370 ;
        RECT 208.700 57.785 208.990 62.370 ;
        RECT 212.880 57.785 213.170 62.370 ;
        RECT 204.580 57.560 204.750 57.785 ;
        RECT 208.760 57.560 208.930 57.785 ;
        RECT 212.940 57.775 213.135 57.785 ;
        RECT 212.940 57.540 213.110 57.775 ;
        RECT 213.510 57.630 213.680 62.370 ;
        RECT 221.980 62.715 224.325 62.850 ;
        RECT 225.125 62.715 227.470 62.850 ;
        RECT 221.980 62.545 227.470 62.715 ;
        RECT 221.980 62.370 224.325 62.545 ;
        RECT 225.125 62.370 227.470 62.545 ;
        RECT 214.840 60.100 217.185 60.130 ;
        RECT 214.660 59.945 217.185 60.100 ;
        RECT 217.985 59.945 220.330 60.130 ;
        RECT 214.660 59.775 220.330 59.945 ;
        RECT 214.660 59.680 217.185 59.775 ;
        RECT 214.840 59.650 217.185 59.680 ;
        RECT 217.985 59.650 220.330 59.775 ;
        RECT 214.840 54.795 215.010 59.650 ;
        RECT 215.350 54.800 215.640 59.650 ;
        RECT 194.865 52.695 195.605 53.475 ;
        RECT 200.410 53.410 201.610 53.610 ;
        RECT 200.410 52.790 202.110 53.410 ;
        RECT 195.080 49.620 195.375 52.695 ;
        RECT 200.410 52.480 201.610 52.790 ;
        RECT 192.480 49.220 194.575 49.250 ;
        RECT 192.480 49.135 194.730 49.220 ;
        RECT 195.710 49.135 195.880 52.110 ;
        RECT 192.480 48.965 195.880 49.135 ;
        RECT 192.480 48.800 194.730 48.965 ;
        RECT 192.480 48.770 194.575 48.800 ;
        RECT 181.160 46.350 183.505 46.530 ;
        RECT 184.560 46.350 187.420 46.530 ;
        RECT 188.485 46.350 190.830 46.530 ;
        RECT 181.160 46.180 190.830 46.350 ;
        RECT 181.160 46.050 183.505 46.180 ;
        RECT 184.560 46.050 187.420 46.180 ;
        RECT 188.485 46.050 190.830 46.180 ;
        RECT 196.865 46.530 197.035 50.885 ;
        RECT 197.375 46.530 197.665 50.880 ;
        RECT 201.555 46.530 201.845 50.880 ;
        RECT 202.185 46.530 202.355 50.885 ;
        RECT 204.010 49.250 204.180 53.850 ;
        RECT 204.520 49.250 204.810 54.080 ;
        RECT 208.700 49.250 208.990 54.080 ;
        RECT 209.330 49.250 209.500 53.910 ;
        RECT 217.440 53.390 217.730 59.340 ;
        RECT 219.530 54.800 219.820 59.650 ;
        RECT 220.160 54.795 220.330 59.650 ;
        RECT 221.980 58.020 222.150 62.370 ;
        RECT 222.490 58.025 222.780 62.370 ;
        RECT 212.730 52.890 217.730 53.390 ;
        RECT 212.730 52.790 213.550 52.890 ;
        RECT 204.010 49.085 206.355 49.250 ;
        RECT 207.155 49.085 209.500 49.250 ;
        RECT 204.010 48.915 209.500 49.085 ;
        RECT 204.010 48.770 206.355 48.915 ;
        RECT 207.155 48.770 209.500 48.915 ;
        RECT 196.865 46.360 199.210 46.530 ;
        RECT 200.010 46.360 202.355 46.530 ;
        RECT 196.865 46.190 202.355 46.360 ;
        RECT 196.865 46.050 199.210 46.190 ;
        RECT 200.010 46.050 202.355 46.190 ;
        RECT 210.660 46.530 210.830 51.280 ;
        RECT 211.230 51.135 211.400 51.370 ;
        RECT 211.205 51.125 211.400 51.135 ;
        RECT 211.170 46.530 211.460 51.125 ;
        RECT 213.260 46.830 213.550 52.790 ;
        RECT 215.410 51.125 215.580 51.370 ;
        RECT 215.350 46.530 215.640 51.125 ;
        RECT 217.440 46.830 217.730 52.890 ;
        RECT 218.480 52.580 219.610 53.580 ;
        RECT 219.590 51.125 219.760 51.370 ;
        RECT 219.530 46.530 219.820 51.125 ;
        RECT 220.160 46.530 220.330 51.180 ;
        RECT 221.980 49.250 222.150 53.665 ;
        RECT 222.490 49.250 222.780 53.660 ;
        RECT 224.580 53.475 224.875 62.065 ;
        RECT 226.670 58.025 226.960 62.370 ;
        RECT 227.300 58.020 227.470 62.370 ;
        RECT 233.510 62.730 235.855 62.850 ;
        RECT 236.920 62.730 239.780 62.850 ;
        RECT 240.835 62.730 243.180 62.850 ;
        RECT 233.510 62.560 243.180 62.730 ;
        RECT 233.510 62.370 235.855 62.560 ;
        RECT 236.920 62.370 239.780 62.560 ;
        RECT 240.835 62.370 243.180 62.560 ;
        RECT 229.760 60.100 231.855 60.130 ;
        RECT 229.605 59.940 231.855 60.100 ;
        RECT 228.455 59.770 231.855 59.940 ;
        RECT 228.455 55.735 228.625 59.770 ;
        RECT 229.605 59.680 231.855 59.770 ;
        RECT 229.760 59.650 231.855 59.680 ;
        RECT 231.055 55.580 231.345 59.650 ;
        RECT 231.685 55.725 231.855 59.650 ;
        RECT 233.510 57.730 233.680 62.370 ;
        RECT 234.020 57.785 234.310 62.370 ;
        RECT 238.200 57.785 238.490 62.370 ;
        RECT 242.380 57.785 242.670 62.370 ;
        RECT 234.080 57.560 234.250 57.785 ;
        RECT 238.260 57.560 238.430 57.785 ;
        RECT 242.440 57.775 242.635 57.785 ;
        RECT 242.440 57.540 242.610 57.775 ;
        RECT 243.010 57.630 243.180 62.370 ;
        RECT 244.340 60.100 246.685 60.130 ;
        RECT 244.160 59.945 246.685 60.100 ;
        RECT 247.485 59.945 249.830 60.130 ;
        RECT 244.160 59.775 249.830 59.945 ;
        RECT 244.160 59.680 246.685 59.775 ;
        RECT 244.340 59.650 246.685 59.680 ;
        RECT 247.485 59.650 249.830 59.775 ;
        RECT 244.340 54.795 244.510 59.650 ;
        RECT 244.850 54.800 245.140 59.650 ;
        RECT 224.365 52.695 225.105 53.475 ;
        RECT 229.910 53.410 231.110 53.610 ;
        RECT 229.910 52.790 231.610 53.410 ;
        RECT 224.580 49.620 224.875 52.695 ;
        RECT 229.910 52.480 231.110 52.790 ;
        RECT 221.980 49.220 224.075 49.250 ;
        RECT 221.980 49.135 224.230 49.220 ;
        RECT 225.210 49.135 225.380 52.110 ;
        RECT 221.980 48.965 225.380 49.135 ;
        RECT 221.980 48.800 224.230 48.965 ;
        RECT 221.980 48.770 224.075 48.800 ;
        RECT 210.660 46.350 213.005 46.530 ;
        RECT 214.060 46.350 216.920 46.530 ;
        RECT 217.985 46.350 220.330 46.530 ;
        RECT 210.660 46.180 220.330 46.350 ;
        RECT 210.660 46.050 213.005 46.180 ;
        RECT 214.060 46.050 216.920 46.180 ;
        RECT 217.985 46.050 220.330 46.180 ;
        RECT 226.365 46.530 226.535 50.885 ;
        RECT 226.875 46.530 227.165 50.880 ;
        RECT 231.055 46.530 231.345 50.880 ;
        RECT 231.685 46.530 231.855 50.885 ;
        RECT 233.510 49.250 233.680 53.850 ;
        RECT 234.020 49.250 234.310 54.080 ;
        RECT 238.200 49.250 238.490 54.080 ;
        RECT 238.830 49.250 239.000 53.910 ;
        RECT 246.940 53.390 247.230 59.340 ;
        RECT 249.030 54.800 249.320 59.650 ;
        RECT 249.660 54.795 249.830 59.650 ;
        RECT 242.230 52.890 247.230 53.390 ;
        RECT 242.230 52.790 243.050 52.890 ;
        RECT 233.510 49.085 235.855 49.250 ;
        RECT 236.655 49.085 239.000 49.250 ;
        RECT 233.510 48.915 239.000 49.085 ;
        RECT 233.510 48.770 235.855 48.915 ;
        RECT 236.655 48.770 239.000 48.915 ;
        RECT 226.365 46.360 228.710 46.530 ;
        RECT 229.510 46.360 231.855 46.530 ;
        RECT 226.365 46.190 231.855 46.360 ;
        RECT 226.365 46.050 228.710 46.190 ;
        RECT 229.510 46.050 231.855 46.190 ;
        RECT 240.160 46.530 240.330 51.280 ;
        RECT 240.730 51.135 240.900 51.370 ;
        RECT 240.705 51.125 240.900 51.135 ;
        RECT 240.670 46.530 240.960 51.125 ;
        RECT 242.760 46.830 243.050 52.790 ;
        RECT 244.910 51.125 245.080 51.370 ;
        RECT 244.850 46.530 245.140 51.125 ;
        RECT 246.940 46.830 247.230 52.890 ;
        RECT 247.980 52.580 249.110 53.580 ;
        RECT 249.090 51.125 249.260 51.370 ;
        RECT 249.030 46.530 249.320 51.125 ;
        RECT 249.660 46.530 249.830 51.180 ;
        RECT 240.160 46.350 242.505 46.530 ;
        RECT 243.560 46.350 246.420 46.530 ;
        RECT 247.485 46.350 249.830 46.530 ;
        RECT 240.160 46.180 249.830 46.350 ;
        RECT 240.160 46.050 242.505 46.180 ;
        RECT 243.560 46.050 246.420 46.180 ;
        RECT 247.485 46.050 249.830 46.180 ;
      LAYER mcon ;
        RECT 90.080 84.160 90.595 84.580 ;
        RECT 90.785 84.160 91.205 84.580 ;
        RECT 91.395 84.160 91.815 84.580 ;
        RECT 92.005 84.160 92.425 84.580 ;
        RECT 93.490 84.160 93.910 84.580 ;
        RECT 94.100 84.160 94.520 84.580 ;
        RECT 94.710 84.160 95.130 84.580 ;
        RECT 95.320 84.160 95.740 84.580 ;
        RECT 95.930 84.160 96.350 84.580 ;
        RECT 97.405 84.160 97.825 84.580 ;
        RECT 98.015 84.160 98.435 84.580 ;
        RECT 98.625 84.160 99.045 84.580 ;
        RECT 99.235 84.160 99.750 84.580 ;
        RECT 90.830 77.110 91.840 78.050 ;
        RECT 108.055 84.160 108.475 84.580 ;
        RECT 108.665 84.160 109.085 84.580 ;
        RECT 109.275 84.160 109.695 84.580 ;
        RECT 109.885 84.160 110.400 84.580 ;
        RECT 111.200 84.160 111.715 84.580 ;
        RECT 111.905 84.160 112.325 84.580 ;
        RECT 112.515 84.160 112.935 84.580 ;
        RECT 113.125 84.160 113.545 84.580 ;
        RECT 100.910 81.440 101.425 81.860 ;
        RECT 101.615 81.440 102.035 81.860 ;
        RECT 102.225 81.440 102.645 81.860 ;
        RECT 102.835 81.440 103.255 81.860 ;
        RECT 104.055 81.440 104.475 81.860 ;
        RECT 104.665 81.440 105.085 81.860 ;
        RECT 105.275 81.440 105.695 81.860 ;
        RECT 105.885 81.440 106.400 81.860 ;
        RECT 96.860 77.270 97.680 77.870 ;
        RECT 119.580 84.160 120.095 84.580 ;
        RECT 120.285 84.160 120.705 84.580 ;
        RECT 120.895 84.160 121.315 84.580 ;
        RECT 121.505 84.160 121.925 84.580 ;
        RECT 122.990 84.160 123.410 84.580 ;
        RECT 123.600 84.160 124.020 84.580 ;
        RECT 124.210 84.160 124.630 84.580 ;
        RECT 124.820 84.160 125.240 84.580 ;
        RECT 125.430 84.160 125.850 84.580 ;
        RECT 126.905 84.160 127.325 84.580 ;
        RECT 127.515 84.160 127.935 84.580 ;
        RECT 128.125 84.160 128.545 84.580 ;
        RECT 128.735 84.160 129.250 84.580 ;
        RECT 116.290 81.440 116.710 81.860 ;
        RECT 116.900 81.440 117.320 81.860 ;
        RECT 117.510 81.440 117.930 81.860 ;
        RECT 108.330 77.280 108.780 77.870 ;
        RECT 108.970 77.280 110.000 77.870 ;
        RECT 114.865 77.215 115.485 77.935 ;
        RECT 90.080 70.560 90.595 70.980 ;
        RECT 90.785 70.560 91.205 70.980 ;
        RECT 91.395 70.560 91.815 70.980 ;
        RECT 92.005 70.560 92.425 70.980 ;
        RECT 93.405 70.560 93.825 70.980 ;
        RECT 94.015 70.560 94.435 70.980 ;
        RECT 94.625 70.560 95.045 70.980 ;
        RECT 95.235 70.560 95.750 70.980 ;
        RECT 108.665 70.560 109.085 70.980 ;
        RECT 109.275 70.560 109.695 70.980 ;
        RECT 109.885 70.560 110.305 70.980 ;
        RECT 96.730 67.840 97.245 68.260 ;
        RECT 97.435 67.840 97.855 68.260 ;
        RECT 98.045 67.840 98.465 68.260 ;
        RECT 98.655 67.840 99.075 68.260 ;
        RECT 100.130 67.840 100.550 68.260 ;
        RECT 100.740 67.840 101.160 68.260 ;
        RECT 101.350 67.840 101.770 68.260 ;
        RECT 101.960 67.840 102.380 68.260 ;
        RECT 102.570 67.840 102.990 68.260 ;
        RECT 104.055 67.840 104.475 68.260 ;
        RECT 104.665 67.840 105.085 68.260 ;
        RECT 105.275 67.840 105.695 68.260 ;
        RECT 105.885 67.840 106.400 68.260 ;
        RECT 120.330 77.110 121.340 78.050 ;
        RECT 137.555 84.160 137.975 84.580 ;
        RECT 138.165 84.160 138.585 84.580 ;
        RECT 138.775 84.160 139.195 84.580 ;
        RECT 139.385 84.160 139.900 84.580 ;
        RECT 140.700 84.160 141.215 84.580 ;
        RECT 141.405 84.160 141.825 84.580 ;
        RECT 142.015 84.160 142.435 84.580 ;
        RECT 142.625 84.160 143.045 84.580 ;
        RECT 130.410 81.440 130.925 81.860 ;
        RECT 131.115 81.440 131.535 81.860 ;
        RECT 131.725 81.440 132.145 81.860 ;
        RECT 132.335 81.440 132.755 81.860 ;
        RECT 133.555 81.440 133.975 81.860 ;
        RECT 134.165 81.440 134.585 81.860 ;
        RECT 134.775 81.440 135.195 81.860 ;
        RECT 135.385 81.440 135.900 81.860 ;
        RECT 126.360 77.270 127.180 77.870 ;
        RECT 149.080 84.160 149.595 84.580 ;
        RECT 149.785 84.160 150.205 84.580 ;
        RECT 150.395 84.160 150.815 84.580 ;
        RECT 151.005 84.160 151.425 84.580 ;
        RECT 152.490 84.160 152.910 84.580 ;
        RECT 153.100 84.160 153.520 84.580 ;
        RECT 153.710 84.160 154.130 84.580 ;
        RECT 154.320 84.160 154.740 84.580 ;
        RECT 154.930 84.160 155.350 84.580 ;
        RECT 156.405 84.160 156.825 84.580 ;
        RECT 157.015 84.160 157.435 84.580 ;
        RECT 157.625 84.160 158.045 84.580 ;
        RECT 158.235 84.160 158.750 84.580 ;
        RECT 145.790 81.440 146.210 81.860 ;
        RECT 146.400 81.440 146.820 81.860 ;
        RECT 147.010 81.440 147.430 81.860 ;
        RECT 137.830 77.280 138.280 77.870 ;
        RECT 138.470 77.280 139.500 77.870 ;
        RECT 144.365 77.215 144.985 77.935 ;
        RECT 119.580 70.560 120.095 70.980 ;
        RECT 120.285 70.560 120.705 70.980 ;
        RECT 120.895 70.560 121.315 70.980 ;
        RECT 121.505 70.560 121.925 70.980 ;
        RECT 122.905 70.560 123.325 70.980 ;
        RECT 123.515 70.560 123.935 70.980 ;
        RECT 124.125 70.560 124.545 70.980 ;
        RECT 124.735 70.560 125.250 70.980 ;
        RECT 112.440 67.840 112.955 68.260 ;
        RECT 113.145 67.840 113.565 68.260 ;
        RECT 113.755 67.840 114.175 68.260 ;
        RECT 114.365 67.840 114.785 68.260 ;
        RECT 115.585 67.840 116.005 68.260 ;
        RECT 116.195 67.840 116.615 68.260 ;
        RECT 116.805 67.840 117.225 68.260 ;
        RECT 117.415 67.840 117.930 68.260 ;
        RECT 138.165 70.560 138.585 70.980 ;
        RECT 138.775 70.560 139.195 70.980 ;
        RECT 139.385 70.560 139.805 70.980 ;
        RECT 126.230 67.840 126.745 68.260 ;
        RECT 126.935 67.840 127.355 68.260 ;
        RECT 127.545 67.840 127.965 68.260 ;
        RECT 128.155 67.840 128.575 68.260 ;
        RECT 129.630 67.840 130.050 68.260 ;
        RECT 130.240 67.840 130.660 68.260 ;
        RECT 130.850 67.840 131.270 68.260 ;
        RECT 131.460 67.840 131.880 68.260 ;
        RECT 132.070 67.840 132.490 68.260 ;
        RECT 133.555 67.840 133.975 68.260 ;
        RECT 134.165 67.840 134.585 68.260 ;
        RECT 134.775 67.840 135.195 68.260 ;
        RECT 135.385 67.840 135.900 68.260 ;
        RECT 149.830 77.110 150.840 78.050 ;
        RECT 167.055 84.160 167.475 84.580 ;
        RECT 167.665 84.160 168.085 84.580 ;
        RECT 168.275 84.160 168.695 84.580 ;
        RECT 168.885 84.160 169.400 84.580 ;
        RECT 170.200 84.160 170.715 84.580 ;
        RECT 170.905 84.160 171.325 84.580 ;
        RECT 171.515 84.160 171.935 84.580 ;
        RECT 172.125 84.160 172.545 84.580 ;
        RECT 159.910 81.440 160.425 81.860 ;
        RECT 160.615 81.440 161.035 81.860 ;
        RECT 161.225 81.440 161.645 81.860 ;
        RECT 161.835 81.440 162.255 81.860 ;
        RECT 163.055 81.440 163.475 81.860 ;
        RECT 163.665 81.440 164.085 81.860 ;
        RECT 164.275 81.440 164.695 81.860 ;
        RECT 164.885 81.440 165.400 81.860 ;
        RECT 155.860 77.270 156.680 77.870 ;
        RECT 178.580 84.160 179.095 84.580 ;
        RECT 179.285 84.160 179.705 84.580 ;
        RECT 179.895 84.160 180.315 84.580 ;
        RECT 180.505 84.160 180.925 84.580 ;
        RECT 181.990 84.160 182.410 84.580 ;
        RECT 182.600 84.160 183.020 84.580 ;
        RECT 183.210 84.160 183.630 84.580 ;
        RECT 183.820 84.160 184.240 84.580 ;
        RECT 184.430 84.160 184.850 84.580 ;
        RECT 185.905 84.160 186.325 84.580 ;
        RECT 186.515 84.160 186.935 84.580 ;
        RECT 187.125 84.160 187.545 84.580 ;
        RECT 187.735 84.160 188.250 84.580 ;
        RECT 175.290 81.440 175.710 81.860 ;
        RECT 175.900 81.440 176.320 81.860 ;
        RECT 176.510 81.440 176.930 81.860 ;
        RECT 167.330 77.280 167.780 77.870 ;
        RECT 167.970 77.280 169.000 77.870 ;
        RECT 173.865 77.215 174.485 77.935 ;
        RECT 149.080 70.560 149.595 70.980 ;
        RECT 149.785 70.560 150.205 70.980 ;
        RECT 150.395 70.560 150.815 70.980 ;
        RECT 151.005 70.560 151.425 70.980 ;
        RECT 152.405 70.560 152.825 70.980 ;
        RECT 153.015 70.560 153.435 70.980 ;
        RECT 153.625 70.560 154.045 70.980 ;
        RECT 154.235 70.560 154.750 70.980 ;
        RECT 141.940 67.840 142.455 68.260 ;
        RECT 142.645 67.840 143.065 68.260 ;
        RECT 143.255 67.840 143.675 68.260 ;
        RECT 143.865 67.840 144.285 68.260 ;
        RECT 145.085 67.840 145.505 68.260 ;
        RECT 145.695 67.840 146.115 68.260 ;
        RECT 146.305 67.840 146.725 68.260 ;
        RECT 146.915 67.840 147.430 68.260 ;
        RECT 167.665 70.560 168.085 70.980 ;
        RECT 168.275 70.560 168.695 70.980 ;
        RECT 168.885 70.560 169.305 70.980 ;
        RECT 155.730 67.840 156.245 68.260 ;
        RECT 156.435 67.840 156.855 68.260 ;
        RECT 157.045 67.840 157.465 68.260 ;
        RECT 157.655 67.840 158.075 68.260 ;
        RECT 159.130 67.840 159.550 68.260 ;
        RECT 159.740 67.840 160.160 68.260 ;
        RECT 160.350 67.840 160.770 68.260 ;
        RECT 160.960 67.840 161.380 68.260 ;
        RECT 161.570 67.840 161.990 68.260 ;
        RECT 163.055 67.840 163.475 68.260 ;
        RECT 163.665 67.840 164.085 68.260 ;
        RECT 164.275 67.840 164.695 68.260 ;
        RECT 164.885 67.840 165.400 68.260 ;
        RECT 179.330 77.110 180.340 78.050 ;
        RECT 196.555 84.160 196.975 84.580 ;
        RECT 197.165 84.160 197.585 84.580 ;
        RECT 197.775 84.160 198.195 84.580 ;
        RECT 198.385 84.160 198.900 84.580 ;
        RECT 199.700 84.160 200.215 84.580 ;
        RECT 200.405 84.160 200.825 84.580 ;
        RECT 201.015 84.160 201.435 84.580 ;
        RECT 201.625 84.160 202.045 84.580 ;
        RECT 189.410 81.440 189.925 81.860 ;
        RECT 190.115 81.440 190.535 81.860 ;
        RECT 190.725 81.440 191.145 81.860 ;
        RECT 191.335 81.440 191.755 81.860 ;
        RECT 192.555 81.440 192.975 81.860 ;
        RECT 193.165 81.440 193.585 81.860 ;
        RECT 193.775 81.440 194.195 81.860 ;
        RECT 194.385 81.440 194.900 81.860 ;
        RECT 185.360 77.270 186.180 77.870 ;
        RECT 208.080 84.160 208.595 84.580 ;
        RECT 208.785 84.160 209.205 84.580 ;
        RECT 209.395 84.160 209.815 84.580 ;
        RECT 210.005 84.160 210.425 84.580 ;
        RECT 211.490 84.160 211.910 84.580 ;
        RECT 212.100 84.160 212.520 84.580 ;
        RECT 212.710 84.160 213.130 84.580 ;
        RECT 213.320 84.160 213.740 84.580 ;
        RECT 213.930 84.160 214.350 84.580 ;
        RECT 215.405 84.160 215.825 84.580 ;
        RECT 216.015 84.160 216.435 84.580 ;
        RECT 216.625 84.160 217.045 84.580 ;
        RECT 217.235 84.160 217.750 84.580 ;
        RECT 204.790 81.440 205.210 81.860 ;
        RECT 205.400 81.440 205.820 81.860 ;
        RECT 206.010 81.440 206.430 81.860 ;
        RECT 196.830 77.280 197.280 77.870 ;
        RECT 197.470 77.280 198.500 77.870 ;
        RECT 203.365 77.215 203.985 77.935 ;
        RECT 178.580 70.560 179.095 70.980 ;
        RECT 179.285 70.560 179.705 70.980 ;
        RECT 179.895 70.560 180.315 70.980 ;
        RECT 180.505 70.560 180.925 70.980 ;
        RECT 181.905 70.560 182.325 70.980 ;
        RECT 182.515 70.560 182.935 70.980 ;
        RECT 183.125 70.560 183.545 70.980 ;
        RECT 183.735 70.560 184.250 70.980 ;
        RECT 171.440 67.840 171.955 68.260 ;
        RECT 172.145 67.840 172.565 68.260 ;
        RECT 172.755 67.840 173.175 68.260 ;
        RECT 173.365 67.840 173.785 68.260 ;
        RECT 174.585 67.840 175.005 68.260 ;
        RECT 175.195 67.840 175.615 68.260 ;
        RECT 175.805 67.840 176.225 68.260 ;
        RECT 176.415 67.840 176.930 68.260 ;
        RECT 197.165 70.560 197.585 70.980 ;
        RECT 197.775 70.560 198.195 70.980 ;
        RECT 198.385 70.560 198.805 70.980 ;
        RECT 185.230 67.840 185.745 68.260 ;
        RECT 185.935 67.840 186.355 68.260 ;
        RECT 186.545 67.840 186.965 68.260 ;
        RECT 187.155 67.840 187.575 68.260 ;
        RECT 188.630 67.840 189.050 68.260 ;
        RECT 189.240 67.840 189.660 68.260 ;
        RECT 189.850 67.840 190.270 68.260 ;
        RECT 190.460 67.840 190.880 68.260 ;
        RECT 191.070 67.840 191.490 68.260 ;
        RECT 192.555 67.840 192.975 68.260 ;
        RECT 193.165 67.840 193.585 68.260 ;
        RECT 193.775 67.840 194.195 68.260 ;
        RECT 194.385 67.840 194.900 68.260 ;
        RECT 208.830 77.110 209.840 78.050 ;
        RECT 226.055 84.160 226.475 84.580 ;
        RECT 226.665 84.160 227.085 84.580 ;
        RECT 227.275 84.160 227.695 84.580 ;
        RECT 227.885 84.160 228.400 84.580 ;
        RECT 229.200 84.160 229.715 84.580 ;
        RECT 229.905 84.160 230.325 84.580 ;
        RECT 230.515 84.160 230.935 84.580 ;
        RECT 231.125 84.160 231.545 84.580 ;
        RECT 218.910 81.440 219.425 81.860 ;
        RECT 219.615 81.440 220.035 81.860 ;
        RECT 220.225 81.440 220.645 81.860 ;
        RECT 220.835 81.440 221.255 81.860 ;
        RECT 222.055 81.440 222.475 81.860 ;
        RECT 222.665 81.440 223.085 81.860 ;
        RECT 223.275 81.440 223.695 81.860 ;
        RECT 223.885 81.440 224.400 81.860 ;
        RECT 214.860 77.270 215.680 77.870 ;
        RECT 234.290 81.440 234.710 81.860 ;
        RECT 234.900 81.440 235.320 81.860 ;
        RECT 235.510 81.440 235.930 81.860 ;
        RECT 226.330 77.280 226.780 77.870 ;
        RECT 226.970 77.280 228.000 77.870 ;
        RECT 232.865 77.215 233.485 77.935 ;
        RECT 208.080 70.560 208.595 70.980 ;
        RECT 208.785 70.560 209.205 70.980 ;
        RECT 209.395 70.560 209.815 70.980 ;
        RECT 210.005 70.560 210.425 70.980 ;
        RECT 211.405 70.560 211.825 70.980 ;
        RECT 212.015 70.560 212.435 70.980 ;
        RECT 212.625 70.560 213.045 70.980 ;
        RECT 213.235 70.560 213.750 70.980 ;
        RECT 200.940 67.840 201.455 68.260 ;
        RECT 201.645 67.840 202.065 68.260 ;
        RECT 202.255 67.840 202.675 68.260 ;
        RECT 202.865 67.840 203.285 68.260 ;
        RECT 204.085 67.840 204.505 68.260 ;
        RECT 204.695 67.840 205.115 68.260 ;
        RECT 205.305 67.840 205.725 68.260 ;
        RECT 205.915 67.840 206.430 68.260 ;
        RECT 226.665 70.560 227.085 70.980 ;
        RECT 227.275 70.560 227.695 70.980 ;
        RECT 227.885 70.560 228.305 70.980 ;
        RECT 214.730 67.840 215.245 68.260 ;
        RECT 215.435 67.840 215.855 68.260 ;
        RECT 216.045 67.840 216.465 68.260 ;
        RECT 216.655 67.840 217.075 68.260 ;
        RECT 218.130 67.840 218.550 68.260 ;
        RECT 218.740 67.840 219.160 68.260 ;
        RECT 219.350 67.840 219.770 68.260 ;
        RECT 219.960 67.840 220.380 68.260 ;
        RECT 220.570 67.840 220.990 68.260 ;
        RECT 222.055 67.840 222.475 68.260 ;
        RECT 222.665 67.840 223.085 68.260 ;
        RECT 223.275 67.840 223.695 68.260 ;
        RECT 223.885 67.840 224.400 68.260 ;
        RECT 230.440 67.840 230.955 68.260 ;
        RECT 231.145 67.840 231.565 68.260 ;
        RECT 231.755 67.840 232.175 68.260 ;
        RECT 232.365 67.840 232.785 68.260 ;
        RECT 233.585 67.840 234.005 68.260 ;
        RECT 234.195 67.840 234.615 68.260 ;
        RECT 234.805 67.840 235.225 68.260 ;
        RECT 235.415 67.840 235.930 68.260 ;
        RECT 244.010 67.940 245.850 68.140 ;
        RECT 247.140 67.480 248.980 67.680 ;
        RECT 74.480 62.400 74.995 62.820 ;
        RECT 75.185 62.400 75.605 62.820 ;
        RECT 75.795 62.400 76.215 62.820 ;
        RECT 76.405 62.400 76.825 62.820 ;
        RECT 77.625 62.400 78.045 62.820 ;
        RECT 78.235 62.400 78.655 62.820 ;
        RECT 78.845 62.400 79.265 62.820 ;
        RECT 79.455 62.400 79.970 62.820 ;
        RECT 86.010 62.400 86.525 62.820 ;
        RECT 86.715 62.400 87.135 62.820 ;
        RECT 87.325 62.400 87.745 62.820 ;
        RECT 87.935 62.400 88.355 62.820 ;
        RECT 89.420 62.400 89.840 62.820 ;
        RECT 90.030 62.400 90.450 62.820 ;
        RECT 90.640 62.400 91.060 62.820 ;
        RECT 91.250 62.400 91.670 62.820 ;
        RECT 91.860 62.400 92.280 62.820 ;
        RECT 93.335 62.400 93.755 62.820 ;
        RECT 93.945 62.400 94.365 62.820 ;
        RECT 94.555 62.400 94.975 62.820 ;
        RECT 95.165 62.400 95.680 62.820 ;
        RECT 82.715 59.680 83.135 60.100 ;
        RECT 83.325 59.680 83.745 60.100 ;
        RECT 83.935 59.680 84.355 60.100 ;
        RECT 103.980 62.400 104.495 62.820 ;
        RECT 104.685 62.400 105.105 62.820 ;
        RECT 105.295 62.400 105.715 62.820 ;
        RECT 105.905 62.400 106.325 62.820 ;
        RECT 107.125 62.400 107.545 62.820 ;
        RECT 107.735 62.400 108.155 62.820 ;
        RECT 108.345 62.400 108.765 62.820 ;
        RECT 108.955 62.400 109.470 62.820 ;
        RECT 97.365 59.680 97.785 60.100 ;
        RECT 97.975 59.680 98.395 60.100 ;
        RECT 98.585 59.680 99.005 60.100 ;
        RECT 99.985 59.680 100.405 60.100 ;
        RECT 100.595 59.680 101.015 60.100 ;
        RECT 101.205 59.680 101.625 60.100 ;
        RECT 101.815 59.680 102.330 60.100 ;
        RECT 76.925 52.725 77.545 53.445 ;
        RECT 82.410 52.790 83.440 53.380 ;
        RECT 83.630 52.790 84.080 53.380 ;
        RECT 75.090 48.800 75.510 49.220 ;
        RECT 75.700 48.800 76.120 49.220 ;
        RECT 76.310 48.800 76.730 49.220 ;
        RECT 86.010 48.800 86.525 49.220 ;
        RECT 86.715 48.800 87.135 49.220 ;
        RECT 87.325 48.800 87.745 49.220 ;
        RECT 87.935 48.800 88.355 49.220 ;
        RECT 89.155 48.800 89.575 49.220 ;
        RECT 89.765 48.800 90.185 49.220 ;
        RECT 90.375 48.800 90.795 49.220 ;
        RECT 90.985 48.800 91.500 49.220 ;
        RECT 78.865 46.080 79.285 46.500 ;
        RECT 79.475 46.080 79.895 46.500 ;
        RECT 80.085 46.080 80.505 46.500 ;
        RECT 80.695 46.080 81.210 46.500 ;
        RECT 82.010 46.080 82.525 46.500 ;
        RECT 82.715 46.080 83.135 46.500 ;
        RECT 83.325 46.080 83.745 46.500 ;
        RECT 83.935 46.080 84.355 46.500 ;
        RECT 100.570 52.610 101.580 53.550 ;
        RECT 115.510 62.400 116.025 62.820 ;
        RECT 116.215 62.400 116.635 62.820 ;
        RECT 116.825 62.400 117.245 62.820 ;
        RECT 117.435 62.400 117.855 62.820 ;
        RECT 118.920 62.400 119.340 62.820 ;
        RECT 119.530 62.400 119.950 62.820 ;
        RECT 120.140 62.400 120.560 62.820 ;
        RECT 120.750 62.400 121.170 62.820 ;
        RECT 121.360 62.400 121.780 62.820 ;
        RECT 122.835 62.400 123.255 62.820 ;
        RECT 123.445 62.400 123.865 62.820 ;
        RECT 124.055 62.400 124.475 62.820 ;
        RECT 124.665 62.400 125.180 62.820 ;
        RECT 112.215 59.680 112.635 60.100 ;
        RECT 112.825 59.680 113.245 60.100 ;
        RECT 113.435 59.680 113.855 60.100 ;
        RECT 133.480 62.400 133.995 62.820 ;
        RECT 134.185 62.400 134.605 62.820 ;
        RECT 134.795 62.400 135.215 62.820 ;
        RECT 135.405 62.400 135.825 62.820 ;
        RECT 136.625 62.400 137.045 62.820 ;
        RECT 137.235 62.400 137.655 62.820 ;
        RECT 137.845 62.400 138.265 62.820 ;
        RECT 138.455 62.400 138.970 62.820 ;
        RECT 126.865 59.680 127.285 60.100 ;
        RECT 127.475 59.680 127.895 60.100 ;
        RECT 128.085 59.680 128.505 60.100 ;
        RECT 129.485 59.680 129.905 60.100 ;
        RECT 130.095 59.680 130.515 60.100 ;
        RECT 130.705 59.680 131.125 60.100 ;
        RECT 131.315 59.680 131.830 60.100 ;
        RECT 106.425 52.725 107.045 53.445 ;
        RECT 111.910 52.790 112.940 53.380 ;
        RECT 113.130 52.790 113.580 53.380 ;
        RECT 104.590 48.800 105.010 49.220 ;
        RECT 105.200 48.800 105.620 49.220 ;
        RECT 105.810 48.800 106.230 49.220 ;
        RECT 92.660 46.080 93.175 46.500 ;
        RECT 93.365 46.080 93.785 46.500 ;
        RECT 93.975 46.080 94.395 46.500 ;
        RECT 94.585 46.080 95.005 46.500 ;
        RECT 96.060 46.080 96.480 46.500 ;
        RECT 96.670 46.080 97.090 46.500 ;
        RECT 97.280 46.080 97.700 46.500 ;
        RECT 97.890 46.080 98.310 46.500 ;
        RECT 98.500 46.080 98.920 46.500 ;
        RECT 99.985 46.080 100.405 46.500 ;
        RECT 100.595 46.080 101.015 46.500 ;
        RECT 101.205 46.080 101.625 46.500 ;
        RECT 101.815 46.080 102.330 46.500 ;
        RECT 115.510 48.800 116.025 49.220 ;
        RECT 116.215 48.800 116.635 49.220 ;
        RECT 116.825 48.800 117.245 49.220 ;
        RECT 117.435 48.800 117.855 49.220 ;
        RECT 118.655 48.800 119.075 49.220 ;
        RECT 119.265 48.800 119.685 49.220 ;
        RECT 119.875 48.800 120.295 49.220 ;
        RECT 120.485 48.800 121.000 49.220 ;
        RECT 108.365 46.080 108.785 46.500 ;
        RECT 108.975 46.080 109.395 46.500 ;
        RECT 109.585 46.080 110.005 46.500 ;
        RECT 110.195 46.080 110.710 46.500 ;
        RECT 111.510 46.080 112.025 46.500 ;
        RECT 112.215 46.080 112.635 46.500 ;
        RECT 112.825 46.080 113.245 46.500 ;
        RECT 113.435 46.080 113.855 46.500 ;
        RECT 130.070 52.610 131.080 53.550 ;
        RECT 145.010 62.400 145.525 62.820 ;
        RECT 145.715 62.400 146.135 62.820 ;
        RECT 146.325 62.400 146.745 62.820 ;
        RECT 146.935 62.400 147.355 62.820 ;
        RECT 148.420 62.400 148.840 62.820 ;
        RECT 149.030 62.400 149.450 62.820 ;
        RECT 149.640 62.400 150.060 62.820 ;
        RECT 150.250 62.400 150.670 62.820 ;
        RECT 150.860 62.400 151.280 62.820 ;
        RECT 152.335 62.400 152.755 62.820 ;
        RECT 152.945 62.400 153.365 62.820 ;
        RECT 153.555 62.400 153.975 62.820 ;
        RECT 154.165 62.400 154.680 62.820 ;
        RECT 141.715 59.680 142.135 60.100 ;
        RECT 142.325 59.680 142.745 60.100 ;
        RECT 142.935 59.680 143.355 60.100 ;
        RECT 162.980 62.400 163.495 62.820 ;
        RECT 163.685 62.400 164.105 62.820 ;
        RECT 164.295 62.400 164.715 62.820 ;
        RECT 164.905 62.400 165.325 62.820 ;
        RECT 166.125 62.400 166.545 62.820 ;
        RECT 166.735 62.400 167.155 62.820 ;
        RECT 167.345 62.400 167.765 62.820 ;
        RECT 167.955 62.400 168.470 62.820 ;
        RECT 156.365 59.680 156.785 60.100 ;
        RECT 156.975 59.680 157.395 60.100 ;
        RECT 157.585 59.680 158.005 60.100 ;
        RECT 158.985 59.680 159.405 60.100 ;
        RECT 159.595 59.680 160.015 60.100 ;
        RECT 160.205 59.680 160.625 60.100 ;
        RECT 160.815 59.680 161.330 60.100 ;
        RECT 135.925 52.725 136.545 53.445 ;
        RECT 141.410 52.790 142.440 53.380 ;
        RECT 142.630 52.790 143.080 53.380 ;
        RECT 134.090 48.800 134.510 49.220 ;
        RECT 134.700 48.800 135.120 49.220 ;
        RECT 135.310 48.800 135.730 49.220 ;
        RECT 122.160 46.080 122.675 46.500 ;
        RECT 122.865 46.080 123.285 46.500 ;
        RECT 123.475 46.080 123.895 46.500 ;
        RECT 124.085 46.080 124.505 46.500 ;
        RECT 125.560 46.080 125.980 46.500 ;
        RECT 126.170 46.080 126.590 46.500 ;
        RECT 126.780 46.080 127.200 46.500 ;
        RECT 127.390 46.080 127.810 46.500 ;
        RECT 128.000 46.080 128.420 46.500 ;
        RECT 129.485 46.080 129.905 46.500 ;
        RECT 130.095 46.080 130.515 46.500 ;
        RECT 130.705 46.080 131.125 46.500 ;
        RECT 131.315 46.080 131.830 46.500 ;
        RECT 145.010 48.800 145.525 49.220 ;
        RECT 145.715 48.800 146.135 49.220 ;
        RECT 146.325 48.800 146.745 49.220 ;
        RECT 146.935 48.800 147.355 49.220 ;
        RECT 148.155 48.800 148.575 49.220 ;
        RECT 148.765 48.800 149.185 49.220 ;
        RECT 149.375 48.800 149.795 49.220 ;
        RECT 149.985 48.800 150.500 49.220 ;
        RECT 137.865 46.080 138.285 46.500 ;
        RECT 138.475 46.080 138.895 46.500 ;
        RECT 139.085 46.080 139.505 46.500 ;
        RECT 139.695 46.080 140.210 46.500 ;
        RECT 141.010 46.080 141.525 46.500 ;
        RECT 141.715 46.080 142.135 46.500 ;
        RECT 142.325 46.080 142.745 46.500 ;
        RECT 142.935 46.080 143.355 46.500 ;
        RECT 159.570 52.610 160.580 53.550 ;
        RECT 174.510 62.400 175.025 62.820 ;
        RECT 175.215 62.400 175.635 62.820 ;
        RECT 175.825 62.400 176.245 62.820 ;
        RECT 176.435 62.400 176.855 62.820 ;
        RECT 177.920 62.400 178.340 62.820 ;
        RECT 178.530 62.400 178.950 62.820 ;
        RECT 179.140 62.400 179.560 62.820 ;
        RECT 179.750 62.400 180.170 62.820 ;
        RECT 180.360 62.400 180.780 62.820 ;
        RECT 181.835 62.400 182.255 62.820 ;
        RECT 182.445 62.400 182.865 62.820 ;
        RECT 183.055 62.400 183.475 62.820 ;
        RECT 183.665 62.400 184.180 62.820 ;
        RECT 171.215 59.680 171.635 60.100 ;
        RECT 171.825 59.680 172.245 60.100 ;
        RECT 172.435 59.680 172.855 60.100 ;
        RECT 192.480 62.400 192.995 62.820 ;
        RECT 193.185 62.400 193.605 62.820 ;
        RECT 193.795 62.400 194.215 62.820 ;
        RECT 194.405 62.400 194.825 62.820 ;
        RECT 195.625 62.400 196.045 62.820 ;
        RECT 196.235 62.400 196.655 62.820 ;
        RECT 196.845 62.400 197.265 62.820 ;
        RECT 197.455 62.400 197.970 62.820 ;
        RECT 185.865 59.680 186.285 60.100 ;
        RECT 186.475 59.680 186.895 60.100 ;
        RECT 187.085 59.680 187.505 60.100 ;
        RECT 188.485 59.680 188.905 60.100 ;
        RECT 189.095 59.680 189.515 60.100 ;
        RECT 189.705 59.680 190.125 60.100 ;
        RECT 190.315 59.680 190.830 60.100 ;
        RECT 165.425 52.725 166.045 53.445 ;
        RECT 170.910 52.790 171.940 53.380 ;
        RECT 172.130 52.790 172.580 53.380 ;
        RECT 163.590 48.800 164.010 49.220 ;
        RECT 164.200 48.800 164.620 49.220 ;
        RECT 164.810 48.800 165.230 49.220 ;
        RECT 151.660 46.080 152.175 46.500 ;
        RECT 152.365 46.080 152.785 46.500 ;
        RECT 152.975 46.080 153.395 46.500 ;
        RECT 153.585 46.080 154.005 46.500 ;
        RECT 155.060 46.080 155.480 46.500 ;
        RECT 155.670 46.080 156.090 46.500 ;
        RECT 156.280 46.080 156.700 46.500 ;
        RECT 156.890 46.080 157.310 46.500 ;
        RECT 157.500 46.080 157.920 46.500 ;
        RECT 158.985 46.080 159.405 46.500 ;
        RECT 159.595 46.080 160.015 46.500 ;
        RECT 160.205 46.080 160.625 46.500 ;
        RECT 160.815 46.080 161.330 46.500 ;
        RECT 174.510 48.800 175.025 49.220 ;
        RECT 175.215 48.800 175.635 49.220 ;
        RECT 175.825 48.800 176.245 49.220 ;
        RECT 176.435 48.800 176.855 49.220 ;
        RECT 177.655 48.800 178.075 49.220 ;
        RECT 178.265 48.800 178.685 49.220 ;
        RECT 178.875 48.800 179.295 49.220 ;
        RECT 179.485 48.800 180.000 49.220 ;
        RECT 167.365 46.080 167.785 46.500 ;
        RECT 167.975 46.080 168.395 46.500 ;
        RECT 168.585 46.080 169.005 46.500 ;
        RECT 169.195 46.080 169.710 46.500 ;
        RECT 170.510 46.080 171.025 46.500 ;
        RECT 171.215 46.080 171.635 46.500 ;
        RECT 171.825 46.080 172.245 46.500 ;
        RECT 172.435 46.080 172.855 46.500 ;
        RECT 189.070 52.610 190.080 53.550 ;
        RECT 204.010 62.400 204.525 62.820 ;
        RECT 204.715 62.400 205.135 62.820 ;
        RECT 205.325 62.400 205.745 62.820 ;
        RECT 205.935 62.400 206.355 62.820 ;
        RECT 207.420 62.400 207.840 62.820 ;
        RECT 208.030 62.400 208.450 62.820 ;
        RECT 208.640 62.400 209.060 62.820 ;
        RECT 209.250 62.400 209.670 62.820 ;
        RECT 209.860 62.400 210.280 62.820 ;
        RECT 211.335 62.400 211.755 62.820 ;
        RECT 211.945 62.400 212.365 62.820 ;
        RECT 212.555 62.400 212.975 62.820 ;
        RECT 213.165 62.400 213.680 62.820 ;
        RECT 200.715 59.680 201.135 60.100 ;
        RECT 201.325 59.680 201.745 60.100 ;
        RECT 201.935 59.680 202.355 60.100 ;
        RECT 221.980 62.400 222.495 62.820 ;
        RECT 222.685 62.400 223.105 62.820 ;
        RECT 223.295 62.400 223.715 62.820 ;
        RECT 223.905 62.400 224.325 62.820 ;
        RECT 225.125 62.400 225.545 62.820 ;
        RECT 225.735 62.400 226.155 62.820 ;
        RECT 226.345 62.400 226.765 62.820 ;
        RECT 226.955 62.400 227.470 62.820 ;
        RECT 215.365 59.680 215.785 60.100 ;
        RECT 215.975 59.680 216.395 60.100 ;
        RECT 216.585 59.680 217.005 60.100 ;
        RECT 217.985 59.680 218.405 60.100 ;
        RECT 218.595 59.680 219.015 60.100 ;
        RECT 219.205 59.680 219.625 60.100 ;
        RECT 219.815 59.680 220.330 60.100 ;
        RECT 194.925 52.725 195.545 53.445 ;
        RECT 200.410 52.790 201.440 53.380 ;
        RECT 201.630 52.790 202.080 53.380 ;
        RECT 193.090 48.800 193.510 49.220 ;
        RECT 193.700 48.800 194.120 49.220 ;
        RECT 194.310 48.800 194.730 49.220 ;
        RECT 181.160 46.080 181.675 46.500 ;
        RECT 181.865 46.080 182.285 46.500 ;
        RECT 182.475 46.080 182.895 46.500 ;
        RECT 183.085 46.080 183.505 46.500 ;
        RECT 184.560 46.080 184.980 46.500 ;
        RECT 185.170 46.080 185.590 46.500 ;
        RECT 185.780 46.080 186.200 46.500 ;
        RECT 186.390 46.080 186.810 46.500 ;
        RECT 187.000 46.080 187.420 46.500 ;
        RECT 188.485 46.080 188.905 46.500 ;
        RECT 189.095 46.080 189.515 46.500 ;
        RECT 189.705 46.080 190.125 46.500 ;
        RECT 190.315 46.080 190.830 46.500 ;
        RECT 204.010 48.800 204.525 49.220 ;
        RECT 204.715 48.800 205.135 49.220 ;
        RECT 205.325 48.800 205.745 49.220 ;
        RECT 205.935 48.800 206.355 49.220 ;
        RECT 207.155 48.800 207.575 49.220 ;
        RECT 207.765 48.800 208.185 49.220 ;
        RECT 208.375 48.800 208.795 49.220 ;
        RECT 208.985 48.800 209.500 49.220 ;
        RECT 196.865 46.080 197.285 46.500 ;
        RECT 197.475 46.080 197.895 46.500 ;
        RECT 198.085 46.080 198.505 46.500 ;
        RECT 198.695 46.080 199.210 46.500 ;
        RECT 200.010 46.080 200.525 46.500 ;
        RECT 200.715 46.080 201.135 46.500 ;
        RECT 201.325 46.080 201.745 46.500 ;
        RECT 201.935 46.080 202.355 46.500 ;
        RECT 218.570 52.610 219.580 53.550 ;
        RECT 233.510 62.400 234.025 62.820 ;
        RECT 234.215 62.400 234.635 62.820 ;
        RECT 234.825 62.400 235.245 62.820 ;
        RECT 235.435 62.400 235.855 62.820 ;
        RECT 236.920 62.400 237.340 62.820 ;
        RECT 237.530 62.400 237.950 62.820 ;
        RECT 238.140 62.400 238.560 62.820 ;
        RECT 238.750 62.400 239.170 62.820 ;
        RECT 239.360 62.400 239.780 62.820 ;
        RECT 240.835 62.400 241.255 62.820 ;
        RECT 241.445 62.400 241.865 62.820 ;
        RECT 242.055 62.400 242.475 62.820 ;
        RECT 242.665 62.400 243.180 62.820 ;
        RECT 230.215 59.680 230.635 60.100 ;
        RECT 230.825 59.680 231.245 60.100 ;
        RECT 231.435 59.680 231.855 60.100 ;
        RECT 244.865 59.680 245.285 60.100 ;
        RECT 245.475 59.680 245.895 60.100 ;
        RECT 246.085 59.680 246.505 60.100 ;
        RECT 247.485 59.680 247.905 60.100 ;
        RECT 248.095 59.680 248.515 60.100 ;
        RECT 248.705 59.680 249.125 60.100 ;
        RECT 249.315 59.680 249.830 60.100 ;
        RECT 224.425 52.725 225.045 53.445 ;
        RECT 229.910 52.790 230.940 53.380 ;
        RECT 231.130 52.790 231.580 53.380 ;
        RECT 222.590 48.800 223.010 49.220 ;
        RECT 223.200 48.800 223.620 49.220 ;
        RECT 223.810 48.800 224.230 49.220 ;
        RECT 210.660 46.080 211.175 46.500 ;
        RECT 211.365 46.080 211.785 46.500 ;
        RECT 211.975 46.080 212.395 46.500 ;
        RECT 212.585 46.080 213.005 46.500 ;
        RECT 214.060 46.080 214.480 46.500 ;
        RECT 214.670 46.080 215.090 46.500 ;
        RECT 215.280 46.080 215.700 46.500 ;
        RECT 215.890 46.080 216.310 46.500 ;
        RECT 216.500 46.080 216.920 46.500 ;
        RECT 217.985 46.080 218.405 46.500 ;
        RECT 218.595 46.080 219.015 46.500 ;
        RECT 219.205 46.080 219.625 46.500 ;
        RECT 219.815 46.080 220.330 46.500 ;
        RECT 233.510 48.800 234.025 49.220 ;
        RECT 234.215 48.800 234.635 49.220 ;
        RECT 234.825 48.800 235.245 49.220 ;
        RECT 235.435 48.800 235.855 49.220 ;
        RECT 236.655 48.800 237.075 49.220 ;
        RECT 237.265 48.800 237.685 49.220 ;
        RECT 237.875 48.800 238.295 49.220 ;
        RECT 238.485 48.800 239.000 49.220 ;
        RECT 226.365 46.080 226.785 46.500 ;
        RECT 226.975 46.080 227.395 46.500 ;
        RECT 227.585 46.080 228.005 46.500 ;
        RECT 228.195 46.080 228.710 46.500 ;
        RECT 229.510 46.080 230.025 46.500 ;
        RECT 230.215 46.080 230.635 46.500 ;
        RECT 230.825 46.080 231.245 46.500 ;
        RECT 231.435 46.080 231.855 46.500 ;
        RECT 248.070 52.610 249.080 53.550 ;
        RECT 240.160 46.080 240.675 46.500 ;
        RECT 240.865 46.080 241.285 46.500 ;
        RECT 241.475 46.080 241.895 46.500 ;
        RECT 242.085 46.080 242.505 46.500 ;
        RECT 243.560 46.080 243.980 46.500 ;
        RECT 244.170 46.080 244.590 46.500 ;
        RECT 244.780 46.080 245.200 46.500 ;
        RECT 245.390 46.080 245.810 46.500 ;
        RECT 246.000 46.080 246.420 46.500 ;
        RECT 247.485 46.080 247.905 46.500 ;
        RECT 248.095 46.080 248.515 46.500 ;
        RECT 248.705 46.080 249.125 46.500 ;
        RECT 249.315 46.080 249.830 46.500 ;
      LAYER met1 ;
        RECT 73.510 84.130 245.000 84.610 ;
        RECT 71.510 81.410 243.950 81.890 ;
        RECT 90.800 77.905 91.930 78.130 ;
        RECT 114.805 77.905 115.545 77.965 ;
        RECT 120.300 77.905 121.430 78.130 ;
        RECT 144.305 77.905 145.045 77.965 ;
        RECT 149.800 77.905 150.930 78.130 ;
        RECT 173.805 77.905 174.545 77.965 ;
        RECT 179.300 77.905 180.430 78.130 ;
        RECT 203.305 77.905 204.045 77.965 ;
        RECT 208.800 77.905 209.930 78.130 ;
        RECT 232.805 77.905 233.545 77.965 ;
        RECT 89.350 77.245 91.930 77.905 ;
        RECT 106.570 77.900 121.430 77.905 ;
        RECT 136.070 77.900 150.930 77.905 ;
        RECT 165.570 77.900 180.430 77.905 ;
        RECT 195.070 77.900 209.930 77.905 ;
        RECT 224.570 77.900 236.950 77.905 ;
        RECT 90.800 77.030 91.930 77.245 ;
        RECT 96.800 77.245 121.430 77.900 ;
        RECT 96.800 77.240 110.060 77.245 ;
        RECT 114.805 77.185 115.545 77.245 ;
        RECT 120.300 77.030 121.430 77.245 ;
        RECT 126.300 77.245 150.930 77.900 ;
        RECT 126.300 77.240 139.560 77.245 ;
        RECT 144.305 77.185 145.045 77.245 ;
        RECT 149.800 77.030 150.930 77.245 ;
        RECT 155.800 77.245 180.430 77.900 ;
        RECT 155.800 77.240 169.060 77.245 ;
        RECT 173.805 77.185 174.545 77.245 ;
        RECT 179.300 77.030 180.430 77.245 ;
        RECT 185.300 77.245 209.930 77.900 ;
        RECT 185.300 77.240 198.560 77.245 ;
        RECT 203.305 77.185 204.045 77.245 ;
        RECT 208.800 77.030 209.930 77.245 ;
        RECT 214.800 77.245 236.950 77.900 ;
        RECT 214.800 77.240 228.060 77.245 ;
        RECT 232.805 77.185 233.545 77.245 ;
        RECT 71.510 73.250 254.240 73.730 ;
        RECT 243.950 72.430 245.910 73.250 ;
        RECT 71.510 70.530 243.950 71.010 ;
        RECT 89.400 68.280 236.900 68.290 ;
        RECT 73.510 67.800 249.040 68.280 ;
        RECT 247.080 67.450 249.040 67.800 ;
        RECT 73.510 62.370 251.950 62.850 ;
        RECT 71.510 59.650 250.950 60.130 ;
        RECT 76.865 53.415 77.605 53.475 ;
        RECT 82.350 53.415 95.610 53.420 ;
        RECT 73.510 52.760 95.610 53.415 ;
        RECT 100.480 53.415 101.610 53.630 ;
        RECT 106.365 53.415 107.105 53.475 ;
        RECT 111.850 53.415 125.110 53.420 ;
        RECT 100.480 52.760 125.110 53.415 ;
        RECT 129.980 53.415 131.110 53.630 ;
        RECT 135.865 53.415 136.605 53.475 ;
        RECT 141.350 53.415 154.610 53.420 ;
        RECT 129.980 52.760 154.610 53.415 ;
        RECT 159.480 53.415 160.610 53.630 ;
        RECT 165.365 53.415 166.105 53.475 ;
        RECT 170.850 53.415 184.110 53.420 ;
        RECT 159.480 52.760 184.110 53.415 ;
        RECT 188.980 53.415 190.110 53.630 ;
        RECT 194.865 53.415 195.605 53.475 ;
        RECT 200.350 53.415 213.610 53.420 ;
        RECT 188.980 52.760 213.610 53.415 ;
        RECT 218.480 53.415 219.610 53.630 ;
        RECT 224.365 53.415 225.105 53.475 ;
        RECT 229.850 53.415 243.110 53.420 ;
        RECT 218.480 52.760 243.110 53.415 ;
        RECT 247.980 53.415 249.110 53.630 ;
        RECT 247.980 53.385 250.510 53.415 ;
        RECT 244.150 52.785 250.510 53.385 ;
        RECT 73.510 52.755 85.840 52.760 ;
        RECT 100.480 52.755 115.340 52.760 ;
        RECT 129.980 52.755 144.840 52.760 ;
        RECT 159.480 52.755 174.340 52.760 ;
        RECT 188.980 52.755 203.840 52.760 ;
        RECT 218.480 52.755 233.340 52.760 ;
        RECT 247.980 52.755 250.510 52.785 ;
        RECT 76.865 52.695 77.605 52.755 ;
        RECT 100.480 52.530 101.610 52.755 ;
        RECT 106.365 52.695 107.105 52.755 ;
        RECT 129.980 52.530 131.110 52.755 ;
        RECT 135.865 52.695 136.605 52.755 ;
        RECT 159.480 52.530 160.610 52.755 ;
        RECT 165.365 52.695 166.105 52.755 ;
        RECT 188.980 52.530 190.110 52.755 ;
        RECT 194.865 52.695 195.605 52.755 ;
        RECT 218.480 52.530 219.610 52.755 ;
        RECT 224.365 52.695 225.105 52.755 ;
        RECT 247.980 52.530 249.110 52.755 ;
        RECT 71.510 48.770 250.950 49.250 ;
        RECT 73.510 46.050 251.950 46.530 ;
      LAYER via ;
        RECT 243.950 84.130 244.950 84.610 ;
        RECT 89.400 77.245 90.295 77.905 ;
        RECT 235.980 77.245 236.900 77.905 ;
        RECT 243.950 67.800 245.950 68.280 ;
        RECT 250.950 62.370 251.900 62.850 ;
        RECT 75.505 52.755 76.205 53.415 ;
        RECT 244.210 52.785 244.910 53.385 ;
        RECT 250.950 46.050 251.920 46.530 ;
      LAYER met2 ;
        RECT 198.000 84.130 200.000 84.610 ;
        RECT 90.000 81.410 92.000 81.890 ;
        RECT 108.000 81.410 110.000 81.890 ;
        RECT 126.000 81.410 128.000 81.890 ;
        RECT 162.000 81.410 164.000 81.890 ;
        RECT 234.000 81.410 236.000 81.890 ;
        RECT 89.400 77.925 90.295 77.955 ;
        RECT 85.930 77.225 90.295 77.925 ;
        RECT 85.930 66.340 86.630 77.225 ;
        RECT 89.400 77.195 90.295 77.225 ;
        RECT 235.980 77.925 236.900 77.955 ;
        RECT 235.980 77.225 241.000 77.925 ;
        RECT 235.980 77.195 236.900 77.225 ;
        RECT 90.000 70.530 92.000 71.010 ;
        RECT 108.000 70.530 110.000 71.010 ;
        RECT 126.000 70.530 128.000 71.010 ;
        RECT 198.000 70.530 200.000 71.010 ;
        RECT 234.000 67.800 236.000 68.280 ;
        RECT 75.510 65.640 86.630 66.340 ;
        RECT 75.510 64.825 76.210 65.640 ;
        RECT 75.505 59.255 76.210 64.825 ;
        RECT 240.300 63.925 241.000 77.225 ;
        RECT 243.950 68.530 244.950 84.660 ;
        RECT 252.000 73.250 254.000 73.730 ;
        RECT 243.950 67.530 251.950 68.530 ;
        RECT 250.950 66.990 251.945 67.530 ;
        RECT 240.300 63.225 244.910 63.925 ;
        RECT 234.000 62.370 236.000 62.850 ;
        RECT 90.000 59.650 92.000 60.130 ;
        RECT 108.000 59.650 110.000 60.130 ;
        RECT 126.000 59.650 128.000 60.130 ;
        RECT 162.000 59.650 164.000 60.130 ;
        RECT 198.000 59.650 200.000 60.130 ;
        RECT 75.505 52.705 76.205 59.255 ;
        RECT 244.210 52.735 244.910 63.225 ;
        RECT 90.000 48.770 92.000 49.250 ;
        RECT 108.000 48.770 110.000 49.250 ;
        RECT 126.000 48.770 128.000 49.250 ;
        RECT 198.000 48.770 200.000 49.250 ;
        RECT 234.000 48.770 236.000 49.250 ;
        RECT 250.950 46.000 251.950 66.990 ;
  END
END vco
END LIBRARY

