VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_adc_wrapper
  CLASS BLOCK ;
  FOREIGN vco_adc_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 600.000 ;
  PIN adc0_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 2.760 900.000 3.360 ;
    END
  END adc0_dat_i[0]
  PIN adc0_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 184.320 900.000 184.920 ;
    END
  END adc0_dat_i[10]
  PIN adc0_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 200.640 900.000 201.240 ;
    END
  END adc0_dat_i[11]
  PIN adc0_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 216.960 900.000 217.560 ;
    END
  END adc0_dat_i[12]
  PIN adc0_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 233.280 900.000 233.880 ;
    END
  END adc0_dat_i[13]
  PIN adc0_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 250.280 900.000 250.880 ;
    END
  END adc0_dat_i[14]
  PIN adc0_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 266.600 900.000 267.200 ;
    END
  END adc0_dat_i[15]
  PIN adc0_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 282.920 900.000 283.520 ;
    END
  END adc0_dat_i[16]
  PIN adc0_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 299.240 900.000 299.840 ;
    END
  END adc0_dat_i[17]
  PIN adc0_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 316.240 900.000 316.840 ;
    END
  END adc0_dat_i[18]
  PIN adc0_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 332.560 900.000 333.160 ;
    END
  END adc0_dat_i[19]
  PIN adc0_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 24.520 900.000 25.120 ;
    END
  END adc0_dat_i[1]
  PIN adc0_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 348.880 900.000 349.480 ;
    END
  END adc0_dat_i[20]
  PIN adc0_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 365.880 900.000 366.480 ;
    END
  END adc0_dat_i[21]
  PIN adc0_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 382.200 900.000 382.800 ;
    END
  END adc0_dat_i[22]
  PIN adc0_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 398.520 900.000 399.120 ;
    END
  END adc0_dat_i[23]
  PIN adc0_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 414.840 900.000 415.440 ;
    END
  END adc0_dat_i[24]
  PIN adc0_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 431.840 900.000 432.440 ;
    END
  END adc0_dat_i[25]
  PIN adc0_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 448.160 900.000 448.760 ;
    END
  END adc0_dat_i[26]
  PIN adc0_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 464.480 900.000 465.080 ;
    END
  END adc0_dat_i[27]
  PIN adc0_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 480.800 900.000 481.400 ;
    END
  END adc0_dat_i[28]
  PIN adc0_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 497.800 900.000 498.400 ;
    END
  END adc0_dat_i[29]
  PIN adc0_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 46.280 900.000 46.880 ;
    END
  END adc0_dat_i[2]
  PIN adc0_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 514.120 900.000 514.720 ;
    END
  END adc0_dat_i[30]
  PIN adc0_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 530.440 900.000 531.040 ;
    END
  END adc0_dat_i[31]
  PIN adc0_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 68.720 900.000 69.320 ;
    END
  END adc0_dat_i[3]
  PIN adc0_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 85.040 900.000 85.640 ;
    END
  END adc0_dat_i[4]
  PIN adc0_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 101.360 900.000 101.960 ;
    END
  END adc0_dat_i[5]
  PIN adc0_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 117.680 900.000 118.280 ;
    END
  END adc0_dat_i[6]
  PIN adc0_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 134.680 900.000 135.280 ;
    END
  END adc0_dat_i[7]
  PIN adc0_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 151.000 900.000 151.600 ;
    END
  END adc0_dat_i[8]
  PIN adc0_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 167.320 900.000 167.920 ;
    END
  END adc0_dat_i[9]
  PIN adc1_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 8.200 900.000 8.800 ;
    END
  END adc1_dat_i[0]
  PIN adc1_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 189.760 900.000 190.360 ;
    END
  END adc1_dat_i[10]
  PIN adc1_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 206.080 900.000 206.680 ;
    END
  END adc1_dat_i[11]
  PIN adc1_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 222.400 900.000 223.000 ;
    END
  END adc1_dat_i[12]
  PIN adc1_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 238.720 900.000 239.320 ;
    END
  END adc1_dat_i[13]
  PIN adc1_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 255.720 900.000 256.320 ;
    END
  END adc1_dat_i[14]
  PIN adc1_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 272.040 900.000 272.640 ;
    END
  END adc1_dat_i[15]
  PIN adc1_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 288.360 900.000 288.960 ;
    END
  END adc1_dat_i[16]
  PIN adc1_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 305.360 900.000 305.960 ;
    END
  END adc1_dat_i[17]
  PIN adc1_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 321.680 900.000 322.280 ;
    END
  END adc1_dat_i[18]
  PIN adc1_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 338.000 900.000 338.600 ;
    END
  END adc1_dat_i[19]
  PIN adc1_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 29.960 900.000 30.560 ;
    END
  END adc1_dat_i[1]
  PIN adc1_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 354.320 900.000 354.920 ;
    END
  END adc1_dat_i[20]
  PIN adc1_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 371.320 900.000 371.920 ;
    END
  END adc1_dat_i[21]
  PIN adc1_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 387.640 900.000 388.240 ;
    END
  END adc1_dat_i[22]
  PIN adc1_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 403.960 900.000 404.560 ;
    END
  END adc1_dat_i[23]
  PIN adc1_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 420.280 900.000 420.880 ;
    END
  END adc1_dat_i[24]
  PIN adc1_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 437.280 900.000 437.880 ;
    END
  END adc1_dat_i[25]
  PIN adc1_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 453.600 900.000 454.200 ;
    END
  END adc1_dat_i[26]
  PIN adc1_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 469.920 900.000 470.520 ;
    END
  END adc1_dat_i[27]
  PIN adc1_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 486.920 900.000 487.520 ;
    END
  END adc1_dat_i[28]
  PIN adc1_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 503.240 900.000 503.840 ;
    END
  END adc1_dat_i[29]
  PIN adc1_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 51.720 900.000 52.320 ;
    END
  END adc1_dat_i[2]
  PIN adc1_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 519.560 900.000 520.160 ;
    END
  END adc1_dat_i[30]
  PIN adc1_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 535.880 900.000 536.480 ;
    END
  END adc1_dat_i[31]
  PIN adc1_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 74.160 900.000 74.760 ;
    END
  END adc1_dat_i[3]
  PIN adc1_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 90.480 900.000 91.080 ;
    END
  END adc1_dat_i[4]
  PIN adc1_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 106.800 900.000 107.400 ;
    END
  END adc1_dat_i[5]
  PIN adc1_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 123.800 900.000 124.400 ;
    END
  END adc1_dat_i[6]
  PIN adc1_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 140.120 900.000 140.720 ;
    END
  END adc1_dat_i[7]
  PIN adc1_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 156.440 900.000 157.040 ;
    END
  END adc1_dat_i[8]
  PIN adc1_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 172.760 900.000 173.360 ;
    END
  END adc1_dat_i[9]
  PIN adc2_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 13.640 900.000 14.240 ;
    END
  END adc2_dat_i[0]
  PIN adc2_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 195.200 900.000 195.800 ;
    END
  END adc2_dat_i[10]
  PIN adc2_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 211.520 900.000 212.120 ;
    END
  END adc2_dat_i[11]
  PIN adc2_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 227.840 900.000 228.440 ;
    END
  END adc2_dat_i[12]
  PIN adc2_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 244.840 900.000 245.440 ;
    END
  END adc2_dat_i[13]
  PIN adc2_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 261.160 900.000 261.760 ;
    END
  END adc2_dat_i[14]
  PIN adc2_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 277.480 900.000 278.080 ;
    END
  END adc2_dat_i[15]
  PIN adc2_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 293.800 900.000 294.400 ;
    END
  END adc2_dat_i[16]
  PIN adc2_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 310.800 900.000 311.400 ;
    END
  END adc2_dat_i[17]
  PIN adc2_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 327.120 900.000 327.720 ;
    END
  END adc2_dat_i[18]
  PIN adc2_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 343.440 900.000 344.040 ;
    END
  END adc2_dat_i[19]
  PIN adc2_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 35.400 900.000 36.000 ;
    END
  END adc2_dat_i[1]
  PIN adc2_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 359.760 900.000 360.360 ;
    END
  END adc2_dat_i[20]
  PIN adc2_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 376.760 900.000 377.360 ;
    END
  END adc2_dat_i[21]
  PIN adc2_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 393.080 900.000 393.680 ;
    END
  END adc2_dat_i[22]
  PIN adc2_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 409.400 900.000 410.000 ;
    END
  END adc2_dat_i[23]
  PIN adc2_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 426.400 900.000 427.000 ;
    END
  END adc2_dat_i[24]
  PIN adc2_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 442.720 900.000 443.320 ;
    END
  END adc2_dat_i[25]
  PIN adc2_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 459.040 900.000 459.640 ;
    END
  END adc2_dat_i[26]
  PIN adc2_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 475.360 900.000 475.960 ;
    END
  END adc2_dat_i[27]
  PIN adc2_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 492.360 900.000 492.960 ;
    END
  END adc2_dat_i[28]
  PIN adc2_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 508.680 900.000 509.280 ;
    END
  END adc2_dat_i[29]
  PIN adc2_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 57.160 900.000 57.760 ;
    END
  END adc2_dat_i[2]
  PIN adc2_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 525.000 900.000 525.600 ;
    END
  END adc2_dat_i[30]
  PIN adc2_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 541.320 900.000 541.920 ;
    END
  END adc2_dat_i[31]
  PIN adc2_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 79.600 900.000 80.200 ;
    END
  END adc2_dat_i[3]
  PIN adc2_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 95.920 900.000 96.520 ;
    END
  END adc2_dat_i[4]
  PIN adc2_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 112.240 900.000 112.840 ;
    END
  END adc2_dat_i[5]
  PIN adc2_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 129.240 900.000 129.840 ;
    END
  END adc2_dat_i[6]
  PIN adc2_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 145.560 900.000 146.160 ;
    END
  END adc2_dat_i[7]
  PIN adc2_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 161.880 900.000 162.480 ;
    END
  END adc2_dat_i[8]
  PIN adc2_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 178.200 900.000 178.800 ;
    END
  END adc2_dat_i[9]
  PIN adc_dvalid_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 19.080 900.000 19.680 ;
    END
  END adc_dvalid_i[0]
  PIN adc_dvalid_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 40.840 900.000 41.440 ;
    END
  END adc_dvalid_i[1]
  PIN adc_dvalid_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 63.280 900.000 63.880 ;
    END
  END adc_dvalid_i[2]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 596.000 5.430 600.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 596.000 224.850 600.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 596.000 246.930 600.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 596.000 268.550 600.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 596.000 290.630 600.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 596.000 312.710 600.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 596.000 334.330 600.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 596.000 356.410 600.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 596.000 378.490 600.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 596.000 400.570 600.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 596.000 422.190 600.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 596.000 27.050 600.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 596.000 444.270 600.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 596.000 466.350 600.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 596.000 488.430 600.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 596.000 510.050 600.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 596.000 532.130 600.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 596.000 554.210 600.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 596.000 576.290 600.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 596.000 597.910 600.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 596.000 619.990 600.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 596.000 642.070 600.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 596.000 49.130 600.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 596.000 663.690 600.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 596.000 685.770 600.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 596.000 707.850 600.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 596.000 729.930 600.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 596.000 751.550 600.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 596.000 773.630 600.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 596.000 795.710 600.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 596.000 817.790 600.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 596.000 71.210 600.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 596.000 92.830 600.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 596.000 114.910 600.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 596.000 136.990 600.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 596.000 159.070 600.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 596.000 180.690 600.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 596.000 202.770 600.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 596.000 16.010 600.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 596.000 235.890 600.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 596.000 257.510 600.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 596.000 279.590 600.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 596.000 301.670 600.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 596.000 323.750 600.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 596.000 345.370 600.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 596.000 367.450 600.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 596.000 389.530 600.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 596.000 411.610 600.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 596.000 433.230 600.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 596.000 38.090 600.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 596.000 455.310 600.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 596.000 477.390 600.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 596.000 499.010 600.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 596.000 521.090 600.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 596.000 543.170 600.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 596.000 565.250 600.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 596.000 586.870 600.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 596.000 608.950 600.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 596.000 631.030 600.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 596.000 653.110 600.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 596.000 60.170 600.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 596.000 674.730 600.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 596.000 696.810 600.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 596.000 718.890 600.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 596.000 740.970 600.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 596.000 762.590 600.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 596.000 784.670 600.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 596.000 806.750 600.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 596.000 828.370 600.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 596.000 82.250 600.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 596.000 103.870 600.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 596.000 125.950 600.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 596.000 148.030 600.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 596.000 169.650 600.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 596.000 191.730 600.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 596.000 213.810 600.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END irq[2]
  PIN mem1_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.120 4.000 21.720 ;
    END
  END mem1_data_i[0]
  PIN mem1_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END mem1_data_i[10]
  PIN mem1_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.760 4.000 292.360 ;
    END
  END mem1_data_i[11]
  PIN mem1_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END mem1_data_i[12]
  PIN mem1_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 321.000 4.000 321.600 ;
    END
  END mem1_data_i[13]
  PIN mem1_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.960 4.000 336.560 ;
    END
  END mem1_data_i[14]
  PIN mem1_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END mem1_data_i[15]
  PIN mem1_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 365.200 4.000 365.800 ;
    END
  END mem1_data_i[16]
  PIN mem1_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.160 4.000 380.760 ;
    END
  END mem1_data_i[17]
  PIN mem1_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.120 4.000 395.720 ;
    END
  END mem1_data_i[18]
  PIN mem1_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END mem1_data_i[19]
  PIN mem1_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END mem1_data_i[1]
  PIN mem1_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 424.360 4.000 424.960 ;
    END
  END mem1_data_i[20]
  PIN mem1_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 439.320 4.000 439.920 ;
    END
  END mem1_data_i[21]
  PIN mem1_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.280 4.000 454.880 ;
    END
  END mem1_data_i[22]
  PIN mem1_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END mem1_data_i[23]
  PIN mem1_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 483.520 4.000 484.120 ;
    END
  END mem1_data_i[24]
  PIN mem1_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 498.480 4.000 499.080 ;
    END
  END mem1_data_i[25]
  PIN mem1_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END mem1_data_i[26]
  PIN mem1_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END mem1_data_i[27]
  PIN mem1_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 542.680 4.000 543.280 ;
    END
  END mem1_data_i[28]
  PIN mem1_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.960 4.000 557.560 ;
    END
  END mem1_data_i[29]
  PIN mem1_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 90.480 4.000 91.080 ;
    END
  END mem1_data_i[2]
  PIN mem1_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.920 4.000 572.520 ;
    END
  END mem1_data_i[30]
  PIN mem1_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.880 4.000 587.480 ;
    END
  END mem1_data_i[31]
  PIN mem1_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END mem1_data_i[3]
  PIN mem1_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END mem1_data_i[4]
  PIN mem1_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.920 4.000 164.520 ;
    END
  END mem1_data_i[5]
  PIN mem1_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 188.400 4.000 189.000 ;
    END
  END mem1_data_i[6]
  PIN mem1_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END mem1_data_i[7]
  PIN mem1_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END mem1_data_i[8]
  PIN mem1_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 262.520 4.000 263.120 ;
    END
  END mem1_data_i[9]
  PIN mem_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END mem_data_i[0]
  PIN mem_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END mem_data_i[10]
  PIN mem_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END mem_data_i[11]
  PIN mem_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 311.480 4.000 312.080 ;
    END
  END mem_data_i[12]
  PIN mem_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END mem_data_i[13]
  PIN mem_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END mem_data_i[14]
  PIN mem_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END mem_data_i[15]
  PIN mem_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END mem_data_i[16]
  PIN mem_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.920 4.000 385.520 ;
    END
  END mem_data_i[17]
  PIN mem_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.880 4.000 400.480 ;
    END
  END mem_data_i[18]
  PIN mem_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END mem_data_i[19]
  PIN mem_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 60.560 4.000 61.160 ;
    END
  END mem_data_i[1]
  PIN mem_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END mem_data_i[20]
  PIN mem_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END mem_data_i[21]
  PIN mem_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END mem_data_i[22]
  PIN mem_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END mem_data_i[23]
  PIN mem_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.280 4.000 488.880 ;
    END
  END mem_data_i[24]
  PIN mem_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.240 4.000 503.840 ;
    END
  END mem_data_i[25]
  PIN mem_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.200 4.000 518.800 ;
    END
  END mem_data_i[26]
  PIN mem_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 532.480 4.000 533.080 ;
    END
  END mem_data_i[27]
  PIN mem_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END mem_data_i[28]
  PIN mem_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 562.400 4.000 563.000 ;
    END
  END mem_data_i[29]
  PIN mem_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END mem_data_i[2]
  PIN mem_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.680 4.000 577.280 ;
    END
  END mem_data_i[30]
  PIN mem_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END mem_data_i[31]
  PIN mem_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mem_data_i[3]
  PIN mem_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.200 4.000 144.800 ;
    END
  END mem_data_i[4]
  PIN mem_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END mem_data_i[5]
  PIN mem_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END mem_data_i[6]
  PIN mem_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 218.320 4.000 218.920 ;
    END
  END mem_data_i[7]
  PIN mem_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.800 4.000 243.400 ;
    END
  END mem_data_i[8]
  PIN mem_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END mem_data_i[9]
  PIN mem_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END mem_data_o[0]
  PIN mem_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END mem_data_o[10]
  PIN mem_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END mem_data_o[11]
  PIN mem_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END mem_data_o[12]
  PIN mem_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.200 4.000 331.800 ;
    END
  END mem_data_o[13]
  PIN mem_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.160 4.000 346.760 ;
    END
  END mem_data_o[14]
  PIN mem_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END mem_data_o[15]
  PIN mem_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END mem_data_o[16]
  PIN mem_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 390.360 4.000 390.960 ;
    END
  END mem_data_o[17]
  PIN mem_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END mem_data_o[18]
  PIN mem_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END mem_data_o[19]
  PIN mem_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END mem_data_o[1]
  PIN mem_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END mem_data_o[20]
  PIN mem_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.840 4.000 449.440 ;
    END
  END mem_data_o[21]
  PIN mem_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.800 4.000 464.400 ;
    END
  END mem_data_o[22]
  PIN mem_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END mem_data_o[23]
  PIN mem_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END mem_data_o[24]
  PIN mem_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END mem_data_o[25]
  PIN mem_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.960 4.000 523.560 ;
    END
  END mem_data_o[26]
  PIN mem_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END mem_data_o[27]
  PIN mem_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.200 4.000 552.800 ;
    END
  END mem_data_o[28]
  PIN mem_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.160 4.000 567.760 ;
    END
  END mem_data_o[29]
  PIN mem_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END mem_data_o[2]
  PIN mem_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END mem_data_o[30]
  PIN mem_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 596.400 4.000 597.000 ;
    END
  END mem_data_o[31]
  PIN mem_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 124.480 4.000 125.080 ;
    END
  END mem_data_o[3]
  PIN mem_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END mem_data_o[4]
  PIN mem_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END mem_data_o[5]
  PIN mem_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 198.600 4.000 199.200 ;
    END
  END mem_data_o[6]
  PIN mem_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END mem_data_o[7]
  PIN mem_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 247.560 4.000 248.160 ;
    END
  END mem_data_o[8]
  PIN mem_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END mem_data_o[9]
  PIN mem_raddr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END mem_raddr_o[0]
  PIN mem_raddr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END mem_raddr_o[1]
  PIN mem_raddr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END mem_raddr_o[2]
  PIN mem_raddr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END mem_raddr_o[3]
  PIN mem_raddr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END mem_raddr_o[4]
  PIN mem_raddr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 178.880 4.000 179.480 ;
    END
  END mem_raddr_o[5]
  PIN mem_raddr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END mem_raddr_o[6]
  PIN mem_raddr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END mem_raddr_o[7]
  PIN mem_raddr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 252.320 4.000 252.920 ;
    END
  END mem_raddr_o[8]
  PIN mem_renb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END mem_renb_o[0]
  PIN mem_renb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END mem_renb_o[1]
  PIN mem_waddr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END mem_waddr_o[0]
  PIN mem_waddr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.280 4.000 80.880 ;
    END
  END mem_waddr_o[1]
  PIN mem_waddr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END mem_waddr_o[2]
  PIN mem_waddr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END mem_waddr_o[3]
  PIN mem_waddr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.160 4.000 159.760 ;
    END
  END mem_waddr_o[4]
  PIN mem_waddr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END mem_waddr_o[5]
  PIN mem_waddr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END mem_waddr_o[6]
  PIN mem_waddr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 232.600 4.000 233.200 ;
    END
  END mem_waddr_o[7]
  PIN mem_waddr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END mem_waddr_o[8]
  PIN mem_wenb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END mem_wenb_o[0]
  PIN mem_wenb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END mem_wenb_o[1]
  PIN oversample_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 547.440 900.000 548.040 ;
    END
  END oversample_o[0]
  PIN oversample_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 552.880 900.000 553.480 ;
    END
  END oversample_o[1]
  PIN oversample_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 558.320 900.000 558.920 ;
    END
  END oversample_o[2]
  PIN oversample_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 563.760 900.000 564.360 ;
    END
  END oversample_o[3]
  PIN oversample_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 569.200 900.000 569.800 ;
    END
  END oversample_o[4]
  PIN oversample_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 574.640 900.000 575.240 ;
    END
  END oversample_o[5]
  PIN oversample_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 580.080 900.000 580.680 ;
    END
  END oversample_o[6]
  PIN oversample_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 585.520 900.000 586.120 ;
    END
  END oversample_o[7]
  PIN oversample_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 590.960 900.000 591.560 ;
    END
  END oversample_o[8]
  PIN oversample_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 596.400 900.000 597.000 ;
    END
  END oversample_o[9]
  PIN sinc3_en_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 596.000 872.530 600.000 ;
    END
  END sinc3_en_o[0]
  PIN sinc3_en_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 596.000 883.570 600.000 ;
    END
  END sinc3_en_o[1]
  PIN sinc3_en_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 596.000 894.610 600.000 ;
    END
  END sinc3_en_o[2]
  PIN vco_enb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 596.000 839.410 600.000 ;
    END
  END vco_enb_o[0]
  PIN vco_enb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 596.000 850.450 600.000 ;
    END
  END vco_enb_o[1]
  PIN vco_enb_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 596.000 861.490 600.000 ;
    END
  END vco_enb_o[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 0.000 854.590 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.910 0.000 813.190 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 0.000 838.030 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 0.000 746.950 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 0.000 796.630 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END wbs_we_i
  PIN wmask_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END wmask_o[0]
  PIN wmask_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END wmask_o[1]
  PIN wmask_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 11.600 4.000 12.200 ;
    END
  END wmask_o[2]
  PIN wmask_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END wmask_o[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 587.760 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 587.760 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 587.760 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 587.760 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 587.520 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 587.520 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 587.520 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 587.520 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 587.520 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 587.520 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 587.520 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 587.520 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 587.520 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 587.520 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 587.520 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 587.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 6.885 895.015 587.605 ;
      LAYER met1 ;
        RECT 3.750 6.840 896.010 587.760 ;
      LAYER met2 ;
        RECT 3.780 595.720 4.870 596.885 ;
        RECT 5.710 595.720 15.450 596.885 ;
        RECT 16.290 595.720 26.490 596.885 ;
        RECT 27.330 595.720 37.530 596.885 ;
        RECT 38.370 595.720 48.570 596.885 ;
        RECT 49.410 595.720 59.610 596.885 ;
        RECT 60.450 595.720 70.650 596.885 ;
        RECT 71.490 595.720 81.690 596.885 ;
        RECT 82.530 595.720 92.270 596.885 ;
        RECT 93.110 595.720 103.310 596.885 ;
        RECT 104.150 595.720 114.350 596.885 ;
        RECT 115.190 595.720 125.390 596.885 ;
        RECT 126.230 595.720 136.430 596.885 ;
        RECT 137.270 595.720 147.470 596.885 ;
        RECT 148.310 595.720 158.510 596.885 ;
        RECT 159.350 595.720 169.090 596.885 ;
        RECT 169.930 595.720 180.130 596.885 ;
        RECT 180.970 595.720 191.170 596.885 ;
        RECT 192.010 595.720 202.210 596.885 ;
        RECT 203.050 595.720 213.250 596.885 ;
        RECT 214.090 595.720 224.290 596.885 ;
        RECT 225.130 595.720 235.330 596.885 ;
        RECT 236.170 595.720 246.370 596.885 ;
        RECT 247.210 595.720 256.950 596.885 ;
        RECT 257.790 595.720 267.990 596.885 ;
        RECT 268.830 595.720 279.030 596.885 ;
        RECT 279.870 595.720 290.070 596.885 ;
        RECT 290.910 595.720 301.110 596.885 ;
        RECT 301.950 595.720 312.150 596.885 ;
        RECT 312.990 595.720 323.190 596.885 ;
        RECT 324.030 595.720 333.770 596.885 ;
        RECT 334.610 595.720 344.810 596.885 ;
        RECT 345.650 595.720 355.850 596.885 ;
        RECT 356.690 595.720 366.890 596.885 ;
        RECT 367.730 595.720 377.930 596.885 ;
        RECT 378.770 595.720 388.970 596.885 ;
        RECT 389.810 595.720 400.010 596.885 ;
        RECT 400.850 595.720 411.050 596.885 ;
        RECT 411.890 595.720 421.630 596.885 ;
        RECT 422.470 595.720 432.670 596.885 ;
        RECT 433.510 595.720 443.710 596.885 ;
        RECT 444.550 595.720 454.750 596.885 ;
        RECT 455.590 595.720 465.790 596.885 ;
        RECT 466.630 595.720 476.830 596.885 ;
        RECT 477.670 595.720 487.870 596.885 ;
        RECT 488.710 595.720 498.450 596.885 ;
        RECT 499.290 595.720 509.490 596.885 ;
        RECT 510.330 595.720 520.530 596.885 ;
        RECT 521.370 595.720 531.570 596.885 ;
        RECT 532.410 595.720 542.610 596.885 ;
        RECT 543.450 595.720 553.650 596.885 ;
        RECT 554.490 595.720 564.690 596.885 ;
        RECT 565.530 595.720 575.730 596.885 ;
        RECT 576.570 595.720 586.310 596.885 ;
        RECT 587.150 595.720 597.350 596.885 ;
        RECT 598.190 595.720 608.390 596.885 ;
        RECT 609.230 595.720 619.430 596.885 ;
        RECT 620.270 595.720 630.470 596.885 ;
        RECT 631.310 595.720 641.510 596.885 ;
        RECT 642.350 595.720 652.550 596.885 ;
        RECT 653.390 595.720 663.130 596.885 ;
        RECT 663.970 595.720 674.170 596.885 ;
        RECT 675.010 595.720 685.210 596.885 ;
        RECT 686.050 595.720 696.250 596.885 ;
        RECT 697.090 595.720 707.290 596.885 ;
        RECT 708.130 595.720 718.330 596.885 ;
        RECT 719.170 595.720 729.370 596.885 ;
        RECT 730.210 595.720 740.410 596.885 ;
        RECT 741.250 595.720 750.990 596.885 ;
        RECT 751.830 595.720 762.030 596.885 ;
        RECT 762.870 595.720 773.070 596.885 ;
        RECT 773.910 595.720 784.110 596.885 ;
        RECT 784.950 595.720 795.150 596.885 ;
        RECT 795.990 595.720 806.190 596.885 ;
        RECT 807.030 595.720 817.230 596.885 ;
        RECT 818.070 595.720 827.810 596.885 ;
        RECT 828.650 595.720 838.850 596.885 ;
        RECT 839.690 595.720 849.890 596.885 ;
        RECT 850.730 595.720 860.930 596.885 ;
        RECT 861.770 595.720 871.970 596.885 ;
        RECT 872.810 595.720 883.010 596.885 ;
        RECT 883.850 595.720 894.050 596.885 ;
        RECT 894.890 595.720 895.980 596.885 ;
        RECT 3.780 4.280 895.980 595.720 ;
        RECT 4.330 2.195 11.310 4.280 ;
        RECT 12.150 2.195 19.590 4.280 ;
        RECT 20.430 2.195 27.870 4.280 ;
        RECT 28.710 2.195 36.150 4.280 ;
        RECT 36.990 2.195 44.430 4.280 ;
        RECT 45.270 2.195 52.710 4.280 ;
        RECT 53.550 2.195 60.990 4.280 ;
        RECT 61.830 2.195 69.270 4.280 ;
        RECT 70.110 2.195 77.550 4.280 ;
        RECT 78.390 2.195 85.830 4.280 ;
        RECT 86.670 2.195 94.110 4.280 ;
        RECT 94.950 2.195 102.390 4.280 ;
        RECT 103.230 2.195 110.670 4.280 ;
        RECT 111.510 2.195 118.950 4.280 ;
        RECT 119.790 2.195 127.230 4.280 ;
        RECT 128.070 2.195 135.510 4.280 ;
        RECT 136.350 2.195 143.790 4.280 ;
        RECT 144.630 2.195 152.070 4.280 ;
        RECT 152.910 2.195 160.350 4.280 ;
        RECT 161.190 2.195 168.630 4.280 ;
        RECT 169.470 2.195 176.910 4.280 ;
        RECT 177.750 2.195 184.730 4.280 ;
        RECT 185.570 2.195 193.010 4.280 ;
        RECT 193.850 2.195 201.290 4.280 ;
        RECT 202.130 2.195 209.570 4.280 ;
        RECT 210.410 2.195 217.850 4.280 ;
        RECT 218.690 2.195 226.130 4.280 ;
        RECT 226.970 2.195 234.410 4.280 ;
        RECT 235.250 2.195 242.690 4.280 ;
        RECT 243.530 2.195 250.970 4.280 ;
        RECT 251.810 2.195 259.250 4.280 ;
        RECT 260.090 2.195 267.530 4.280 ;
        RECT 268.370 2.195 275.810 4.280 ;
        RECT 276.650 2.195 284.090 4.280 ;
        RECT 284.930 2.195 292.370 4.280 ;
        RECT 293.210 2.195 300.650 4.280 ;
        RECT 301.490 2.195 308.930 4.280 ;
        RECT 309.770 2.195 317.210 4.280 ;
        RECT 318.050 2.195 325.490 4.280 ;
        RECT 326.330 2.195 333.770 4.280 ;
        RECT 334.610 2.195 342.050 4.280 ;
        RECT 342.890 2.195 350.330 4.280 ;
        RECT 351.170 2.195 358.610 4.280 ;
        RECT 359.450 2.195 366.430 4.280 ;
        RECT 367.270 2.195 374.710 4.280 ;
        RECT 375.550 2.195 382.990 4.280 ;
        RECT 383.830 2.195 391.270 4.280 ;
        RECT 392.110 2.195 399.550 4.280 ;
        RECT 400.390 2.195 407.830 4.280 ;
        RECT 408.670 2.195 416.110 4.280 ;
        RECT 416.950 2.195 424.390 4.280 ;
        RECT 425.230 2.195 432.670 4.280 ;
        RECT 433.510 2.195 440.950 4.280 ;
        RECT 441.790 2.195 449.230 4.280 ;
        RECT 450.070 2.195 457.510 4.280 ;
        RECT 458.350 2.195 465.790 4.280 ;
        RECT 466.630 2.195 474.070 4.280 ;
        RECT 474.910 2.195 482.350 4.280 ;
        RECT 483.190 2.195 490.630 4.280 ;
        RECT 491.470 2.195 498.910 4.280 ;
        RECT 499.750 2.195 507.190 4.280 ;
        RECT 508.030 2.195 515.470 4.280 ;
        RECT 516.310 2.195 523.750 4.280 ;
        RECT 524.590 2.195 532.030 4.280 ;
        RECT 532.870 2.195 540.310 4.280 ;
        RECT 541.150 2.195 548.130 4.280 ;
        RECT 548.970 2.195 556.410 4.280 ;
        RECT 557.250 2.195 564.690 4.280 ;
        RECT 565.530 2.195 572.970 4.280 ;
        RECT 573.810 2.195 581.250 4.280 ;
        RECT 582.090 2.195 589.530 4.280 ;
        RECT 590.370 2.195 597.810 4.280 ;
        RECT 598.650 2.195 606.090 4.280 ;
        RECT 606.930 2.195 614.370 4.280 ;
        RECT 615.210 2.195 622.650 4.280 ;
        RECT 623.490 2.195 630.930 4.280 ;
        RECT 631.770 2.195 639.210 4.280 ;
        RECT 640.050 2.195 647.490 4.280 ;
        RECT 648.330 2.195 655.770 4.280 ;
        RECT 656.610 2.195 664.050 4.280 ;
        RECT 664.890 2.195 672.330 4.280 ;
        RECT 673.170 2.195 680.610 4.280 ;
        RECT 681.450 2.195 688.890 4.280 ;
        RECT 689.730 2.195 697.170 4.280 ;
        RECT 698.010 2.195 705.450 4.280 ;
        RECT 706.290 2.195 713.730 4.280 ;
        RECT 714.570 2.195 722.010 4.280 ;
        RECT 722.850 2.195 729.830 4.280 ;
        RECT 730.670 2.195 738.110 4.280 ;
        RECT 738.950 2.195 746.390 4.280 ;
        RECT 747.230 2.195 754.670 4.280 ;
        RECT 755.510 2.195 762.950 4.280 ;
        RECT 763.790 2.195 771.230 4.280 ;
        RECT 772.070 2.195 779.510 4.280 ;
        RECT 780.350 2.195 787.790 4.280 ;
        RECT 788.630 2.195 796.070 4.280 ;
        RECT 796.910 2.195 804.350 4.280 ;
        RECT 805.190 2.195 812.630 4.280 ;
        RECT 813.470 2.195 820.910 4.280 ;
        RECT 821.750 2.195 829.190 4.280 ;
        RECT 830.030 2.195 837.470 4.280 ;
        RECT 838.310 2.195 845.750 4.280 ;
        RECT 846.590 2.195 854.030 4.280 ;
        RECT 854.870 2.195 862.310 4.280 ;
        RECT 863.150 2.195 870.590 4.280 ;
        RECT 871.430 2.195 878.870 4.280 ;
        RECT 879.710 2.195 887.150 4.280 ;
        RECT 887.990 2.195 895.430 4.280 ;
      LAYER met3 ;
        RECT 4.400 596.000 895.600 596.865 ;
        RECT 4.000 592.640 896.000 596.000 ;
        RECT 4.400 591.960 896.000 592.640 ;
        RECT 4.400 591.240 895.600 591.960 ;
        RECT 4.000 590.560 895.600 591.240 ;
        RECT 4.000 587.880 896.000 590.560 ;
        RECT 4.400 586.520 896.000 587.880 ;
        RECT 4.400 586.480 895.600 586.520 ;
        RECT 4.000 585.120 895.600 586.480 ;
        RECT 4.000 583.120 896.000 585.120 ;
        RECT 4.400 581.720 896.000 583.120 ;
        RECT 4.000 581.080 896.000 581.720 ;
        RECT 4.000 579.680 895.600 581.080 ;
        RECT 4.000 577.680 896.000 579.680 ;
        RECT 4.400 576.280 896.000 577.680 ;
        RECT 4.000 575.640 896.000 576.280 ;
        RECT 4.000 574.240 895.600 575.640 ;
        RECT 4.000 572.920 896.000 574.240 ;
        RECT 4.400 571.520 896.000 572.920 ;
        RECT 4.000 570.200 896.000 571.520 ;
        RECT 4.000 568.800 895.600 570.200 ;
        RECT 4.000 568.160 896.000 568.800 ;
        RECT 4.400 566.760 896.000 568.160 ;
        RECT 4.000 564.760 896.000 566.760 ;
        RECT 4.000 563.400 895.600 564.760 ;
        RECT 4.400 563.360 895.600 563.400 ;
        RECT 4.400 562.000 896.000 563.360 ;
        RECT 4.000 559.320 896.000 562.000 ;
        RECT 4.000 557.960 895.600 559.320 ;
        RECT 4.400 557.920 895.600 557.960 ;
        RECT 4.400 556.560 896.000 557.920 ;
        RECT 4.000 553.880 896.000 556.560 ;
        RECT 4.000 553.200 895.600 553.880 ;
        RECT 4.400 552.480 895.600 553.200 ;
        RECT 4.400 551.800 896.000 552.480 ;
        RECT 4.000 548.440 896.000 551.800 ;
        RECT 4.400 547.040 895.600 548.440 ;
        RECT 4.000 543.680 896.000 547.040 ;
        RECT 4.400 542.320 896.000 543.680 ;
        RECT 4.400 542.280 895.600 542.320 ;
        RECT 4.000 540.920 895.600 542.280 ;
        RECT 4.000 538.920 896.000 540.920 ;
        RECT 4.400 537.520 896.000 538.920 ;
        RECT 4.000 536.880 896.000 537.520 ;
        RECT 4.000 535.480 895.600 536.880 ;
        RECT 4.000 533.480 896.000 535.480 ;
        RECT 4.400 532.080 896.000 533.480 ;
        RECT 4.000 531.440 896.000 532.080 ;
        RECT 4.000 530.040 895.600 531.440 ;
        RECT 4.000 528.720 896.000 530.040 ;
        RECT 4.400 527.320 896.000 528.720 ;
        RECT 4.000 526.000 896.000 527.320 ;
        RECT 4.000 524.600 895.600 526.000 ;
        RECT 4.000 523.960 896.000 524.600 ;
        RECT 4.400 522.560 896.000 523.960 ;
        RECT 4.000 520.560 896.000 522.560 ;
        RECT 4.000 519.200 895.600 520.560 ;
        RECT 4.400 519.160 895.600 519.200 ;
        RECT 4.400 517.800 896.000 519.160 ;
        RECT 4.000 515.120 896.000 517.800 ;
        RECT 4.000 513.760 895.600 515.120 ;
        RECT 4.400 513.720 895.600 513.760 ;
        RECT 4.400 512.360 896.000 513.720 ;
        RECT 4.000 509.680 896.000 512.360 ;
        RECT 4.000 509.000 895.600 509.680 ;
        RECT 4.400 508.280 895.600 509.000 ;
        RECT 4.400 507.600 896.000 508.280 ;
        RECT 4.000 504.240 896.000 507.600 ;
        RECT 4.400 502.840 895.600 504.240 ;
        RECT 4.000 499.480 896.000 502.840 ;
        RECT 4.400 498.800 896.000 499.480 ;
        RECT 4.400 498.080 895.600 498.800 ;
        RECT 4.000 497.400 895.600 498.080 ;
        RECT 4.000 494.040 896.000 497.400 ;
        RECT 4.400 493.360 896.000 494.040 ;
        RECT 4.400 492.640 895.600 493.360 ;
        RECT 4.000 491.960 895.600 492.640 ;
        RECT 4.000 489.280 896.000 491.960 ;
        RECT 4.400 487.920 896.000 489.280 ;
        RECT 4.400 487.880 895.600 487.920 ;
        RECT 4.000 486.520 895.600 487.880 ;
        RECT 4.000 484.520 896.000 486.520 ;
        RECT 4.400 483.120 896.000 484.520 ;
        RECT 4.000 481.800 896.000 483.120 ;
        RECT 4.000 480.400 895.600 481.800 ;
        RECT 4.000 479.760 896.000 480.400 ;
        RECT 4.400 478.360 896.000 479.760 ;
        RECT 4.000 476.360 896.000 478.360 ;
        RECT 4.000 475.000 895.600 476.360 ;
        RECT 4.400 474.960 895.600 475.000 ;
        RECT 4.400 473.600 896.000 474.960 ;
        RECT 4.000 470.920 896.000 473.600 ;
        RECT 4.000 469.560 895.600 470.920 ;
        RECT 4.400 469.520 895.600 469.560 ;
        RECT 4.400 468.160 896.000 469.520 ;
        RECT 4.000 465.480 896.000 468.160 ;
        RECT 4.000 464.800 895.600 465.480 ;
        RECT 4.400 464.080 895.600 464.800 ;
        RECT 4.400 463.400 896.000 464.080 ;
        RECT 4.000 460.040 896.000 463.400 ;
        RECT 4.400 458.640 895.600 460.040 ;
        RECT 4.000 455.280 896.000 458.640 ;
        RECT 4.400 454.600 896.000 455.280 ;
        RECT 4.400 453.880 895.600 454.600 ;
        RECT 4.000 453.200 895.600 453.880 ;
        RECT 4.000 449.840 896.000 453.200 ;
        RECT 4.400 449.160 896.000 449.840 ;
        RECT 4.400 448.440 895.600 449.160 ;
        RECT 4.000 447.760 895.600 448.440 ;
        RECT 4.000 445.080 896.000 447.760 ;
        RECT 4.400 443.720 896.000 445.080 ;
        RECT 4.400 443.680 895.600 443.720 ;
        RECT 4.000 442.320 895.600 443.680 ;
        RECT 4.000 440.320 896.000 442.320 ;
        RECT 4.400 438.920 896.000 440.320 ;
        RECT 4.000 438.280 896.000 438.920 ;
        RECT 4.000 436.880 895.600 438.280 ;
        RECT 4.000 435.560 896.000 436.880 ;
        RECT 4.400 434.160 896.000 435.560 ;
        RECT 4.000 432.840 896.000 434.160 ;
        RECT 4.000 431.440 895.600 432.840 ;
        RECT 4.000 430.120 896.000 431.440 ;
        RECT 4.400 428.720 896.000 430.120 ;
        RECT 4.000 427.400 896.000 428.720 ;
        RECT 4.000 426.000 895.600 427.400 ;
        RECT 4.000 425.360 896.000 426.000 ;
        RECT 4.400 423.960 896.000 425.360 ;
        RECT 4.000 421.280 896.000 423.960 ;
        RECT 4.000 420.600 895.600 421.280 ;
        RECT 4.400 419.880 895.600 420.600 ;
        RECT 4.400 419.200 896.000 419.880 ;
        RECT 4.000 415.840 896.000 419.200 ;
        RECT 4.400 414.440 895.600 415.840 ;
        RECT 4.000 411.080 896.000 414.440 ;
        RECT 4.400 410.400 896.000 411.080 ;
        RECT 4.400 409.680 895.600 410.400 ;
        RECT 4.000 409.000 895.600 409.680 ;
        RECT 4.000 405.640 896.000 409.000 ;
        RECT 4.400 404.960 896.000 405.640 ;
        RECT 4.400 404.240 895.600 404.960 ;
        RECT 4.000 403.560 895.600 404.240 ;
        RECT 4.000 400.880 896.000 403.560 ;
        RECT 4.400 399.520 896.000 400.880 ;
        RECT 4.400 399.480 895.600 399.520 ;
        RECT 4.000 398.120 895.600 399.480 ;
        RECT 4.000 396.120 896.000 398.120 ;
        RECT 4.400 394.720 896.000 396.120 ;
        RECT 4.000 394.080 896.000 394.720 ;
        RECT 4.000 392.680 895.600 394.080 ;
        RECT 4.000 391.360 896.000 392.680 ;
        RECT 4.400 389.960 896.000 391.360 ;
        RECT 4.000 388.640 896.000 389.960 ;
        RECT 4.000 387.240 895.600 388.640 ;
        RECT 4.000 385.920 896.000 387.240 ;
        RECT 4.400 384.520 896.000 385.920 ;
        RECT 4.000 383.200 896.000 384.520 ;
        RECT 4.000 381.800 895.600 383.200 ;
        RECT 4.000 381.160 896.000 381.800 ;
        RECT 4.400 379.760 896.000 381.160 ;
        RECT 4.000 377.760 896.000 379.760 ;
        RECT 4.000 376.400 895.600 377.760 ;
        RECT 4.400 376.360 895.600 376.400 ;
        RECT 4.400 375.000 896.000 376.360 ;
        RECT 4.000 372.320 896.000 375.000 ;
        RECT 4.000 371.640 895.600 372.320 ;
        RECT 4.400 370.920 895.600 371.640 ;
        RECT 4.400 370.240 896.000 370.920 ;
        RECT 4.000 366.880 896.000 370.240 ;
        RECT 4.000 366.200 895.600 366.880 ;
        RECT 4.400 365.480 895.600 366.200 ;
        RECT 4.400 364.800 896.000 365.480 ;
        RECT 4.000 361.440 896.000 364.800 ;
        RECT 4.400 360.760 896.000 361.440 ;
        RECT 4.400 360.040 895.600 360.760 ;
        RECT 4.000 359.360 895.600 360.040 ;
        RECT 4.000 356.680 896.000 359.360 ;
        RECT 4.400 355.320 896.000 356.680 ;
        RECT 4.400 355.280 895.600 355.320 ;
        RECT 4.000 353.920 895.600 355.280 ;
        RECT 4.000 351.920 896.000 353.920 ;
        RECT 4.400 350.520 896.000 351.920 ;
        RECT 4.000 349.880 896.000 350.520 ;
        RECT 4.000 348.480 895.600 349.880 ;
        RECT 4.000 347.160 896.000 348.480 ;
        RECT 4.400 345.760 896.000 347.160 ;
        RECT 4.000 344.440 896.000 345.760 ;
        RECT 4.000 343.040 895.600 344.440 ;
        RECT 4.000 341.720 896.000 343.040 ;
        RECT 4.400 340.320 896.000 341.720 ;
        RECT 4.000 339.000 896.000 340.320 ;
        RECT 4.000 337.600 895.600 339.000 ;
        RECT 4.000 336.960 896.000 337.600 ;
        RECT 4.400 335.560 896.000 336.960 ;
        RECT 4.000 333.560 896.000 335.560 ;
        RECT 4.000 332.200 895.600 333.560 ;
        RECT 4.400 332.160 895.600 332.200 ;
        RECT 4.400 330.800 896.000 332.160 ;
        RECT 4.000 328.120 896.000 330.800 ;
        RECT 4.000 327.440 895.600 328.120 ;
        RECT 4.400 326.720 895.600 327.440 ;
        RECT 4.400 326.040 896.000 326.720 ;
        RECT 4.000 322.680 896.000 326.040 ;
        RECT 4.000 322.000 895.600 322.680 ;
        RECT 4.400 321.280 895.600 322.000 ;
        RECT 4.400 320.600 896.000 321.280 ;
        RECT 4.000 317.240 896.000 320.600 ;
        RECT 4.400 315.840 895.600 317.240 ;
        RECT 4.000 312.480 896.000 315.840 ;
        RECT 4.400 311.800 896.000 312.480 ;
        RECT 4.400 311.080 895.600 311.800 ;
        RECT 4.000 310.400 895.600 311.080 ;
        RECT 4.000 307.720 896.000 310.400 ;
        RECT 4.400 306.360 896.000 307.720 ;
        RECT 4.400 306.320 895.600 306.360 ;
        RECT 4.000 304.960 895.600 306.320 ;
        RECT 4.000 302.960 896.000 304.960 ;
        RECT 4.400 301.560 896.000 302.960 ;
        RECT 4.000 300.240 896.000 301.560 ;
        RECT 4.000 298.840 895.600 300.240 ;
        RECT 4.000 297.520 896.000 298.840 ;
        RECT 4.400 296.120 896.000 297.520 ;
        RECT 4.000 294.800 896.000 296.120 ;
        RECT 4.000 293.400 895.600 294.800 ;
        RECT 4.000 292.760 896.000 293.400 ;
        RECT 4.400 291.360 896.000 292.760 ;
        RECT 4.000 289.360 896.000 291.360 ;
        RECT 4.000 288.000 895.600 289.360 ;
        RECT 4.400 287.960 895.600 288.000 ;
        RECT 4.400 286.600 896.000 287.960 ;
        RECT 4.000 283.920 896.000 286.600 ;
        RECT 4.000 283.240 895.600 283.920 ;
        RECT 4.400 282.520 895.600 283.240 ;
        RECT 4.400 281.840 896.000 282.520 ;
        RECT 4.000 278.480 896.000 281.840 ;
        RECT 4.000 277.800 895.600 278.480 ;
        RECT 4.400 277.080 895.600 277.800 ;
        RECT 4.400 276.400 896.000 277.080 ;
        RECT 4.000 273.040 896.000 276.400 ;
        RECT 4.400 271.640 895.600 273.040 ;
        RECT 4.000 268.280 896.000 271.640 ;
        RECT 4.400 267.600 896.000 268.280 ;
        RECT 4.400 266.880 895.600 267.600 ;
        RECT 4.000 266.200 895.600 266.880 ;
        RECT 4.000 263.520 896.000 266.200 ;
        RECT 4.400 262.160 896.000 263.520 ;
        RECT 4.400 262.120 895.600 262.160 ;
        RECT 4.000 260.760 895.600 262.120 ;
        RECT 4.000 258.080 896.000 260.760 ;
        RECT 4.400 256.720 896.000 258.080 ;
        RECT 4.400 256.680 895.600 256.720 ;
        RECT 4.000 255.320 895.600 256.680 ;
        RECT 4.000 253.320 896.000 255.320 ;
        RECT 4.400 251.920 896.000 253.320 ;
        RECT 4.000 251.280 896.000 251.920 ;
        RECT 4.000 249.880 895.600 251.280 ;
        RECT 4.000 248.560 896.000 249.880 ;
        RECT 4.400 247.160 896.000 248.560 ;
        RECT 4.000 245.840 896.000 247.160 ;
        RECT 4.000 244.440 895.600 245.840 ;
        RECT 4.000 243.800 896.000 244.440 ;
        RECT 4.400 242.400 896.000 243.800 ;
        RECT 4.000 239.720 896.000 242.400 ;
        RECT 4.000 239.040 895.600 239.720 ;
        RECT 4.400 238.320 895.600 239.040 ;
        RECT 4.400 237.640 896.000 238.320 ;
        RECT 4.000 234.280 896.000 237.640 ;
        RECT 4.000 233.600 895.600 234.280 ;
        RECT 4.400 232.880 895.600 233.600 ;
        RECT 4.400 232.200 896.000 232.880 ;
        RECT 4.000 228.840 896.000 232.200 ;
        RECT 4.400 227.440 895.600 228.840 ;
        RECT 4.000 224.080 896.000 227.440 ;
        RECT 4.400 223.400 896.000 224.080 ;
        RECT 4.400 222.680 895.600 223.400 ;
        RECT 4.000 222.000 895.600 222.680 ;
        RECT 4.000 219.320 896.000 222.000 ;
        RECT 4.400 217.960 896.000 219.320 ;
        RECT 4.400 217.920 895.600 217.960 ;
        RECT 4.000 216.560 895.600 217.920 ;
        RECT 4.000 213.880 896.000 216.560 ;
        RECT 4.400 212.520 896.000 213.880 ;
        RECT 4.400 212.480 895.600 212.520 ;
        RECT 4.000 211.120 895.600 212.480 ;
        RECT 4.000 209.120 896.000 211.120 ;
        RECT 4.400 207.720 896.000 209.120 ;
        RECT 4.000 207.080 896.000 207.720 ;
        RECT 4.000 205.680 895.600 207.080 ;
        RECT 4.000 204.360 896.000 205.680 ;
        RECT 4.400 202.960 896.000 204.360 ;
        RECT 4.000 201.640 896.000 202.960 ;
        RECT 4.000 200.240 895.600 201.640 ;
        RECT 4.000 199.600 896.000 200.240 ;
        RECT 4.400 198.200 896.000 199.600 ;
        RECT 4.000 196.200 896.000 198.200 ;
        RECT 4.000 194.800 895.600 196.200 ;
        RECT 4.000 194.160 896.000 194.800 ;
        RECT 4.400 192.760 896.000 194.160 ;
        RECT 4.000 190.760 896.000 192.760 ;
        RECT 4.000 189.400 895.600 190.760 ;
        RECT 4.400 189.360 895.600 189.400 ;
        RECT 4.400 188.000 896.000 189.360 ;
        RECT 4.000 185.320 896.000 188.000 ;
        RECT 4.000 184.640 895.600 185.320 ;
        RECT 4.400 183.920 895.600 184.640 ;
        RECT 4.400 183.240 896.000 183.920 ;
        RECT 4.000 179.880 896.000 183.240 ;
        RECT 4.400 179.200 896.000 179.880 ;
        RECT 4.400 178.480 895.600 179.200 ;
        RECT 4.000 177.800 895.600 178.480 ;
        RECT 4.000 175.120 896.000 177.800 ;
        RECT 4.400 173.760 896.000 175.120 ;
        RECT 4.400 173.720 895.600 173.760 ;
        RECT 4.000 172.360 895.600 173.720 ;
        RECT 4.000 169.680 896.000 172.360 ;
        RECT 4.400 168.320 896.000 169.680 ;
        RECT 4.400 168.280 895.600 168.320 ;
        RECT 4.000 166.920 895.600 168.280 ;
        RECT 4.000 164.920 896.000 166.920 ;
        RECT 4.400 163.520 896.000 164.920 ;
        RECT 4.000 162.880 896.000 163.520 ;
        RECT 4.000 161.480 895.600 162.880 ;
        RECT 4.000 160.160 896.000 161.480 ;
        RECT 4.400 158.760 896.000 160.160 ;
        RECT 4.000 157.440 896.000 158.760 ;
        RECT 4.000 156.040 895.600 157.440 ;
        RECT 4.000 155.400 896.000 156.040 ;
        RECT 4.400 154.000 896.000 155.400 ;
        RECT 4.000 152.000 896.000 154.000 ;
        RECT 4.000 150.600 895.600 152.000 ;
        RECT 4.000 149.960 896.000 150.600 ;
        RECT 4.400 148.560 896.000 149.960 ;
        RECT 4.000 146.560 896.000 148.560 ;
        RECT 4.000 145.200 895.600 146.560 ;
        RECT 4.400 145.160 895.600 145.200 ;
        RECT 4.400 143.800 896.000 145.160 ;
        RECT 4.000 141.120 896.000 143.800 ;
        RECT 4.000 140.440 895.600 141.120 ;
        RECT 4.400 139.720 895.600 140.440 ;
        RECT 4.400 139.040 896.000 139.720 ;
        RECT 4.000 135.680 896.000 139.040 ;
        RECT 4.400 134.280 895.600 135.680 ;
        RECT 4.000 130.240 896.000 134.280 ;
        RECT 4.400 128.840 895.600 130.240 ;
        RECT 4.000 125.480 896.000 128.840 ;
        RECT 4.400 124.800 896.000 125.480 ;
        RECT 4.400 124.080 895.600 124.800 ;
        RECT 4.000 123.400 895.600 124.080 ;
        RECT 4.000 120.720 896.000 123.400 ;
        RECT 4.400 119.320 896.000 120.720 ;
        RECT 4.000 118.680 896.000 119.320 ;
        RECT 4.000 117.280 895.600 118.680 ;
        RECT 4.000 115.960 896.000 117.280 ;
        RECT 4.400 114.560 896.000 115.960 ;
        RECT 4.000 113.240 896.000 114.560 ;
        RECT 4.000 111.840 895.600 113.240 ;
        RECT 4.000 111.200 896.000 111.840 ;
        RECT 4.400 109.800 896.000 111.200 ;
        RECT 4.000 107.800 896.000 109.800 ;
        RECT 4.000 106.400 895.600 107.800 ;
        RECT 4.000 105.760 896.000 106.400 ;
        RECT 4.400 104.360 896.000 105.760 ;
        RECT 4.000 102.360 896.000 104.360 ;
        RECT 4.000 101.000 895.600 102.360 ;
        RECT 4.400 100.960 895.600 101.000 ;
        RECT 4.400 99.600 896.000 100.960 ;
        RECT 4.000 96.920 896.000 99.600 ;
        RECT 4.000 96.240 895.600 96.920 ;
        RECT 4.400 95.520 895.600 96.240 ;
        RECT 4.400 94.840 896.000 95.520 ;
        RECT 4.000 91.480 896.000 94.840 ;
        RECT 4.400 90.080 895.600 91.480 ;
        RECT 4.000 86.040 896.000 90.080 ;
        RECT 4.400 84.640 895.600 86.040 ;
        RECT 4.000 81.280 896.000 84.640 ;
        RECT 4.400 80.600 896.000 81.280 ;
        RECT 4.400 79.880 895.600 80.600 ;
        RECT 4.000 79.200 895.600 79.880 ;
        RECT 4.000 76.520 896.000 79.200 ;
        RECT 4.400 75.160 896.000 76.520 ;
        RECT 4.400 75.120 895.600 75.160 ;
        RECT 4.000 73.760 895.600 75.120 ;
        RECT 4.000 71.760 896.000 73.760 ;
        RECT 4.400 70.360 896.000 71.760 ;
        RECT 4.000 69.720 896.000 70.360 ;
        RECT 4.000 68.320 895.600 69.720 ;
        RECT 4.000 66.320 896.000 68.320 ;
        RECT 4.400 64.920 896.000 66.320 ;
        RECT 4.000 64.280 896.000 64.920 ;
        RECT 4.000 62.880 895.600 64.280 ;
        RECT 4.000 61.560 896.000 62.880 ;
        RECT 4.400 60.160 896.000 61.560 ;
        RECT 4.000 58.160 896.000 60.160 ;
        RECT 4.000 56.800 895.600 58.160 ;
        RECT 4.400 56.760 895.600 56.800 ;
        RECT 4.400 55.400 896.000 56.760 ;
        RECT 4.000 52.720 896.000 55.400 ;
        RECT 4.000 52.040 895.600 52.720 ;
        RECT 4.400 51.320 895.600 52.040 ;
        RECT 4.400 50.640 896.000 51.320 ;
        RECT 4.000 47.280 896.000 50.640 ;
        RECT 4.400 45.880 895.600 47.280 ;
        RECT 4.000 41.840 896.000 45.880 ;
        RECT 4.400 40.440 895.600 41.840 ;
        RECT 4.000 37.080 896.000 40.440 ;
        RECT 4.400 36.400 896.000 37.080 ;
        RECT 4.400 35.680 895.600 36.400 ;
        RECT 4.000 35.000 895.600 35.680 ;
        RECT 4.000 32.320 896.000 35.000 ;
        RECT 4.400 30.960 896.000 32.320 ;
        RECT 4.400 30.920 895.600 30.960 ;
        RECT 4.000 29.560 895.600 30.920 ;
        RECT 4.000 27.560 896.000 29.560 ;
        RECT 4.400 26.160 896.000 27.560 ;
        RECT 4.000 25.520 896.000 26.160 ;
        RECT 4.000 24.120 895.600 25.520 ;
        RECT 4.000 22.120 896.000 24.120 ;
        RECT 4.400 20.720 896.000 22.120 ;
        RECT 4.000 20.080 896.000 20.720 ;
        RECT 4.000 18.680 895.600 20.080 ;
        RECT 4.000 17.360 896.000 18.680 ;
        RECT 4.400 15.960 896.000 17.360 ;
        RECT 4.000 14.640 896.000 15.960 ;
        RECT 4.000 13.240 895.600 14.640 ;
        RECT 4.000 12.600 896.000 13.240 ;
        RECT 4.400 11.200 896.000 12.600 ;
        RECT 4.000 9.200 896.000 11.200 ;
        RECT 4.000 7.840 895.600 9.200 ;
        RECT 4.400 7.800 895.600 7.840 ;
        RECT 4.400 6.440 896.000 7.800 ;
        RECT 4.000 3.760 896.000 6.440 ;
        RECT 4.000 3.080 895.600 3.760 ;
        RECT 4.400 2.360 895.600 3.080 ;
        RECT 4.400 2.215 896.000 2.360 ;
  END
END vco_adc_wrapper
END LIBRARY

