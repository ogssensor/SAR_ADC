VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_adc_wrapper
  CLASS BLOCK ;
  FOREIGN vco_adc_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 800.000 ;
  PIN adc0_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 3.440 900.000 4.040 ;
    END
  END adc0_dat_i[0]
  PIN adc0_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 245.520 900.000 246.120 ;
    END
  END adc0_dat_i[10]
  PIN adc0_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 267.280 900.000 267.880 ;
    END
  END adc0_dat_i[11]
  PIN adc0_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 289.040 900.000 289.640 ;
    END
  END adc0_dat_i[12]
  PIN adc0_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 311.480 900.000 312.080 ;
    END
  END adc0_dat_i[13]
  PIN adc0_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 333.240 900.000 333.840 ;
    END
  END adc0_dat_i[14]
  PIN adc0_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 355.000 900.000 355.600 ;
    END
  END adc0_dat_i[15]
  PIN adc0_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 377.440 900.000 378.040 ;
    END
  END adc0_dat_i[16]
  PIN adc0_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 399.200 900.000 399.800 ;
    END
  END adc0_dat_i[17]
  PIN adc0_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 420.960 900.000 421.560 ;
    END
  END adc0_dat_i[18]
  PIN adc0_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 443.400 900.000 444.000 ;
    END
  END adc0_dat_i[19]
  PIN adc0_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 32.680 900.000 33.280 ;
    END
  END adc0_dat_i[1]
  PIN adc0_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 465.160 900.000 465.760 ;
    END
  END adc0_dat_i[20]
  PIN adc0_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 487.600 900.000 488.200 ;
    END
  END adc0_dat_i[21]
  PIN adc0_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 509.360 900.000 509.960 ;
    END
  END adc0_dat_i[22]
  PIN adc0_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 531.120 900.000 531.720 ;
    END
  END adc0_dat_i[23]
  PIN adc0_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 553.560 900.000 554.160 ;
    END
  END adc0_dat_i[24]
  PIN adc0_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 575.320 900.000 575.920 ;
    END
  END adc0_dat_i[25]
  PIN adc0_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 597.080 900.000 597.680 ;
    END
  END adc0_dat_i[26]
  PIN adc0_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 619.520 900.000 620.120 ;
    END
  END adc0_dat_i[27]
  PIN adc0_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 641.280 900.000 641.880 ;
    END
  END adc0_dat_i[28]
  PIN adc0_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 663.720 900.000 664.320 ;
    END
  END adc0_dat_i[29]
  PIN adc0_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 61.920 900.000 62.520 ;
    END
  END adc0_dat_i[2]
  PIN adc0_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 685.480 900.000 686.080 ;
    END
  END adc0_dat_i[30]
  PIN adc0_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 707.240 900.000 707.840 ;
    END
  END adc0_dat_i[31]
  PIN adc0_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 91.160 900.000 91.760 ;
    END
  END adc0_dat_i[3]
  PIN adc0_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 112.920 900.000 113.520 ;
    END
  END adc0_dat_i[4]
  PIN adc0_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 135.360 900.000 135.960 ;
    END
  END adc0_dat_i[5]
  PIN adc0_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 157.120 900.000 157.720 ;
    END
  END adc0_dat_i[6]
  PIN adc0_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 178.880 900.000 179.480 ;
    END
  END adc0_dat_i[7]
  PIN adc0_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 201.320 900.000 201.920 ;
    END
  END adc0_dat_i[8]
  PIN adc0_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 223.080 900.000 223.680 ;
    END
  END adc0_dat_i[9]
  PIN adc1_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 10.240 900.000 10.840 ;
    END
  END adc1_dat_i[0]
  PIN adc1_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 252.320 900.000 252.920 ;
    END
  END adc1_dat_i[10]
  PIN adc1_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 274.760 900.000 275.360 ;
    END
  END adc1_dat_i[11]
  PIN adc1_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 296.520 900.000 297.120 ;
    END
  END adc1_dat_i[12]
  PIN adc1_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 318.280 900.000 318.880 ;
    END
  END adc1_dat_i[13]
  PIN adc1_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 340.720 900.000 341.320 ;
    END
  END adc1_dat_i[14]
  PIN adc1_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 362.480 900.000 363.080 ;
    END
  END adc1_dat_i[15]
  PIN adc1_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 384.920 900.000 385.520 ;
    END
  END adc1_dat_i[16]
  PIN adc1_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 406.680 900.000 407.280 ;
    END
  END adc1_dat_i[17]
  PIN adc1_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 428.440 900.000 429.040 ;
    END
  END adc1_dat_i[18]
  PIN adc1_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 450.880 900.000 451.480 ;
    END
  END adc1_dat_i[19]
  PIN adc1_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 39.480 900.000 40.080 ;
    END
  END adc1_dat_i[1]
  PIN adc1_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 472.640 900.000 473.240 ;
    END
  END adc1_dat_i[20]
  PIN adc1_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 494.400 900.000 495.000 ;
    END
  END adc1_dat_i[21]
  PIN adc1_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 516.840 900.000 517.440 ;
    END
  END adc1_dat_i[22]
  PIN adc1_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 538.600 900.000 539.200 ;
    END
  END adc1_dat_i[23]
  PIN adc1_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 560.360 900.000 560.960 ;
    END
  END adc1_dat_i[24]
  PIN adc1_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 582.800 900.000 583.400 ;
    END
  END adc1_dat_i[25]
  PIN adc1_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 604.560 900.000 605.160 ;
    END
  END adc1_dat_i[26]
  PIN adc1_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 627.000 900.000 627.600 ;
    END
  END adc1_dat_i[27]
  PIN adc1_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 648.760 900.000 649.360 ;
    END
  END adc1_dat_i[28]
  PIN adc1_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 670.520 900.000 671.120 ;
    END
  END adc1_dat_i[29]
  PIN adc1_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 69.400 900.000 70.000 ;
    END
  END adc1_dat_i[2]
  PIN adc1_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 692.960 900.000 693.560 ;
    END
  END adc1_dat_i[30]
  PIN adc1_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 714.720 900.000 715.320 ;
    END
  END adc1_dat_i[31]
  PIN adc1_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 98.640 900.000 99.240 ;
    END
  END adc1_dat_i[3]
  PIN adc1_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 120.400 900.000 121.000 ;
    END
  END adc1_dat_i[4]
  PIN adc1_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 142.160 900.000 142.760 ;
    END
  END adc1_dat_i[5]
  PIN adc1_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 164.600 900.000 165.200 ;
    END
  END adc1_dat_i[6]
  PIN adc1_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 186.360 900.000 186.960 ;
    END
  END adc1_dat_i[7]
  PIN adc1_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 208.800 900.000 209.400 ;
    END
  END adc1_dat_i[8]
  PIN adc1_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 230.560 900.000 231.160 ;
    END
  END adc1_dat_i[9]
  PIN adc2_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 17.720 900.000 18.320 ;
    END
  END adc2_dat_i[0]
  PIN adc2_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 259.800 900.000 260.400 ;
    END
  END adc2_dat_i[10]
  PIN adc2_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 281.560 900.000 282.160 ;
    END
  END adc2_dat_i[11]
  PIN adc2_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 304.000 900.000 304.600 ;
    END
  END adc2_dat_i[12]
  PIN adc2_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 325.760 900.000 326.360 ;
    END
  END adc2_dat_i[13]
  PIN adc2_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 348.200 900.000 348.800 ;
    END
  END adc2_dat_i[14]
  PIN adc2_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 369.960 900.000 370.560 ;
    END
  END adc2_dat_i[15]
  PIN adc2_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 391.720 900.000 392.320 ;
    END
  END adc2_dat_i[16]
  PIN adc2_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 414.160 900.000 414.760 ;
    END
  END adc2_dat_i[17]
  PIN adc2_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 435.920 900.000 436.520 ;
    END
  END adc2_dat_i[18]
  PIN adc2_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 457.680 900.000 458.280 ;
    END
  END adc2_dat_i[19]
  PIN adc2_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 46.960 900.000 47.560 ;
    END
  END adc2_dat_i[1]
  PIN adc2_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 480.120 900.000 480.720 ;
    END
  END adc2_dat_i[20]
  PIN adc2_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 501.880 900.000 502.480 ;
    END
  END adc2_dat_i[21]
  PIN adc2_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 524.320 900.000 524.920 ;
    END
  END adc2_dat_i[22]
  PIN adc2_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 546.080 900.000 546.680 ;
    END
  END adc2_dat_i[23]
  PIN adc2_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 567.840 900.000 568.440 ;
    END
  END adc2_dat_i[24]
  PIN adc2_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 590.280 900.000 590.880 ;
    END
  END adc2_dat_i[25]
  PIN adc2_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 612.040 900.000 612.640 ;
    END
  END adc2_dat_i[26]
  PIN adc2_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 633.800 900.000 634.400 ;
    END
  END adc2_dat_i[27]
  PIN adc2_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 656.240 900.000 656.840 ;
    END
  END adc2_dat_i[28]
  PIN adc2_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 678.000 900.000 678.600 ;
    END
  END adc2_dat_i[29]
  PIN adc2_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 76.200 900.000 76.800 ;
    END
  END adc2_dat_i[2]
  PIN adc2_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 699.760 900.000 700.360 ;
    END
  END adc2_dat_i[30]
  PIN adc2_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 722.200 900.000 722.800 ;
    END
  END adc2_dat_i[31]
  PIN adc2_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 106.120 900.000 106.720 ;
    END
  END adc2_dat_i[3]
  PIN adc2_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 127.880 900.000 128.480 ;
    END
  END adc2_dat_i[4]
  PIN adc2_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 149.640 900.000 150.240 ;
    END
  END adc2_dat_i[5]
  PIN adc2_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 172.080 900.000 172.680 ;
    END
  END adc2_dat_i[6]
  PIN adc2_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 193.840 900.000 194.440 ;
    END
  END adc2_dat_i[7]
  PIN adc2_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 215.600 900.000 216.200 ;
    END
  END adc2_dat_i[8]
  PIN adc2_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 238.040 900.000 238.640 ;
    END
  END adc2_dat_i[9]
  PIN adc_dvalid_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 25.200 900.000 25.800 ;
    END
  END adc_dvalid_i[0]
  PIN adc_dvalid_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 54.440 900.000 55.040 ;
    END
  END adc_dvalid_i[1]
  PIN adc_dvalid_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 83.680 900.000 84.280 ;
    END
  END adc_dvalid_i[2]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 796.000 5.430 800.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 796.000 224.850 800.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 796.000 246.930 800.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 796.000 268.550 800.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 796.000 290.630 800.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 796.000 312.710 800.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 796.000 334.330 800.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 796.000 356.410 800.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 796.000 378.490 800.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 796.000 400.570 800.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 796.000 422.190 800.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 796.000 27.050 800.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 796.000 444.270 800.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 796.000 466.350 800.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 796.000 488.430 800.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 796.000 510.050 800.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 796.000 532.130 800.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 796.000 554.210 800.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 796.000 576.290 800.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 796.000 597.910 800.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 796.000 619.990 800.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 796.000 642.070 800.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 796.000 49.130 800.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 796.000 663.690 800.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 796.000 685.770 800.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 796.000 707.850 800.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 796.000 729.930 800.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 796.000 751.550 800.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 796.000 773.630 800.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 796.000 795.710 800.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 796.000 817.790 800.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 796.000 71.210 800.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 796.000 92.830 800.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 796.000 114.910 800.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 796.000 136.990 800.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 796.000 159.070 800.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 796.000 180.690 800.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 796.000 202.770 800.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 796.000 16.010 800.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 796.000 235.890 800.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 796.000 257.510 800.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 796.000 279.590 800.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 796.000 301.670 800.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 796.000 323.750 800.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 796.000 345.370 800.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 796.000 367.450 800.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 796.000 389.530 800.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 796.000 411.610 800.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 796.000 433.230 800.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 796.000 38.090 800.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 796.000 455.310 800.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 796.000 477.390 800.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 796.000 499.010 800.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 796.000 521.090 800.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 796.000 543.170 800.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 796.000 565.250 800.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 796.000 586.870 800.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 796.000 608.950 800.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 796.000 631.030 800.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 796.000 653.110 800.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 796.000 60.170 800.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 796.000 674.730 800.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 796.000 696.810 800.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 796.000 718.890 800.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 796.000 740.970 800.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 796.000 762.590 800.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 796.000 784.670 800.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 796.000 806.750 800.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 796.000 828.370 800.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 796.000 82.250 800.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 796.000 103.870 800.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 796.000 125.950 800.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 796.000 148.030 800.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 796.000 169.650 800.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 796.000 191.730 800.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 796.000 213.810 800.000 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.150 0.000 879.430 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END irq[2]
  PIN mem1_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 28.600 4.000 29.200 ;
    END
  END mem1_data_i[0]
  PIN mem1_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END mem1_data_i[10]
  PIN mem1_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.000 4.000 389.600 ;
    END
  END mem1_data_i[11]
  PIN mem1_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END mem1_data_i[12]
  PIN mem1_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END mem1_data_i[13]
  PIN mem1_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END mem1_data_i[14]
  PIN mem1_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.880 4.000 468.480 ;
    END
  END mem1_data_i[15]
  PIN mem1_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END mem1_data_i[16]
  PIN mem1_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END mem1_data_i[17]
  PIN mem1_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.040 4.000 527.640 ;
    END
  END mem1_data_i[18]
  PIN mem1_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END mem1_data_i[19]
  PIN mem1_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END mem1_data_i[1]
  PIN mem1_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END mem1_data_i[20]
  PIN mem1_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END mem1_data_i[21]
  PIN mem1_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 605.240 4.000 605.840 ;
    END
  END mem1_data_i[22]
  PIN mem1_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 624.960 4.000 625.560 ;
    END
  END mem1_data_i[23]
  PIN mem1_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END mem1_data_i[24]
  PIN mem1_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 664.400 4.000 665.000 ;
    END
  END mem1_data_i[25]
  PIN mem1_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.120 4.000 684.720 ;
    END
  END mem1_data_i[26]
  PIN mem1_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 703.840 4.000 704.440 ;
    END
  END mem1_data_i[27]
  PIN mem1_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 723.560 4.000 724.160 ;
    END
  END mem1_data_i[28]
  PIN mem1_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END mem1_data_i[29]
  PIN mem1_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 120.400 4.000 121.000 ;
    END
  END mem1_data_i[2]
  PIN mem1_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 763.000 4.000 763.600 ;
    END
  END mem1_data_i[30]
  PIN mem1_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 782.720 4.000 783.320 ;
    END
  END mem1_data_i[31]
  PIN mem1_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END mem1_data_i[3]
  PIN mem1_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END mem1_data_i[4]
  PIN mem1_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END mem1_data_i[5]
  PIN mem1_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END mem1_data_i[6]
  PIN mem1_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 284.280 4.000 284.880 ;
    END
  END mem1_data_i[7]
  PIN mem1_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END mem1_data_i[8]
  PIN mem1_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END mem1_data_i[9]
  PIN mem_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END mem_data_i[0]
  PIN mem_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.080 4.000 376.680 ;
    END
  END mem_data_i[10]
  PIN mem_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END mem_data_i[11]
  PIN mem_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END mem_data_i[12]
  PIN mem_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END mem_data_i[13]
  PIN mem_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END mem_data_i[14]
  PIN mem_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.680 4.000 475.280 ;
    END
  END mem_data_i[15]
  PIN mem_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.720 4.000 494.320 ;
    END
  END mem_data_i[16]
  PIN mem_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 513.440 4.000 514.040 ;
    END
  END mem_data_i[17]
  PIN mem_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.160 4.000 533.760 ;
    END
  END mem_data_i[18]
  PIN mem_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END mem_data_i[19]
  PIN mem_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END mem_data_i[1]
  PIN mem_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END mem_data_i[20]
  PIN mem_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 592.320 4.000 592.920 ;
    END
  END mem_data_i[21]
  PIN mem_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 612.040 4.000 612.640 ;
    END
  END mem_data_i[22]
  PIN mem_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.760 4.000 632.360 ;
    END
  END mem_data_i[23]
  PIN mem_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 651.480 4.000 652.080 ;
    END
  END mem_data_i[24]
  PIN mem_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.200 4.000 671.800 ;
    END
  END mem_data_i[25]
  PIN mem_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END mem_data_i[26]
  PIN mem_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 710.640 4.000 711.240 ;
    END
  END mem_data_i[27]
  PIN mem_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 729.680 4.000 730.280 ;
    END
  END mem_data_i[28]
  PIN mem_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 749.400 4.000 750.000 ;
    END
  END mem_data_i[29]
  PIN mem_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.200 4.000 127.800 ;
    END
  END mem_data_i[2]
  PIN mem_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 769.120 4.000 769.720 ;
    END
  END mem_data_i[30]
  PIN mem_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.840 4.000 789.440 ;
    END
  END mem_data_i[31]
  PIN mem_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END mem_data_i[3]
  PIN mem_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 192.480 4.000 193.080 ;
    END
  END mem_data_i[4]
  PIN mem_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.120 4.000 225.720 ;
    END
  END mem_data_i[5]
  PIN mem_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END mem_data_i[6]
  PIN mem_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END mem_data_i[7]
  PIN mem_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END mem_data_i[8]
  PIN mem_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 356.360 4.000 356.960 ;
    END
  END mem_data_i[9]
  PIN mem_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 41.520 4.000 42.120 ;
    END
  END mem_data_o[0]
  PIN mem_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END mem_data_o[10]
  PIN mem_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END mem_data_o[11]
  PIN mem_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END mem_data_o[12]
  PIN mem_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END mem_data_o[13]
  PIN mem_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END mem_data_o[14]
  PIN mem_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END mem_data_o[15]
  PIN mem_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 500.520 4.000 501.120 ;
    END
  END mem_data_o[16]
  PIN mem_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.240 4.000 520.840 ;
    END
  END mem_data_o[17]
  PIN mem_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END mem_data_o[18]
  PIN mem_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END mem_data_o[19]
  PIN mem_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END mem_data_o[1]
  PIN mem_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 579.400 4.000 580.000 ;
    END
  END mem_data_o[20]
  PIN mem_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END mem_data_o[21]
  PIN mem_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 618.840 4.000 619.440 ;
    END
  END mem_data_o[22]
  PIN mem_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END mem_data_o[23]
  PIN mem_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 657.600 4.000 658.200 ;
    END
  END mem_data_o[24]
  PIN mem_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 677.320 4.000 677.920 ;
    END
  END mem_data_o[25]
  PIN mem_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.040 4.000 697.640 ;
    END
  END mem_data_o[26]
  PIN mem_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 716.760 4.000 717.360 ;
    END
  END mem_data_o[27]
  PIN mem_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 736.480 4.000 737.080 ;
    END
  END mem_data_o[28]
  PIN mem_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 756.200 4.000 756.800 ;
    END
  END mem_data_o[29]
  PIN mem_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END mem_data_o[2]
  PIN mem_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 775.920 4.000 776.520 ;
    END
  END mem_data_o[30]
  PIN mem_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END mem_data_o[31]
  PIN mem_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 165.960 4.000 166.560 ;
    END
  END mem_data_o[3]
  PIN mem_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.280 4.000 199.880 ;
    END
  END mem_data_o[4]
  PIN mem_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END mem_data_o[5]
  PIN mem_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END mem_data_o[6]
  PIN mem_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.200 4.000 297.800 ;
    END
  END mem_data_o[7]
  PIN mem_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.840 4.000 330.440 ;
    END
  END mem_data_o[8]
  PIN mem_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.160 4.000 363.760 ;
    END
  END mem_data_o[9]
  PIN mem_raddr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END mem_raddr_o[0]
  PIN mem_raddr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END mem_raddr_o[1]
  PIN mem_raddr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END mem_raddr_o[2]
  PIN mem_raddr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 172.760 4.000 173.360 ;
    END
  END mem_raddr_o[3]
  PIN mem_raddr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 205.400 4.000 206.000 ;
    END
  END mem_raddr_o[4]
  PIN mem_raddr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END mem_raddr_o[5]
  PIN mem_raddr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 271.360 4.000 271.960 ;
    END
  END mem_raddr_o[6]
  PIN mem_raddr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.000 4.000 304.600 ;
    END
  END mem_raddr_o[7]
  PIN mem_raddr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 336.640 4.000 337.240 ;
    END
  END mem_raddr_o[8]
  PIN mem_renb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END mem_renb_o[0]
  PIN mem_renb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END mem_renb_o[1]
  PIN mem_waddr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END mem_waddr_o[0]
  PIN mem_waddr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END mem_waddr_o[1]
  PIN mem_waddr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.920 4.000 147.520 ;
    END
  END mem_waddr_o[2]
  PIN mem_waddr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 179.560 4.000 180.160 ;
    END
  END mem_waddr_o[3]
  PIN mem_waddr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END mem_waddr_o[4]
  PIN mem_waddr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END mem_waddr_o[5]
  PIN mem_waddr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END mem_waddr_o[6]
  PIN mem_waddr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.800 4.000 311.400 ;
    END
  END mem_waddr_o[7]
  PIN mem_waddr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END mem_waddr_o[8]
  PIN mem_wenb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END mem_wenb_o[0]
  PIN mem_wenb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END mem_wenb_o[1]
  PIN oversample_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 729.680 900.000 730.280 ;
    END
  END oversample_o[0]
  PIN oversample_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 736.480 900.000 737.080 ;
    END
  END oversample_o[1]
  PIN oversample_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 743.960 900.000 744.560 ;
    END
  END oversample_o[2]
  PIN oversample_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 751.440 900.000 752.040 ;
    END
  END oversample_o[3]
  PIN oversample_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 758.920 900.000 759.520 ;
    END
  END oversample_o[4]
  PIN oversample_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 766.400 900.000 767.000 ;
    END
  END oversample_o[5]
  PIN oversample_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 773.200 900.000 773.800 ;
    END
  END oversample_o[6]
  PIN oversample_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 780.680 900.000 781.280 ;
    END
  END oversample_o[7]
  PIN oversample_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 788.160 900.000 788.760 ;
    END
  END oversample_o[8]
  PIN oversample_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 795.640 900.000 796.240 ;
    END
  END oversample_o[9]
  PIN sinc3_en_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 796.000 872.530 800.000 ;
    END
  END sinc3_en_o[0]
  PIN sinc3_en_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 796.000 883.570 800.000 ;
    END
  END sinc3_en_o[1]
  PIN sinc3_en_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 796.000 894.610 800.000 ;
    END
  END sinc3_en_o[2]
  PIN vco_enb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 796.000 839.410 800.000 ;
    END
  END vco_enb_o[0]
  PIN vco_enb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 796.000 850.450 800.000 ;
    END
  END vco_enb_o[1]
  PIN vco_enb_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 796.000 861.490 800.000 ;
    END
  END vco_enb_o[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 0.000 334.330 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.890 0.000 359.170 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 408.110 0.000 408.390 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.790 0.000 458.070 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.630 0.000 482.910 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 0.000 507.750 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 532.310 0.000 532.590 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.690 0.000 556.970 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.110 0.000 86.390 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 0.000 631.490 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.050 0.000 656.330 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.730 0.000 706.010 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.110 0.000 730.390 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.950 0.000 755.230 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 779.790 0.000 780.070 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.630 0.000 804.910 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.470 0.000 829.750 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.310 0.000 854.590 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 0.000 152.630 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.690 0.000 234.970 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.530 0.000 259.810 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.710 0.000 366.990 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 0.000 391.830 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.390 0.000 416.670 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.230 0.000 441.510 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.590 0.000 540.870 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 0.000 565.250 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.390 0.000 94.670 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.490 0.000 639.770 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 0.000 664.610 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.170 0.000 689.450 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.010 0.000 714.290 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.390 0.000 738.670 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.230 0.000 763.510 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.910 0.000 813.190 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.510 0.000 127.790 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 837.750 0.000 838.030 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.590 0.000 862.870 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 0.000 218.410 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.490 0.000 317.770 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 0.000 69.830 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 350.610 0.000 350.890 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.990 0.000 375.270 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.830 0.000 400.110 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.670 0.000 424.950 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 0.000 449.790 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.350 0.000 474.630 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 0.000 499.470 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.030 0.000 524.310 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.410 0.000 548.690 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 0.000 573.530 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.930 0.000 623.210 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.770 0.000 648.050 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.610 0.000 672.890 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 0.000 697.730 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.290 0.000 722.570 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.670 0.000 746.950 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.510 0.000 771.790 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 0.000 796.630 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.190 0.000 821.470 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.910 0.000 169.190 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.410 0.000 226.690 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 0.000 111.230 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 0.000 144.350 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 0.000 177.470 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 0.000 44.990 4.000 ;
    END
  END wbs_we_i
  PIN wmask_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END wmask_o[0]
  PIN wmask_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.880 4.000 9.480 ;
    END
  END wmask_o[1]
  PIN wmask_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 15.680 4.000 16.280 ;
    END
  END wmask_o[2]
  PIN wmask_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 21.800 4.000 22.400 ;
    END
  END wmask_o[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 789.040 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 788.800 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 788.800 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 788.800 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 788.800 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 788.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 788.800 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 788.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 788.800 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 788.800 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 788.800 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 788.800 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 788.800 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 7.225 895.015 788.885 ;
      LAYER met1 ;
        RECT 3.750 7.180 896.010 789.040 ;
      LAYER met2 ;
        RECT 3.780 795.720 4.870 796.125 ;
        RECT 5.710 795.720 15.450 796.125 ;
        RECT 16.290 795.720 26.490 796.125 ;
        RECT 27.330 795.720 37.530 796.125 ;
        RECT 38.370 795.720 48.570 796.125 ;
        RECT 49.410 795.720 59.610 796.125 ;
        RECT 60.450 795.720 70.650 796.125 ;
        RECT 71.490 795.720 81.690 796.125 ;
        RECT 82.530 795.720 92.270 796.125 ;
        RECT 93.110 795.720 103.310 796.125 ;
        RECT 104.150 795.720 114.350 796.125 ;
        RECT 115.190 795.720 125.390 796.125 ;
        RECT 126.230 795.720 136.430 796.125 ;
        RECT 137.270 795.720 147.470 796.125 ;
        RECT 148.310 795.720 158.510 796.125 ;
        RECT 159.350 795.720 169.090 796.125 ;
        RECT 169.930 795.720 180.130 796.125 ;
        RECT 180.970 795.720 191.170 796.125 ;
        RECT 192.010 795.720 202.210 796.125 ;
        RECT 203.050 795.720 213.250 796.125 ;
        RECT 214.090 795.720 224.290 796.125 ;
        RECT 225.130 795.720 235.330 796.125 ;
        RECT 236.170 795.720 246.370 796.125 ;
        RECT 247.210 795.720 256.950 796.125 ;
        RECT 257.790 795.720 267.990 796.125 ;
        RECT 268.830 795.720 279.030 796.125 ;
        RECT 279.870 795.720 290.070 796.125 ;
        RECT 290.910 795.720 301.110 796.125 ;
        RECT 301.950 795.720 312.150 796.125 ;
        RECT 312.990 795.720 323.190 796.125 ;
        RECT 324.030 795.720 333.770 796.125 ;
        RECT 334.610 795.720 344.810 796.125 ;
        RECT 345.650 795.720 355.850 796.125 ;
        RECT 356.690 795.720 366.890 796.125 ;
        RECT 367.730 795.720 377.930 796.125 ;
        RECT 378.770 795.720 388.970 796.125 ;
        RECT 389.810 795.720 400.010 796.125 ;
        RECT 400.850 795.720 411.050 796.125 ;
        RECT 411.890 795.720 421.630 796.125 ;
        RECT 422.470 795.720 432.670 796.125 ;
        RECT 433.510 795.720 443.710 796.125 ;
        RECT 444.550 795.720 454.750 796.125 ;
        RECT 455.590 795.720 465.790 796.125 ;
        RECT 466.630 795.720 476.830 796.125 ;
        RECT 477.670 795.720 487.870 796.125 ;
        RECT 488.710 795.720 498.450 796.125 ;
        RECT 499.290 795.720 509.490 796.125 ;
        RECT 510.330 795.720 520.530 796.125 ;
        RECT 521.370 795.720 531.570 796.125 ;
        RECT 532.410 795.720 542.610 796.125 ;
        RECT 543.450 795.720 553.650 796.125 ;
        RECT 554.490 795.720 564.690 796.125 ;
        RECT 565.530 795.720 575.730 796.125 ;
        RECT 576.570 795.720 586.310 796.125 ;
        RECT 587.150 795.720 597.350 796.125 ;
        RECT 598.190 795.720 608.390 796.125 ;
        RECT 609.230 795.720 619.430 796.125 ;
        RECT 620.270 795.720 630.470 796.125 ;
        RECT 631.310 795.720 641.510 796.125 ;
        RECT 642.350 795.720 652.550 796.125 ;
        RECT 653.390 795.720 663.130 796.125 ;
        RECT 663.970 795.720 674.170 796.125 ;
        RECT 675.010 795.720 685.210 796.125 ;
        RECT 686.050 795.720 696.250 796.125 ;
        RECT 697.090 795.720 707.290 796.125 ;
        RECT 708.130 795.720 718.330 796.125 ;
        RECT 719.170 795.720 729.370 796.125 ;
        RECT 730.210 795.720 740.410 796.125 ;
        RECT 741.250 795.720 750.990 796.125 ;
        RECT 751.830 795.720 762.030 796.125 ;
        RECT 762.870 795.720 773.070 796.125 ;
        RECT 773.910 795.720 784.110 796.125 ;
        RECT 784.950 795.720 795.150 796.125 ;
        RECT 795.990 795.720 806.190 796.125 ;
        RECT 807.030 795.720 817.230 796.125 ;
        RECT 818.070 795.720 827.810 796.125 ;
        RECT 828.650 795.720 838.850 796.125 ;
        RECT 839.690 795.720 849.890 796.125 ;
        RECT 850.730 795.720 860.930 796.125 ;
        RECT 861.770 795.720 871.970 796.125 ;
        RECT 872.810 795.720 883.010 796.125 ;
        RECT 883.850 795.720 894.050 796.125 ;
        RECT 894.890 795.720 895.980 796.125 ;
        RECT 3.780 4.280 895.980 795.720 ;
        RECT 4.330 2.875 11.310 4.280 ;
        RECT 12.150 2.875 19.590 4.280 ;
        RECT 20.430 2.875 27.870 4.280 ;
        RECT 28.710 2.875 36.150 4.280 ;
        RECT 36.990 2.875 44.430 4.280 ;
        RECT 45.270 2.875 52.710 4.280 ;
        RECT 53.550 2.875 60.990 4.280 ;
        RECT 61.830 2.875 69.270 4.280 ;
        RECT 70.110 2.875 77.550 4.280 ;
        RECT 78.390 2.875 85.830 4.280 ;
        RECT 86.670 2.875 94.110 4.280 ;
        RECT 94.950 2.875 102.390 4.280 ;
        RECT 103.230 2.875 110.670 4.280 ;
        RECT 111.510 2.875 118.950 4.280 ;
        RECT 119.790 2.875 127.230 4.280 ;
        RECT 128.070 2.875 135.510 4.280 ;
        RECT 136.350 2.875 143.790 4.280 ;
        RECT 144.630 2.875 152.070 4.280 ;
        RECT 152.910 2.875 160.350 4.280 ;
        RECT 161.190 2.875 168.630 4.280 ;
        RECT 169.470 2.875 176.910 4.280 ;
        RECT 177.750 2.875 184.730 4.280 ;
        RECT 185.570 2.875 193.010 4.280 ;
        RECT 193.850 2.875 201.290 4.280 ;
        RECT 202.130 2.875 209.570 4.280 ;
        RECT 210.410 2.875 217.850 4.280 ;
        RECT 218.690 2.875 226.130 4.280 ;
        RECT 226.970 2.875 234.410 4.280 ;
        RECT 235.250 2.875 242.690 4.280 ;
        RECT 243.530 2.875 250.970 4.280 ;
        RECT 251.810 2.875 259.250 4.280 ;
        RECT 260.090 2.875 267.530 4.280 ;
        RECT 268.370 2.875 275.810 4.280 ;
        RECT 276.650 2.875 284.090 4.280 ;
        RECT 284.930 2.875 292.370 4.280 ;
        RECT 293.210 2.875 300.650 4.280 ;
        RECT 301.490 2.875 308.930 4.280 ;
        RECT 309.770 2.875 317.210 4.280 ;
        RECT 318.050 2.875 325.490 4.280 ;
        RECT 326.330 2.875 333.770 4.280 ;
        RECT 334.610 2.875 342.050 4.280 ;
        RECT 342.890 2.875 350.330 4.280 ;
        RECT 351.170 2.875 358.610 4.280 ;
        RECT 359.450 2.875 366.430 4.280 ;
        RECT 367.270 2.875 374.710 4.280 ;
        RECT 375.550 2.875 382.990 4.280 ;
        RECT 383.830 2.875 391.270 4.280 ;
        RECT 392.110 2.875 399.550 4.280 ;
        RECT 400.390 2.875 407.830 4.280 ;
        RECT 408.670 2.875 416.110 4.280 ;
        RECT 416.950 2.875 424.390 4.280 ;
        RECT 425.230 2.875 432.670 4.280 ;
        RECT 433.510 2.875 440.950 4.280 ;
        RECT 441.790 2.875 449.230 4.280 ;
        RECT 450.070 2.875 457.510 4.280 ;
        RECT 458.350 2.875 465.790 4.280 ;
        RECT 466.630 2.875 474.070 4.280 ;
        RECT 474.910 2.875 482.350 4.280 ;
        RECT 483.190 2.875 490.630 4.280 ;
        RECT 491.470 2.875 498.910 4.280 ;
        RECT 499.750 2.875 507.190 4.280 ;
        RECT 508.030 2.875 515.470 4.280 ;
        RECT 516.310 2.875 523.750 4.280 ;
        RECT 524.590 2.875 532.030 4.280 ;
        RECT 532.870 2.875 540.310 4.280 ;
        RECT 541.150 2.875 548.130 4.280 ;
        RECT 548.970 2.875 556.410 4.280 ;
        RECT 557.250 2.875 564.690 4.280 ;
        RECT 565.530 2.875 572.970 4.280 ;
        RECT 573.810 2.875 581.250 4.280 ;
        RECT 582.090 2.875 589.530 4.280 ;
        RECT 590.370 2.875 597.810 4.280 ;
        RECT 598.650 2.875 606.090 4.280 ;
        RECT 606.930 2.875 614.370 4.280 ;
        RECT 615.210 2.875 622.650 4.280 ;
        RECT 623.490 2.875 630.930 4.280 ;
        RECT 631.770 2.875 639.210 4.280 ;
        RECT 640.050 2.875 647.490 4.280 ;
        RECT 648.330 2.875 655.770 4.280 ;
        RECT 656.610 2.875 664.050 4.280 ;
        RECT 664.890 2.875 672.330 4.280 ;
        RECT 673.170 2.875 680.610 4.280 ;
        RECT 681.450 2.875 688.890 4.280 ;
        RECT 689.730 2.875 697.170 4.280 ;
        RECT 698.010 2.875 705.450 4.280 ;
        RECT 706.290 2.875 713.730 4.280 ;
        RECT 714.570 2.875 722.010 4.280 ;
        RECT 722.850 2.875 729.830 4.280 ;
        RECT 730.670 2.875 738.110 4.280 ;
        RECT 738.950 2.875 746.390 4.280 ;
        RECT 747.230 2.875 754.670 4.280 ;
        RECT 755.510 2.875 762.950 4.280 ;
        RECT 763.790 2.875 771.230 4.280 ;
        RECT 772.070 2.875 779.510 4.280 ;
        RECT 780.350 2.875 787.790 4.280 ;
        RECT 788.630 2.875 796.070 4.280 ;
        RECT 796.910 2.875 804.350 4.280 ;
        RECT 805.190 2.875 812.630 4.280 ;
        RECT 813.470 2.875 820.910 4.280 ;
        RECT 821.750 2.875 829.190 4.280 ;
        RECT 830.030 2.875 837.470 4.280 ;
        RECT 838.310 2.875 845.750 4.280 ;
        RECT 846.590 2.875 854.030 4.280 ;
        RECT 854.870 2.875 862.310 4.280 ;
        RECT 863.150 2.875 870.590 4.280 ;
        RECT 871.430 2.875 878.870 4.280 ;
        RECT 879.710 2.875 887.150 4.280 ;
        RECT 887.990 2.875 895.430 4.280 ;
      LAYER met3 ;
        RECT 4.400 795.240 895.600 796.105 ;
        RECT 4.000 789.840 896.000 795.240 ;
        RECT 4.400 789.160 896.000 789.840 ;
        RECT 4.400 788.440 895.600 789.160 ;
        RECT 4.000 787.760 895.600 788.440 ;
        RECT 4.000 783.720 896.000 787.760 ;
        RECT 4.400 782.320 896.000 783.720 ;
        RECT 4.000 781.680 896.000 782.320 ;
        RECT 4.000 780.280 895.600 781.680 ;
        RECT 4.000 776.920 896.000 780.280 ;
        RECT 4.400 775.520 896.000 776.920 ;
        RECT 4.000 774.200 896.000 775.520 ;
        RECT 4.000 772.800 895.600 774.200 ;
        RECT 4.000 770.120 896.000 772.800 ;
        RECT 4.400 768.720 896.000 770.120 ;
        RECT 4.000 767.400 896.000 768.720 ;
        RECT 4.000 766.000 895.600 767.400 ;
        RECT 4.000 764.000 896.000 766.000 ;
        RECT 4.400 762.600 896.000 764.000 ;
        RECT 4.000 759.920 896.000 762.600 ;
        RECT 4.000 758.520 895.600 759.920 ;
        RECT 4.000 757.200 896.000 758.520 ;
        RECT 4.400 755.800 896.000 757.200 ;
        RECT 4.000 752.440 896.000 755.800 ;
        RECT 4.000 751.040 895.600 752.440 ;
        RECT 4.000 750.400 896.000 751.040 ;
        RECT 4.400 749.000 896.000 750.400 ;
        RECT 4.000 744.960 896.000 749.000 ;
        RECT 4.000 744.280 895.600 744.960 ;
        RECT 4.400 743.560 895.600 744.280 ;
        RECT 4.400 742.880 896.000 743.560 ;
        RECT 4.000 737.480 896.000 742.880 ;
        RECT 4.400 736.080 895.600 737.480 ;
        RECT 4.000 730.680 896.000 736.080 ;
        RECT 4.400 729.280 895.600 730.680 ;
        RECT 4.000 724.560 896.000 729.280 ;
        RECT 4.400 723.200 896.000 724.560 ;
        RECT 4.400 723.160 895.600 723.200 ;
        RECT 4.000 721.800 895.600 723.160 ;
        RECT 4.000 717.760 896.000 721.800 ;
        RECT 4.400 716.360 896.000 717.760 ;
        RECT 4.000 715.720 896.000 716.360 ;
        RECT 4.000 714.320 895.600 715.720 ;
        RECT 4.000 711.640 896.000 714.320 ;
        RECT 4.400 710.240 896.000 711.640 ;
        RECT 4.000 708.240 896.000 710.240 ;
        RECT 4.000 706.840 895.600 708.240 ;
        RECT 4.000 704.840 896.000 706.840 ;
        RECT 4.400 703.440 896.000 704.840 ;
        RECT 4.000 700.760 896.000 703.440 ;
        RECT 4.000 699.360 895.600 700.760 ;
        RECT 4.000 698.040 896.000 699.360 ;
        RECT 4.400 696.640 896.000 698.040 ;
        RECT 4.000 693.960 896.000 696.640 ;
        RECT 4.000 692.560 895.600 693.960 ;
        RECT 4.000 691.920 896.000 692.560 ;
        RECT 4.400 690.520 896.000 691.920 ;
        RECT 4.000 686.480 896.000 690.520 ;
        RECT 4.000 685.120 895.600 686.480 ;
        RECT 4.400 685.080 895.600 685.120 ;
        RECT 4.400 683.720 896.000 685.080 ;
        RECT 4.000 679.000 896.000 683.720 ;
        RECT 4.000 678.320 895.600 679.000 ;
        RECT 4.400 677.600 895.600 678.320 ;
        RECT 4.400 676.920 896.000 677.600 ;
        RECT 4.000 672.200 896.000 676.920 ;
        RECT 4.400 671.520 896.000 672.200 ;
        RECT 4.400 670.800 895.600 671.520 ;
        RECT 4.000 670.120 895.600 670.800 ;
        RECT 4.000 665.400 896.000 670.120 ;
        RECT 4.400 664.720 896.000 665.400 ;
        RECT 4.400 664.000 895.600 664.720 ;
        RECT 4.000 663.320 895.600 664.000 ;
        RECT 4.000 658.600 896.000 663.320 ;
        RECT 4.400 657.240 896.000 658.600 ;
        RECT 4.400 657.200 895.600 657.240 ;
        RECT 4.000 655.840 895.600 657.200 ;
        RECT 4.000 652.480 896.000 655.840 ;
        RECT 4.400 651.080 896.000 652.480 ;
        RECT 4.000 649.760 896.000 651.080 ;
        RECT 4.000 648.360 895.600 649.760 ;
        RECT 4.000 645.680 896.000 648.360 ;
        RECT 4.400 644.280 896.000 645.680 ;
        RECT 4.000 642.280 896.000 644.280 ;
        RECT 4.000 640.880 895.600 642.280 ;
        RECT 4.000 639.560 896.000 640.880 ;
        RECT 4.400 638.160 896.000 639.560 ;
        RECT 4.000 634.800 896.000 638.160 ;
        RECT 4.000 633.400 895.600 634.800 ;
        RECT 4.000 632.760 896.000 633.400 ;
        RECT 4.400 631.360 896.000 632.760 ;
        RECT 4.000 628.000 896.000 631.360 ;
        RECT 4.000 626.600 895.600 628.000 ;
        RECT 4.000 625.960 896.000 626.600 ;
        RECT 4.400 624.560 896.000 625.960 ;
        RECT 4.000 620.520 896.000 624.560 ;
        RECT 4.000 619.840 895.600 620.520 ;
        RECT 4.400 619.120 895.600 619.840 ;
        RECT 4.400 618.440 896.000 619.120 ;
        RECT 4.000 613.040 896.000 618.440 ;
        RECT 4.400 611.640 895.600 613.040 ;
        RECT 4.000 606.240 896.000 611.640 ;
        RECT 4.400 605.560 896.000 606.240 ;
        RECT 4.400 604.840 895.600 605.560 ;
        RECT 4.000 604.160 895.600 604.840 ;
        RECT 4.000 600.120 896.000 604.160 ;
        RECT 4.400 598.720 896.000 600.120 ;
        RECT 4.000 598.080 896.000 598.720 ;
        RECT 4.000 596.680 895.600 598.080 ;
        RECT 4.000 593.320 896.000 596.680 ;
        RECT 4.400 591.920 896.000 593.320 ;
        RECT 4.000 591.280 896.000 591.920 ;
        RECT 4.000 589.880 895.600 591.280 ;
        RECT 4.000 586.520 896.000 589.880 ;
        RECT 4.400 585.120 896.000 586.520 ;
        RECT 4.000 583.800 896.000 585.120 ;
        RECT 4.000 582.400 895.600 583.800 ;
        RECT 4.000 580.400 896.000 582.400 ;
        RECT 4.400 579.000 896.000 580.400 ;
        RECT 4.000 576.320 896.000 579.000 ;
        RECT 4.000 574.920 895.600 576.320 ;
        RECT 4.000 573.600 896.000 574.920 ;
        RECT 4.400 572.200 896.000 573.600 ;
        RECT 4.000 568.840 896.000 572.200 ;
        RECT 4.000 567.440 895.600 568.840 ;
        RECT 4.000 566.800 896.000 567.440 ;
        RECT 4.400 565.400 896.000 566.800 ;
        RECT 4.000 561.360 896.000 565.400 ;
        RECT 4.000 560.680 895.600 561.360 ;
        RECT 4.400 559.960 895.600 560.680 ;
        RECT 4.400 559.280 896.000 559.960 ;
        RECT 4.000 554.560 896.000 559.280 ;
        RECT 4.000 553.880 895.600 554.560 ;
        RECT 4.400 553.160 895.600 553.880 ;
        RECT 4.400 552.480 896.000 553.160 ;
        RECT 4.000 547.760 896.000 552.480 ;
        RECT 4.400 547.080 896.000 547.760 ;
        RECT 4.400 546.360 895.600 547.080 ;
        RECT 4.000 545.680 895.600 546.360 ;
        RECT 4.000 540.960 896.000 545.680 ;
        RECT 4.400 539.600 896.000 540.960 ;
        RECT 4.400 539.560 895.600 539.600 ;
        RECT 4.000 538.200 895.600 539.560 ;
        RECT 4.000 534.160 896.000 538.200 ;
        RECT 4.400 532.760 896.000 534.160 ;
        RECT 4.000 532.120 896.000 532.760 ;
        RECT 4.000 530.720 895.600 532.120 ;
        RECT 4.000 528.040 896.000 530.720 ;
        RECT 4.400 526.640 896.000 528.040 ;
        RECT 4.000 525.320 896.000 526.640 ;
        RECT 4.000 523.920 895.600 525.320 ;
        RECT 4.000 521.240 896.000 523.920 ;
        RECT 4.400 519.840 896.000 521.240 ;
        RECT 4.000 517.840 896.000 519.840 ;
        RECT 4.000 516.440 895.600 517.840 ;
        RECT 4.000 514.440 896.000 516.440 ;
        RECT 4.400 513.040 896.000 514.440 ;
        RECT 4.000 510.360 896.000 513.040 ;
        RECT 4.000 508.960 895.600 510.360 ;
        RECT 4.000 508.320 896.000 508.960 ;
        RECT 4.400 506.920 896.000 508.320 ;
        RECT 4.000 502.880 896.000 506.920 ;
        RECT 4.000 501.520 895.600 502.880 ;
        RECT 4.400 501.480 895.600 501.520 ;
        RECT 4.400 500.120 896.000 501.480 ;
        RECT 4.000 495.400 896.000 500.120 ;
        RECT 4.000 494.720 895.600 495.400 ;
        RECT 4.400 494.000 895.600 494.720 ;
        RECT 4.400 493.320 896.000 494.000 ;
        RECT 4.000 488.600 896.000 493.320 ;
        RECT 4.400 487.200 895.600 488.600 ;
        RECT 4.000 481.800 896.000 487.200 ;
        RECT 4.400 481.120 896.000 481.800 ;
        RECT 4.400 480.400 895.600 481.120 ;
        RECT 4.000 479.720 895.600 480.400 ;
        RECT 4.000 475.680 896.000 479.720 ;
        RECT 4.400 474.280 896.000 475.680 ;
        RECT 4.000 473.640 896.000 474.280 ;
        RECT 4.000 472.240 895.600 473.640 ;
        RECT 4.000 468.880 896.000 472.240 ;
        RECT 4.400 467.480 896.000 468.880 ;
        RECT 4.000 466.160 896.000 467.480 ;
        RECT 4.000 464.760 895.600 466.160 ;
        RECT 4.000 462.080 896.000 464.760 ;
        RECT 4.400 460.680 896.000 462.080 ;
        RECT 4.000 458.680 896.000 460.680 ;
        RECT 4.000 457.280 895.600 458.680 ;
        RECT 4.000 455.960 896.000 457.280 ;
        RECT 4.400 454.560 896.000 455.960 ;
        RECT 4.000 451.880 896.000 454.560 ;
        RECT 4.000 450.480 895.600 451.880 ;
        RECT 4.000 449.160 896.000 450.480 ;
        RECT 4.400 447.760 896.000 449.160 ;
        RECT 4.000 444.400 896.000 447.760 ;
        RECT 4.000 443.000 895.600 444.400 ;
        RECT 4.000 442.360 896.000 443.000 ;
        RECT 4.400 440.960 896.000 442.360 ;
        RECT 4.000 436.920 896.000 440.960 ;
        RECT 4.000 436.240 895.600 436.920 ;
        RECT 4.400 435.520 895.600 436.240 ;
        RECT 4.400 434.840 896.000 435.520 ;
        RECT 4.000 429.440 896.000 434.840 ;
        RECT 4.400 428.040 895.600 429.440 ;
        RECT 4.000 422.640 896.000 428.040 ;
        RECT 4.400 421.960 896.000 422.640 ;
        RECT 4.400 421.240 895.600 421.960 ;
        RECT 4.000 420.560 895.600 421.240 ;
        RECT 4.000 416.520 896.000 420.560 ;
        RECT 4.400 415.160 896.000 416.520 ;
        RECT 4.400 415.120 895.600 415.160 ;
        RECT 4.000 413.760 895.600 415.120 ;
        RECT 4.000 409.720 896.000 413.760 ;
        RECT 4.400 408.320 896.000 409.720 ;
        RECT 4.000 407.680 896.000 408.320 ;
        RECT 4.000 406.280 895.600 407.680 ;
        RECT 4.000 403.600 896.000 406.280 ;
        RECT 4.400 402.200 896.000 403.600 ;
        RECT 4.000 400.200 896.000 402.200 ;
        RECT 4.000 398.800 895.600 400.200 ;
        RECT 4.000 396.800 896.000 398.800 ;
        RECT 4.400 395.400 896.000 396.800 ;
        RECT 4.000 392.720 896.000 395.400 ;
        RECT 4.000 391.320 895.600 392.720 ;
        RECT 4.000 390.000 896.000 391.320 ;
        RECT 4.400 388.600 896.000 390.000 ;
        RECT 4.000 385.920 896.000 388.600 ;
        RECT 4.000 384.520 895.600 385.920 ;
        RECT 4.000 383.880 896.000 384.520 ;
        RECT 4.400 382.480 896.000 383.880 ;
        RECT 4.000 378.440 896.000 382.480 ;
        RECT 4.000 377.080 895.600 378.440 ;
        RECT 4.400 377.040 895.600 377.080 ;
        RECT 4.400 375.680 896.000 377.040 ;
        RECT 4.000 370.960 896.000 375.680 ;
        RECT 4.000 370.280 895.600 370.960 ;
        RECT 4.400 369.560 895.600 370.280 ;
        RECT 4.400 368.880 896.000 369.560 ;
        RECT 4.000 364.160 896.000 368.880 ;
        RECT 4.400 363.480 896.000 364.160 ;
        RECT 4.400 362.760 895.600 363.480 ;
        RECT 4.000 362.080 895.600 362.760 ;
        RECT 4.000 357.360 896.000 362.080 ;
        RECT 4.400 356.000 896.000 357.360 ;
        RECT 4.400 355.960 895.600 356.000 ;
        RECT 4.000 354.600 895.600 355.960 ;
        RECT 4.000 350.560 896.000 354.600 ;
        RECT 4.400 349.200 896.000 350.560 ;
        RECT 4.400 349.160 895.600 349.200 ;
        RECT 4.000 347.800 895.600 349.160 ;
        RECT 4.000 344.440 896.000 347.800 ;
        RECT 4.400 343.040 896.000 344.440 ;
        RECT 4.000 341.720 896.000 343.040 ;
        RECT 4.000 340.320 895.600 341.720 ;
        RECT 4.000 337.640 896.000 340.320 ;
        RECT 4.400 336.240 896.000 337.640 ;
        RECT 4.000 334.240 896.000 336.240 ;
        RECT 4.000 332.840 895.600 334.240 ;
        RECT 4.000 330.840 896.000 332.840 ;
        RECT 4.400 329.440 896.000 330.840 ;
        RECT 4.000 326.760 896.000 329.440 ;
        RECT 4.000 325.360 895.600 326.760 ;
        RECT 4.000 324.720 896.000 325.360 ;
        RECT 4.400 323.320 896.000 324.720 ;
        RECT 4.000 319.280 896.000 323.320 ;
        RECT 4.000 317.920 895.600 319.280 ;
        RECT 4.400 317.880 895.600 317.920 ;
        RECT 4.400 316.520 896.000 317.880 ;
        RECT 4.000 312.480 896.000 316.520 ;
        RECT 4.000 311.800 895.600 312.480 ;
        RECT 4.400 311.080 895.600 311.800 ;
        RECT 4.400 310.400 896.000 311.080 ;
        RECT 4.000 305.000 896.000 310.400 ;
        RECT 4.400 303.600 895.600 305.000 ;
        RECT 4.000 298.200 896.000 303.600 ;
        RECT 4.400 297.520 896.000 298.200 ;
        RECT 4.400 296.800 895.600 297.520 ;
        RECT 4.000 296.120 895.600 296.800 ;
        RECT 4.000 292.080 896.000 296.120 ;
        RECT 4.400 290.680 896.000 292.080 ;
        RECT 4.000 290.040 896.000 290.680 ;
        RECT 4.000 288.640 895.600 290.040 ;
        RECT 4.000 285.280 896.000 288.640 ;
        RECT 4.400 283.880 896.000 285.280 ;
        RECT 4.000 282.560 896.000 283.880 ;
        RECT 4.000 281.160 895.600 282.560 ;
        RECT 4.000 278.480 896.000 281.160 ;
        RECT 4.400 277.080 896.000 278.480 ;
        RECT 4.000 275.760 896.000 277.080 ;
        RECT 4.000 274.360 895.600 275.760 ;
        RECT 4.000 272.360 896.000 274.360 ;
        RECT 4.400 270.960 896.000 272.360 ;
        RECT 4.000 268.280 896.000 270.960 ;
        RECT 4.000 266.880 895.600 268.280 ;
        RECT 4.000 265.560 896.000 266.880 ;
        RECT 4.400 264.160 896.000 265.560 ;
        RECT 4.000 260.800 896.000 264.160 ;
        RECT 4.000 259.400 895.600 260.800 ;
        RECT 4.000 258.760 896.000 259.400 ;
        RECT 4.400 257.360 896.000 258.760 ;
        RECT 4.000 253.320 896.000 257.360 ;
        RECT 4.000 252.640 895.600 253.320 ;
        RECT 4.400 251.920 895.600 252.640 ;
        RECT 4.400 251.240 896.000 251.920 ;
        RECT 4.000 246.520 896.000 251.240 ;
        RECT 4.000 245.840 895.600 246.520 ;
        RECT 4.400 245.120 895.600 245.840 ;
        RECT 4.400 244.440 896.000 245.120 ;
        RECT 4.000 239.720 896.000 244.440 ;
        RECT 4.400 239.040 896.000 239.720 ;
        RECT 4.400 238.320 895.600 239.040 ;
        RECT 4.000 237.640 895.600 238.320 ;
        RECT 4.000 232.920 896.000 237.640 ;
        RECT 4.400 231.560 896.000 232.920 ;
        RECT 4.400 231.520 895.600 231.560 ;
        RECT 4.000 230.160 895.600 231.520 ;
        RECT 4.000 226.120 896.000 230.160 ;
        RECT 4.400 224.720 896.000 226.120 ;
        RECT 4.000 224.080 896.000 224.720 ;
        RECT 4.000 222.680 895.600 224.080 ;
        RECT 4.000 220.000 896.000 222.680 ;
        RECT 4.400 218.600 896.000 220.000 ;
        RECT 4.000 216.600 896.000 218.600 ;
        RECT 4.000 215.200 895.600 216.600 ;
        RECT 4.000 213.200 896.000 215.200 ;
        RECT 4.400 211.800 896.000 213.200 ;
        RECT 4.000 209.800 896.000 211.800 ;
        RECT 4.000 208.400 895.600 209.800 ;
        RECT 4.000 206.400 896.000 208.400 ;
        RECT 4.400 205.000 896.000 206.400 ;
        RECT 4.000 202.320 896.000 205.000 ;
        RECT 4.000 200.920 895.600 202.320 ;
        RECT 4.000 200.280 896.000 200.920 ;
        RECT 4.400 198.880 896.000 200.280 ;
        RECT 4.000 194.840 896.000 198.880 ;
        RECT 4.000 193.480 895.600 194.840 ;
        RECT 4.400 193.440 895.600 193.480 ;
        RECT 4.400 192.080 896.000 193.440 ;
        RECT 4.000 187.360 896.000 192.080 ;
        RECT 4.000 186.680 895.600 187.360 ;
        RECT 4.400 185.960 895.600 186.680 ;
        RECT 4.400 185.280 896.000 185.960 ;
        RECT 4.000 180.560 896.000 185.280 ;
        RECT 4.400 179.880 896.000 180.560 ;
        RECT 4.400 179.160 895.600 179.880 ;
        RECT 4.000 178.480 895.600 179.160 ;
        RECT 4.000 173.760 896.000 178.480 ;
        RECT 4.400 173.080 896.000 173.760 ;
        RECT 4.400 172.360 895.600 173.080 ;
        RECT 4.000 171.680 895.600 172.360 ;
        RECT 4.000 166.960 896.000 171.680 ;
        RECT 4.400 165.600 896.000 166.960 ;
        RECT 4.400 165.560 895.600 165.600 ;
        RECT 4.000 164.200 895.600 165.560 ;
        RECT 4.000 160.840 896.000 164.200 ;
        RECT 4.400 159.440 896.000 160.840 ;
        RECT 4.000 158.120 896.000 159.440 ;
        RECT 4.000 156.720 895.600 158.120 ;
        RECT 4.000 154.040 896.000 156.720 ;
        RECT 4.400 152.640 896.000 154.040 ;
        RECT 4.000 150.640 896.000 152.640 ;
        RECT 4.000 149.240 895.600 150.640 ;
        RECT 4.000 147.920 896.000 149.240 ;
        RECT 4.400 146.520 896.000 147.920 ;
        RECT 4.000 143.160 896.000 146.520 ;
        RECT 4.000 141.760 895.600 143.160 ;
        RECT 4.000 141.120 896.000 141.760 ;
        RECT 4.400 139.720 896.000 141.120 ;
        RECT 4.000 136.360 896.000 139.720 ;
        RECT 4.000 134.960 895.600 136.360 ;
        RECT 4.000 134.320 896.000 134.960 ;
        RECT 4.400 132.920 896.000 134.320 ;
        RECT 4.000 128.880 896.000 132.920 ;
        RECT 4.000 128.200 895.600 128.880 ;
        RECT 4.400 127.480 895.600 128.200 ;
        RECT 4.400 126.800 896.000 127.480 ;
        RECT 4.000 121.400 896.000 126.800 ;
        RECT 4.400 120.000 895.600 121.400 ;
        RECT 4.000 114.600 896.000 120.000 ;
        RECT 4.400 113.920 896.000 114.600 ;
        RECT 4.400 113.200 895.600 113.920 ;
        RECT 4.000 112.520 895.600 113.200 ;
        RECT 4.000 108.480 896.000 112.520 ;
        RECT 4.400 107.120 896.000 108.480 ;
        RECT 4.400 107.080 895.600 107.120 ;
        RECT 4.000 105.720 895.600 107.080 ;
        RECT 4.000 101.680 896.000 105.720 ;
        RECT 4.400 100.280 896.000 101.680 ;
        RECT 4.000 99.640 896.000 100.280 ;
        RECT 4.000 98.240 895.600 99.640 ;
        RECT 4.000 94.880 896.000 98.240 ;
        RECT 4.400 93.480 896.000 94.880 ;
        RECT 4.000 92.160 896.000 93.480 ;
        RECT 4.000 90.760 895.600 92.160 ;
        RECT 4.000 88.760 896.000 90.760 ;
        RECT 4.400 87.360 896.000 88.760 ;
        RECT 4.000 84.680 896.000 87.360 ;
        RECT 4.000 83.280 895.600 84.680 ;
        RECT 4.000 81.960 896.000 83.280 ;
        RECT 4.400 80.560 896.000 81.960 ;
        RECT 4.000 77.200 896.000 80.560 ;
        RECT 4.000 75.840 895.600 77.200 ;
        RECT 4.400 75.800 895.600 75.840 ;
        RECT 4.400 74.440 896.000 75.800 ;
        RECT 4.000 70.400 896.000 74.440 ;
        RECT 4.000 69.040 895.600 70.400 ;
        RECT 4.400 69.000 895.600 69.040 ;
        RECT 4.400 67.640 896.000 69.000 ;
        RECT 4.000 62.920 896.000 67.640 ;
        RECT 4.000 62.240 895.600 62.920 ;
        RECT 4.400 61.520 895.600 62.240 ;
        RECT 4.400 60.840 896.000 61.520 ;
        RECT 4.000 56.120 896.000 60.840 ;
        RECT 4.400 55.440 896.000 56.120 ;
        RECT 4.400 54.720 895.600 55.440 ;
        RECT 4.000 54.040 895.600 54.720 ;
        RECT 4.000 49.320 896.000 54.040 ;
        RECT 4.400 47.960 896.000 49.320 ;
        RECT 4.400 47.920 895.600 47.960 ;
        RECT 4.000 46.560 895.600 47.920 ;
        RECT 4.000 42.520 896.000 46.560 ;
        RECT 4.400 41.120 896.000 42.520 ;
        RECT 4.000 40.480 896.000 41.120 ;
        RECT 4.000 39.080 895.600 40.480 ;
        RECT 4.000 36.400 896.000 39.080 ;
        RECT 4.400 35.000 896.000 36.400 ;
        RECT 4.000 33.680 896.000 35.000 ;
        RECT 4.000 32.280 895.600 33.680 ;
        RECT 4.000 29.600 896.000 32.280 ;
        RECT 4.400 28.200 896.000 29.600 ;
        RECT 4.000 26.200 896.000 28.200 ;
        RECT 4.000 24.800 895.600 26.200 ;
        RECT 4.000 22.800 896.000 24.800 ;
        RECT 4.400 21.400 896.000 22.800 ;
        RECT 4.000 18.720 896.000 21.400 ;
        RECT 4.000 17.320 895.600 18.720 ;
        RECT 4.000 16.680 896.000 17.320 ;
        RECT 4.400 15.280 896.000 16.680 ;
        RECT 4.000 11.240 896.000 15.280 ;
        RECT 4.000 9.880 895.600 11.240 ;
        RECT 4.400 9.840 895.600 9.880 ;
        RECT 4.400 8.480 896.000 9.840 ;
        RECT 4.000 4.440 896.000 8.480 ;
        RECT 4.000 3.760 895.600 4.440 ;
        RECT 4.400 3.040 895.600 3.760 ;
        RECT 4.400 2.895 896.000 3.040 ;
      LAYER met4 ;
        RECT 887.175 30.775 889.345 759.385 ;
  END
END vco_adc_wrapper
END LIBRARY

