VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ring_osc
  CLASS BLOCK ;
  FOREIGN ring_osc ;
  ORIGIN -0.500 0.290 ;
  SIZE 183.000 BY 38.660 ;
  OBS
      LAYER pwell ;
        RECT 18.390 32.310 28.420 38.370 ;
      LAYER nwell ;
        RECT 3.630 28.505 6.310 30.340 ;
        RECT 7.800 28.505 9.560 30.340 ;
      LAYER pwell ;
        RECT 4.310 27.985 6.115 28.215 ;
        RECT 3.825 27.305 6.115 27.985 ;
        RECT 3.970 27.115 4.140 27.305 ;
        RECT 8.135 27.115 8.305 27.285 ;
      LAYER nwell ;
        RECT 18.390 24.245 24.240 30.120 ;
        RECT 29.220 29.780 35.070 35.635 ;
      LAYER pwell ;
        RECT 36.365 32.270 42.215 38.370 ;
      LAYER nwell ;
        RECT 42.840 30.310 46.600 35.585 ;
      LAYER pwell ;
        RECT 47.890 32.310 57.920 38.370 ;
        RECT 25.040 21.460 35.070 27.860 ;
      LAYER nwell ;
        RECT 36.365 24.250 40.125 29.560 ;
      LAYER pwell ;
        RECT 40.745 26.625 46.595 27.565 ;
        RECT 40.745 26.575 46.600 26.625 ;
        RECT 40.750 21.465 46.600 26.575 ;
      LAYER nwell ;
        RECT 47.890 24.245 53.740 30.120 ;
        RECT 58.720 29.780 64.570 35.635 ;
      LAYER pwell ;
        RECT 65.865 32.270 71.715 38.370 ;
      LAYER nwell ;
        RECT 72.340 30.310 76.100 35.585 ;
      LAYER pwell ;
        RECT 77.390 32.310 87.420 38.370 ;
        RECT 54.540 21.460 64.570 27.860 ;
      LAYER nwell ;
        RECT 65.865 24.250 69.625 29.560 ;
      LAYER pwell ;
        RECT 70.245 26.625 76.095 27.565 ;
        RECT 70.245 26.575 76.100 26.625 ;
        RECT 70.250 21.465 76.100 26.575 ;
      LAYER nwell ;
        RECT 77.390 24.245 83.240 30.120 ;
        RECT 88.220 29.780 94.070 35.635 ;
      LAYER pwell ;
        RECT 95.365 32.270 101.215 38.370 ;
      LAYER nwell ;
        RECT 101.840 30.310 105.600 35.585 ;
      LAYER pwell ;
        RECT 106.890 32.310 116.920 38.370 ;
        RECT 84.040 21.460 94.070 27.860 ;
      LAYER nwell ;
        RECT 95.365 24.250 99.125 29.560 ;
      LAYER pwell ;
        RECT 99.745 26.625 105.595 27.565 ;
        RECT 99.745 26.575 105.600 26.625 ;
        RECT 99.750 21.465 105.600 26.575 ;
      LAYER nwell ;
        RECT 106.890 24.245 112.740 30.120 ;
        RECT 117.720 29.780 123.570 35.635 ;
      LAYER pwell ;
        RECT 124.865 32.270 130.715 38.370 ;
      LAYER nwell ;
        RECT 131.340 30.310 135.100 35.585 ;
      LAYER pwell ;
        RECT 136.390 32.310 146.420 38.370 ;
        RECT 113.540 21.460 123.570 27.860 ;
      LAYER nwell ;
        RECT 124.865 24.250 128.625 29.560 ;
      LAYER pwell ;
        RECT 129.245 26.625 135.095 27.565 ;
        RECT 129.245 26.575 135.100 26.625 ;
        RECT 129.250 21.465 135.100 26.575 ;
      LAYER nwell ;
        RECT 136.390 24.245 142.240 30.120 ;
        RECT 147.220 29.780 153.070 35.635 ;
      LAYER pwell ;
        RECT 154.365 32.270 160.215 38.370 ;
      LAYER nwell ;
        RECT 160.840 30.310 164.600 35.585 ;
      LAYER pwell ;
        RECT 143.040 21.460 153.070 27.860 ;
      LAYER nwell ;
        RECT 154.365 24.250 158.125 29.560 ;
      LAYER pwell ;
        RECT 158.745 26.625 164.595 27.565 ;
        RECT 158.745 26.575 164.600 26.625 ;
        RECT 158.750 21.465 164.600 26.575 ;
        RECT 2.790 11.505 8.640 16.615 ;
        RECT 2.790 11.455 8.645 11.505 ;
        RECT 2.795 10.515 8.645 11.455 ;
      LAYER nwell ;
        RECT 9.265 8.520 13.025 13.830 ;
      LAYER pwell ;
        RECT 14.320 10.220 24.350 16.620 ;
      LAYER nwell ;
        RECT 2.790 2.495 6.550 7.770 ;
      LAYER pwell ;
        RECT 7.175 -0.290 13.025 5.810 ;
      LAYER nwell ;
        RECT 14.320 2.445 20.170 8.300 ;
        RECT 25.150 7.960 31.000 13.835 ;
      LAYER pwell ;
        RECT 32.290 11.505 38.140 16.615 ;
        RECT 32.290 11.455 38.145 11.505 ;
        RECT 32.295 10.515 38.145 11.455 ;
      LAYER nwell ;
        RECT 38.765 8.520 42.525 13.830 ;
      LAYER pwell ;
        RECT 43.820 10.220 53.850 16.620 ;
        RECT 20.970 -0.290 31.000 5.770 ;
      LAYER nwell ;
        RECT 32.290 2.495 36.050 7.770 ;
      LAYER pwell ;
        RECT 36.675 -0.290 42.525 5.810 ;
      LAYER nwell ;
        RECT 43.820 2.445 49.670 8.300 ;
        RECT 54.650 7.960 60.500 13.835 ;
      LAYER pwell ;
        RECT 61.790 11.505 67.640 16.615 ;
        RECT 61.790 11.455 67.645 11.505 ;
        RECT 61.795 10.515 67.645 11.455 ;
      LAYER nwell ;
        RECT 68.265 8.520 72.025 13.830 ;
      LAYER pwell ;
        RECT 73.320 10.220 83.350 16.620 ;
        RECT 50.470 -0.290 60.500 5.770 ;
      LAYER nwell ;
        RECT 61.790 2.495 65.550 7.770 ;
      LAYER pwell ;
        RECT 66.175 -0.290 72.025 5.810 ;
      LAYER nwell ;
        RECT 73.320 2.445 79.170 8.300 ;
        RECT 84.150 7.960 90.000 13.835 ;
      LAYER pwell ;
        RECT 91.290 11.505 97.140 16.615 ;
        RECT 91.290 11.455 97.145 11.505 ;
        RECT 91.295 10.515 97.145 11.455 ;
      LAYER nwell ;
        RECT 97.765 8.520 101.525 13.830 ;
      LAYER pwell ;
        RECT 102.820 10.220 112.850 16.620 ;
        RECT 79.970 -0.290 90.000 5.770 ;
      LAYER nwell ;
        RECT 91.290 2.495 95.050 7.770 ;
      LAYER pwell ;
        RECT 95.675 -0.290 101.525 5.810 ;
      LAYER nwell ;
        RECT 102.820 2.445 108.670 8.300 ;
        RECT 113.650 7.960 119.500 13.835 ;
      LAYER pwell ;
        RECT 120.790 11.505 126.640 16.615 ;
        RECT 120.790 11.455 126.645 11.505 ;
        RECT 120.795 10.515 126.645 11.455 ;
      LAYER nwell ;
        RECT 127.265 8.520 131.025 13.830 ;
      LAYER pwell ;
        RECT 132.320 10.220 142.350 16.620 ;
        RECT 109.470 -0.290 119.500 5.770 ;
      LAYER nwell ;
        RECT 120.790 2.495 124.550 7.770 ;
      LAYER pwell ;
        RECT 125.175 -0.290 131.025 5.810 ;
      LAYER nwell ;
        RECT 132.320 2.445 138.170 8.300 ;
        RECT 143.150 7.960 149.000 13.835 ;
      LAYER pwell ;
        RECT 150.290 11.505 156.140 16.615 ;
        RECT 150.290 11.455 156.145 11.505 ;
        RECT 150.295 10.515 156.145 11.455 ;
      LAYER nwell ;
        RECT 156.765 8.520 160.525 13.830 ;
      LAYER pwell ;
        RECT 161.820 10.220 171.850 16.620 ;
        RECT 138.970 -0.290 149.000 5.770 ;
      LAYER nwell ;
        RECT 150.290 2.495 154.050 7.770 ;
      LAYER pwell ;
        RECT 154.675 -0.290 160.525 5.810 ;
      LAYER nwell ;
        RECT 161.820 2.445 167.670 8.300 ;
        RECT 172.650 7.960 178.500 13.835 ;
      LAYER pwell ;
        RECT 168.470 -0.290 178.500 5.770 ;
      LAYER li1 ;
        RECT 18.570 37.840 20.915 38.320 ;
        RECT 21.980 37.840 24.840 38.320 ;
        RECT 25.895 37.840 28.240 38.320 ;
        RECT 36.545 37.840 38.890 38.320 ;
        RECT 39.690 37.840 42.035 38.320 ;
        RECT 48.070 37.840 50.415 38.320 ;
        RECT 51.480 37.840 54.340 38.320 ;
        RECT 55.395 37.840 57.740 38.320 ;
        RECT 66.045 37.840 68.390 38.320 ;
        RECT 69.190 37.840 71.535 38.320 ;
        RECT 77.570 37.840 79.915 38.320 ;
        RECT 80.980 37.840 83.840 38.320 ;
        RECT 84.895 37.840 87.240 38.320 ;
        RECT 95.545 37.840 97.890 38.320 ;
        RECT 98.690 37.840 101.035 38.320 ;
        RECT 107.070 37.840 109.415 38.320 ;
        RECT 110.480 37.840 113.340 38.320 ;
        RECT 114.395 37.840 116.740 38.320 ;
        RECT 125.045 37.840 127.390 38.320 ;
        RECT 128.190 37.840 130.535 38.320 ;
        RECT 136.570 37.840 138.915 38.320 ;
        RECT 139.980 37.840 142.840 38.320 ;
        RECT 143.895 37.840 146.240 38.320 ;
        RECT 154.545 37.840 156.890 38.320 ;
        RECT 157.690 37.840 160.035 38.320 ;
        RECT 19.080 33.245 19.370 37.840 ;
        RECT 19.140 33.000 19.310 33.245 ;
        RECT 19.290 30.790 20.420 31.790 ;
        RECT 21.170 31.480 21.460 37.540 ;
        RECT 23.260 33.245 23.550 37.840 ;
        RECT 23.320 33.000 23.490 33.245 ;
        RECT 25.350 31.580 25.640 37.540 ;
        RECT 27.440 33.245 27.730 37.840 ;
        RECT 29.400 35.455 31.745 35.600 ;
        RECT 32.545 35.455 34.890 35.600 ;
        RECT 29.400 35.285 34.890 35.455 ;
        RECT 29.400 35.120 31.745 35.285 ;
        RECT 32.545 35.120 34.890 35.285 ;
        RECT 27.500 33.235 27.695 33.245 ;
        RECT 27.500 33.000 27.670 33.235 ;
        RECT 25.350 31.480 26.170 31.580 ;
        RECT 21.170 30.980 26.170 31.480 ;
        RECT 4.340 30.005 5.310 30.160 ;
        RECT 8.340 30.005 9.310 30.160 ;
        RECT 3.820 29.835 6.120 30.005 ;
        RECT 7.990 29.835 9.370 30.005 ;
        RECT 3.905 29.265 4.165 29.665 ;
        RECT 4.335 29.435 5.270 29.835 ;
        RECT 5.440 29.325 6.035 29.665 ;
        RECT 3.905 29.095 5.270 29.265 ;
        RECT 3.905 28.195 4.365 28.925 ;
        RECT 4.535 28.025 5.270 29.095 ;
        RECT 3.905 27.855 5.270 28.025 ;
        RECT 5.440 28.005 5.615 29.325 ;
        RECT 6.330 29.155 7.780 29.375 ;
        RECT 5.795 29.075 7.780 29.155 ;
        RECT 8.265 29.110 8.595 29.835 ;
        RECT 5.795 28.855 6.630 29.075 ;
        RECT 7.480 28.940 7.780 29.075 ;
        RECT 5.795 28.175 6.035 28.855 ;
        RECT 5.440 27.875 6.035 28.005 ;
        RECT 6.860 27.875 7.160 28.710 ;
        RECT 7.480 28.640 8.595 28.940 ;
        RECT 3.905 27.455 4.165 27.855 ;
        RECT 4.335 27.285 5.270 27.685 ;
        RECT 5.440 27.575 7.160 27.875 ;
        RECT 5.440 27.455 6.035 27.575 ;
        RECT 8.075 27.455 8.595 28.640 ;
        RECT 8.765 28.115 9.285 29.665 ;
        RECT 8.765 27.285 9.105 27.945 ;
        RECT 3.820 27.115 6.120 27.285 ;
        RECT 7.990 27.115 9.370 27.285 ;
        RECT 18.570 24.720 18.740 29.575 ;
        RECT 19.080 24.720 19.370 29.570 ;
        RECT 21.170 25.030 21.460 30.980 ;
        RECT 29.400 30.460 29.570 35.120 ;
        RECT 29.910 30.290 30.200 35.120 ;
        RECT 32.000 29.850 32.290 34.850 ;
        RECT 34.090 30.290 34.380 35.120 ;
        RECT 34.720 30.520 34.890 35.120 ;
        RECT 37.055 33.490 37.345 37.840 ;
        RECT 37.290 31.580 38.490 31.890 ;
        RECT 36.790 30.960 38.490 31.580 ;
        RECT 37.290 30.760 38.490 30.960 ;
        RECT 39.140 29.850 39.435 37.530 ;
        RECT 41.235 33.490 41.525 37.840 ;
        RECT 44.325 35.570 46.420 35.600 ;
        RECT 44.170 35.405 46.420 35.570 ;
        RECT 43.020 35.235 46.420 35.405 ;
        RECT 43.020 32.260 43.190 35.235 ;
        RECT 44.170 35.150 46.420 35.235 ;
        RECT 44.325 35.120 46.420 35.150 ;
        RECT 43.525 31.675 43.820 34.750 ;
        RECT 43.295 30.895 44.035 31.675 ;
        RECT 23.260 24.720 23.550 29.570 ;
        RECT 23.890 24.720 24.060 29.575 ;
        RECT 29.360 29.350 41.955 29.850 ;
        RECT 29.360 27.910 29.860 29.350 ;
        RECT 30.890 28.320 34.890 28.920 ;
        RECT 32.890 28.200 34.890 28.320 ;
        RECT 27.820 27.620 32.290 27.910 ;
        RECT 32.890 27.620 34.090 28.200 ;
        RECT 25.790 26.595 25.960 26.830 ;
        RECT 25.765 26.585 25.960 26.595 ;
        RECT 18.570 24.595 20.915 24.720 ;
        RECT 21.715 24.690 24.060 24.720 ;
        RECT 21.715 24.595 24.240 24.690 ;
        RECT 18.570 24.425 24.240 24.595 ;
        RECT 18.570 24.240 20.915 24.425 ;
        RECT 21.715 24.270 24.240 24.425 ;
        RECT 21.715 24.240 24.060 24.270 ;
        RECT 25.730 22.000 26.020 26.585 ;
        RECT 27.820 22.290 28.110 27.620 ;
        RECT 29.970 26.585 30.140 26.810 ;
        RECT 29.910 22.000 30.200 26.585 ;
        RECT 32.000 22.290 32.290 27.620 ;
        RECT 34.150 26.585 34.320 26.810 ;
        RECT 34.090 22.000 34.380 26.585 ;
        RECT 36.545 24.720 36.715 28.645 ;
        RECT 37.055 24.720 37.345 28.790 ;
        RECT 39.145 25.085 39.440 29.350 ;
        RECT 36.545 24.690 38.640 24.720 ;
        RECT 36.545 24.600 38.795 24.690 ;
        RECT 39.775 24.600 39.945 28.635 ;
        RECT 41.455 28.200 41.955 29.350 ;
        RECT 36.545 24.430 39.945 24.600 ;
        RECT 36.545 24.270 38.795 24.430 ;
        RECT 36.545 24.240 38.640 24.270 ;
        RECT 41.440 22.000 41.730 26.345 ;
        RECT 43.525 22.305 43.820 30.895 ;
        RECT 45.620 30.710 45.910 35.120 ;
        RECT 46.250 30.705 46.420 35.120 ;
        RECT 48.580 33.245 48.870 37.840 ;
        RECT 48.640 33.000 48.810 33.245 ;
        RECT 48.790 30.790 49.920 31.790 ;
        RECT 50.670 31.480 50.960 37.540 ;
        RECT 52.760 33.245 53.050 37.840 ;
        RECT 52.820 33.000 52.990 33.245 ;
        RECT 54.850 31.580 55.140 37.540 ;
        RECT 56.940 33.245 57.230 37.840 ;
        RECT 58.900 35.455 61.245 35.600 ;
        RECT 62.045 35.455 64.390 35.600 ;
        RECT 58.900 35.285 64.390 35.455 ;
        RECT 58.900 35.120 61.245 35.285 ;
        RECT 62.045 35.120 64.390 35.285 ;
        RECT 57.000 33.235 57.195 33.245 ;
        RECT 57.000 33.000 57.170 33.235 ;
        RECT 54.850 31.480 55.670 31.580 ;
        RECT 50.670 30.980 55.670 31.480 ;
        RECT 44.440 28.860 45.620 29.060 ;
        RECT 44.440 28.260 46.120 28.860 ;
        RECT 44.440 27.980 45.620 28.260 ;
        RECT 45.620 22.000 45.910 26.345 ;
        RECT 48.070 24.720 48.240 29.575 ;
        RECT 48.580 24.720 48.870 29.570 ;
        RECT 50.670 25.030 50.960 30.980 ;
        RECT 58.900 30.460 59.070 35.120 ;
        RECT 59.410 30.290 59.700 35.120 ;
        RECT 61.500 29.850 61.790 34.850 ;
        RECT 63.590 30.290 63.880 35.120 ;
        RECT 64.220 30.520 64.390 35.120 ;
        RECT 66.555 33.490 66.845 37.840 ;
        RECT 66.790 31.580 67.990 31.890 ;
        RECT 66.290 30.960 67.990 31.580 ;
        RECT 66.790 30.760 67.990 30.960 ;
        RECT 68.640 29.850 68.935 37.530 ;
        RECT 70.735 33.490 71.025 37.840 ;
        RECT 73.825 35.570 75.920 35.600 ;
        RECT 73.670 35.405 75.920 35.570 ;
        RECT 72.520 35.235 75.920 35.405 ;
        RECT 72.520 32.260 72.690 35.235 ;
        RECT 73.670 35.150 75.920 35.235 ;
        RECT 73.825 35.120 75.920 35.150 ;
        RECT 73.025 31.675 73.320 34.750 ;
        RECT 72.795 30.895 73.535 31.675 ;
        RECT 52.760 24.720 53.050 29.570 ;
        RECT 53.390 24.720 53.560 29.575 ;
        RECT 58.860 29.350 71.455 29.850 ;
        RECT 58.860 27.910 59.360 29.350 ;
        RECT 60.390 28.320 64.390 28.920 ;
        RECT 62.390 28.200 64.390 28.320 ;
        RECT 57.320 27.620 61.790 27.910 ;
        RECT 62.390 27.620 63.590 28.200 ;
        RECT 55.290 26.595 55.460 26.830 ;
        RECT 55.265 26.585 55.460 26.595 ;
        RECT 48.070 24.595 50.415 24.720 ;
        RECT 51.215 24.690 53.560 24.720 ;
        RECT 51.215 24.595 53.740 24.690 ;
        RECT 48.070 24.425 53.740 24.595 ;
        RECT 48.070 24.240 50.415 24.425 ;
        RECT 51.215 24.270 53.740 24.425 ;
        RECT 51.215 24.240 53.560 24.270 ;
        RECT 55.230 22.000 55.520 26.585 ;
        RECT 57.320 22.290 57.610 27.620 ;
        RECT 59.470 26.585 59.640 26.810 ;
        RECT 59.410 22.000 59.700 26.585 ;
        RECT 61.500 22.290 61.790 27.620 ;
        RECT 63.650 26.585 63.820 26.810 ;
        RECT 63.590 22.000 63.880 26.585 ;
        RECT 66.045 24.720 66.215 28.645 ;
        RECT 66.555 24.720 66.845 28.790 ;
        RECT 68.645 25.085 68.940 29.350 ;
        RECT 66.045 24.690 68.140 24.720 ;
        RECT 66.045 24.600 68.295 24.690 ;
        RECT 69.275 24.600 69.445 28.635 ;
        RECT 70.955 28.200 71.455 29.350 ;
        RECT 66.045 24.430 69.445 24.600 ;
        RECT 66.045 24.270 68.295 24.430 ;
        RECT 66.045 24.240 68.140 24.270 ;
        RECT 70.940 22.000 71.230 26.345 ;
        RECT 73.025 22.305 73.320 30.895 ;
        RECT 75.120 30.710 75.410 35.120 ;
        RECT 75.750 30.705 75.920 35.120 ;
        RECT 78.080 33.245 78.370 37.840 ;
        RECT 78.140 33.000 78.310 33.245 ;
        RECT 78.290 30.790 79.420 31.790 ;
        RECT 80.170 31.480 80.460 37.540 ;
        RECT 82.260 33.245 82.550 37.840 ;
        RECT 82.320 33.000 82.490 33.245 ;
        RECT 84.350 31.580 84.640 37.540 ;
        RECT 86.440 33.245 86.730 37.840 ;
        RECT 88.400 35.455 90.745 35.600 ;
        RECT 91.545 35.455 93.890 35.600 ;
        RECT 88.400 35.285 93.890 35.455 ;
        RECT 88.400 35.120 90.745 35.285 ;
        RECT 91.545 35.120 93.890 35.285 ;
        RECT 86.500 33.235 86.695 33.245 ;
        RECT 86.500 33.000 86.670 33.235 ;
        RECT 84.350 31.480 85.170 31.580 ;
        RECT 80.170 30.980 85.170 31.480 ;
        RECT 73.940 28.860 75.120 29.060 ;
        RECT 73.940 28.260 75.620 28.860 ;
        RECT 73.940 27.980 75.120 28.260 ;
        RECT 75.120 22.000 75.410 26.345 ;
        RECT 77.570 24.720 77.740 29.575 ;
        RECT 78.080 24.720 78.370 29.570 ;
        RECT 80.170 25.030 80.460 30.980 ;
        RECT 88.400 30.460 88.570 35.120 ;
        RECT 88.910 30.290 89.200 35.120 ;
        RECT 91.000 29.850 91.290 34.850 ;
        RECT 93.090 30.290 93.380 35.120 ;
        RECT 93.720 30.520 93.890 35.120 ;
        RECT 96.055 33.490 96.345 37.840 ;
        RECT 96.290 31.580 97.490 31.890 ;
        RECT 95.790 30.960 97.490 31.580 ;
        RECT 96.290 30.760 97.490 30.960 ;
        RECT 98.140 29.850 98.435 37.530 ;
        RECT 100.235 33.490 100.525 37.840 ;
        RECT 103.325 35.570 105.420 35.600 ;
        RECT 103.170 35.405 105.420 35.570 ;
        RECT 102.020 35.235 105.420 35.405 ;
        RECT 102.020 32.260 102.190 35.235 ;
        RECT 103.170 35.150 105.420 35.235 ;
        RECT 103.325 35.120 105.420 35.150 ;
        RECT 102.525 31.675 102.820 34.750 ;
        RECT 102.295 30.895 103.035 31.675 ;
        RECT 82.260 24.720 82.550 29.570 ;
        RECT 82.890 24.720 83.060 29.575 ;
        RECT 88.360 29.350 100.955 29.850 ;
        RECT 88.360 27.910 88.860 29.350 ;
        RECT 89.890 28.320 93.890 28.920 ;
        RECT 91.890 28.200 93.890 28.320 ;
        RECT 86.820 27.620 91.290 27.910 ;
        RECT 91.890 27.620 93.090 28.200 ;
        RECT 84.790 26.595 84.960 26.830 ;
        RECT 84.765 26.585 84.960 26.595 ;
        RECT 77.570 24.595 79.915 24.720 ;
        RECT 80.715 24.690 83.060 24.720 ;
        RECT 80.715 24.595 83.240 24.690 ;
        RECT 77.570 24.425 83.240 24.595 ;
        RECT 77.570 24.240 79.915 24.425 ;
        RECT 80.715 24.270 83.240 24.425 ;
        RECT 80.715 24.240 83.060 24.270 ;
        RECT 84.730 22.000 85.020 26.585 ;
        RECT 86.820 22.290 87.110 27.620 ;
        RECT 88.970 26.585 89.140 26.810 ;
        RECT 88.910 22.000 89.200 26.585 ;
        RECT 91.000 22.290 91.290 27.620 ;
        RECT 93.150 26.585 93.320 26.810 ;
        RECT 93.090 22.000 93.380 26.585 ;
        RECT 95.545 24.720 95.715 28.645 ;
        RECT 96.055 24.720 96.345 28.790 ;
        RECT 98.145 25.085 98.440 29.350 ;
        RECT 95.545 24.690 97.640 24.720 ;
        RECT 95.545 24.600 97.795 24.690 ;
        RECT 98.775 24.600 98.945 28.635 ;
        RECT 100.455 28.200 100.955 29.350 ;
        RECT 95.545 24.430 98.945 24.600 ;
        RECT 95.545 24.270 97.795 24.430 ;
        RECT 95.545 24.240 97.640 24.270 ;
        RECT 100.440 22.000 100.730 26.345 ;
        RECT 102.525 22.305 102.820 30.895 ;
        RECT 104.620 30.710 104.910 35.120 ;
        RECT 105.250 30.705 105.420 35.120 ;
        RECT 107.580 33.245 107.870 37.840 ;
        RECT 107.640 33.000 107.810 33.245 ;
        RECT 107.790 30.790 108.920 31.790 ;
        RECT 109.670 31.480 109.960 37.540 ;
        RECT 111.760 33.245 112.050 37.840 ;
        RECT 111.820 33.000 111.990 33.245 ;
        RECT 113.850 31.580 114.140 37.540 ;
        RECT 115.940 33.245 116.230 37.840 ;
        RECT 117.900 35.455 120.245 35.600 ;
        RECT 121.045 35.455 123.390 35.600 ;
        RECT 117.900 35.285 123.390 35.455 ;
        RECT 117.900 35.120 120.245 35.285 ;
        RECT 121.045 35.120 123.390 35.285 ;
        RECT 116.000 33.235 116.195 33.245 ;
        RECT 116.000 33.000 116.170 33.235 ;
        RECT 113.850 31.480 114.670 31.580 ;
        RECT 109.670 30.980 114.670 31.480 ;
        RECT 103.440 28.860 104.620 29.060 ;
        RECT 103.440 28.260 105.120 28.860 ;
        RECT 103.440 27.980 104.620 28.260 ;
        RECT 104.620 22.000 104.910 26.345 ;
        RECT 107.070 24.720 107.240 29.575 ;
        RECT 107.580 24.720 107.870 29.570 ;
        RECT 109.670 25.030 109.960 30.980 ;
        RECT 117.900 30.460 118.070 35.120 ;
        RECT 118.410 30.290 118.700 35.120 ;
        RECT 120.500 29.850 120.790 34.850 ;
        RECT 122.590 30.290 122.880 35.120 ;
        RECT 123.220 30.520 123.390 35.120 ;
        RECT 125.555 33.490 125.845 37.840 ;
        RECT 125.790 31.580 126.990 31.890 ;
        RECT 125.290 30.960 126.990 31.580 ;
        RECT 125.790 30.760 126.990 30.960 ;
        RECT 127.640 29.850 127.935 37.530 ;
        RECT 129.735 33.490 130.025 37.840 ;
        RECT 132.825 35.570 134.920 35.600 ;
        RECT 132.670 35.405 134.920 35.570 ;
        RECT 131.520 35.235 134.920 35.405 ;
        RECT 131.520 32.260 131.690 35.235 ;
        RECT 132.670 35.150 134.920 35.235 ;
        RECT 132.825 35.120 134.920 35.150 ;
        RECT 132.025 31.675 132.320 34.750 ;
        RECT 131.795 30.895 132.535 31.675 ;
        RECT 111.760 24.720 112.050 29.570 ;
        RECT 112.390 24.720 112.560 29.575 ;
        RECT 117.860 29.350 130.455 29.850 ;
        RECT 117.860 27.910 118.360 29.350 ;
        RECT 119.390 28.320 123.390 28.920 ;
        RECT 121.390 28.200 123.390 28.320 ;
        RECT 116.320 27.620 120.790 27.910 ;
        RECT 121.390 27.620 122.590 28.200 ;
        RECT 114.290 26.595 114.460 26.830 ;
        RECT 114.265 26.585 114.460 26.595 ;
        RECT 107.070 24.595 109.415 24.720 ;
        RECT 110.215 24.690 112.560 24.720 ;
        RECT 110.215 24.595 112.740 24.690 ;
        RECT 107.070 24.425 112.740 24.595 ;
        RECT 107.070 24.240 109.415 24.425 ;
        RECT 110.215 24.270 112.740 24.425 ;
        RECT 110.215 24.240 112.560 24.270 ;
        RECT 114.230 22.000 114.520 26.585 ;
        RECT 116.320 22.290 116.610 27.620 ;
        RECT 118.470 26.585 118.640 26.810 ;
        RECT 118.410 22.000 118.700 26.585 ;
        RECT 120.500 22.290 120.790 27.620 ;
        RECT 122.650 26.585 122.820 26.810 ;
        RECT 122.590 22.000 122.880 26.585 ;
        RECT 125.045 24.720 125.215 28.645 ;
        RECT 125.555 24.720 125.845 28.790 ;
        RECT 127.645 25.085 127.940 29.350 ;
        RECT 125.045 24.690 127.140 24.720 ;
        RECT 125.045 24.600 127.295 24.690 ;
        RECT 128.275 24.600 128.445 28.635 ;
        RECT 129.955 28.200 130.455 29.350 ;
        RECT 125.045 24.430 128.445 24.600 ;
        RECT 125.045 24.270 127.295 24.430 ;
        RECT 125.045 24.240 127.140 24.270 ;
        RECT 129.940 22.000 130.230 26.345 ;
        RECT 132.025 22.305 132.320 30.895 ;
        RECT 134.120 30.710 134.410 35.120 ;
        RECT 134.750 30.705 134.920 35.120 ;
        RECT 137.080 33.245 137.370 37.840 ;
        RECT 137.140 33.000 137.310 33.245 ;
        RECT 137.290 30.790 138.420 31.790 ;
        RECT 139.170 31.480 139.460 37.540 ;
        RECT 141.260 33.245 141.550 37.840 ;
        RECT 141.320 33.000 141.490 33.245 ;
        RECT 143.350 31.580 143.640 37.540 ;
        RECT 145.440 33.245 145.730 37.840 ;
        RECT 147.400 35.455 149.745 35.600 ;
        RECT 150.545 35.455 152.890 35.600 ;
        RECT 147.400 35.285 152.890 35.455 ;
        RECT 147.400 35.120 149.745 35.285 ;
        RECT 150.545 35.120 152.890 35.285 ;
        RECT 145.500 33.235 145.695 33.245 ;
        RECT 145.500 33.000 145.670 33.235 ;
        RECT 143.350 31.480 144.170 31.580 ;
        RECT 139.170 30.980 144.170 31.480 ;
        RECT 132.940 28.860 134.120 29.060 ;
        RECT 132.940 28.260 134.620 28.860 ;
        RECT 132.940 27.980 134.120 28.260 ;
        RECT 134.120 22.000 134.410 26.345 ;
        RECT 136.570 24.720 136.740 29.575 ;
        RECT 137.080 24.720 137.370 29.570 ;
        RECT 139.170 25.030 139.460 30.980 ;
        RECT 147.400 30.460 147.570 35.120 ;
        RECT 147.910 30.290 148.200 35.120 ;
        RECT 150.000 29.850 150.290 34.850 ;
        RECT 152.090 30.290 152.380 35.120 ;
        RECT 152.720 30.520 152.890 35.120 ;
        RECT 155.055 33.490 155.345 37.840 ;
        RECT 155.290 31.580 156.490 31.890 ;
        RECT 154.790 30.960 156.490 31.580 ;
        RECT 155.290 30.760 156.490 30.960 ;
        RECT 157.140 29.850 157.435 37.530 ;
        RECT 159.235 33.490 159.525 37.840 ;
        RECT 162.325 35.570 164.420 35.600 ;
        RECT 162.170 35.405 164.420 35.570 ;
        RECT 161.020 35.235 164.420 35.405 ;
        RECT 161.020 32.260 161.190 35.235 ;
        RECT 162.170 35.150 164.420 35.235 ;
        RECT 162.325 35.120 164.420 35.150 ;
        RECT 161.525 31.675 161.820 34.750 ;
        RECT 161.295 30.895 162.035 31.675 ;
        RECT 141.260 24.720 141.550 29.570 ;
        RECT 141.890 24.720 142.060 29.575 ;
        RECT 147.360 29.350 159.955 29.850 ;
        RECT 147.360 27.910 147.860 29.350 ;
        RECT 148.890 28.320 152.890 28.920 ;
        RECT 150.890 28.200 152.890 28.320 ;
        RECT 145.820 27.620 150.290 27.910 ;
        RECT 150.890 27.620 152.090 28.200 ;
        RECT 143.790 26.595 143.960 26.830 ;
        RECT 143.765 26.585 143.960 26.595 ;
        RECT 136.570 24.595 138.915 24.720 ;
        RECT 139.715 24.690 142.060 24.720 ;
        RECT 139.715 24.595 142.240 24.690 ;
        RECT 136.570 24.425 142.240 24.595 ;
        RECT 136.570 24.240 138.915 24.425 ;
        RECT 139.715 24.270 142.240 24.425 ;
        RECT 139.715 24.240 142.060 24.270 ;
        RECT 143.730 22.000 144.020 26.585 ;
        RECT 145.820 22.290 146.110 27.620 ;
        RECT 147.970 26.585 148.140 26.810 ;
        RECT 147.910 22.000 148.200 26.585 ;
        RECT 150.000 22.290 150.290 27.620 ;
        RECT 152.150 26.585 152.320 26.810 ;
        RECT 152.090 22.000 152.380 26.585 ;
        RECT 154.545 24.720 154.715 28.645 ;
        RECT 155.055 24.720 155.345 28.790 ;
        RECT 157.145 25.085 157.440 29.350 ;
        RECT 154.545 24.690 156.640 24.720 ;
        RECT 154.545 24.600 156.795 24.690 ;
        RECT 157.775 24.600 157.945 28.635 ;
        RECT 159.455 28.200 159.955 29.350 ;
        RECT 154.545 24.430 157.945 24.600 ;
        RECT 154.545 24.270 156.795 24.430 ;
        RECT 154.545 24.240 156.640 24.270 ;
        RECT 159.440 22.000 159.730 26.345 ;
        RECT 161.525 22.305 161.820 30.895 ;
        RECT 163.620 30.710 163.910 35.120 ;
        RECT 164.250 30.705 164.420 35.120 ;
        RECT 162.440 28.860 163.620 29.060 ;
        RECT 162.440 28.260 164.120 28.860 ;
        RECT 162.440 27.980 163.620 28.260 ;
        RECT 163.620 22.000 163.910 26.345 ;
        RECT 25.220 21.520 27.570 22.000 ;
        RECT 28.620 21.520 31.480 22.000 ;
        RECT 32.545 21.520 34.890 22.000 ;
        RECT 40.930 21.970 43.270 22.000 ;
        RECT 44.080 21.970 46.420 22.000 ;
        RECT 40.930 21.550 43.275 21.970 ;
        RECT 44.075 21.550 46.420 21.970 ;
        RECT 40.930 21.520 43.270 21.550 ;
        RECT 44.080 21.520 46.420 21.550 ;
        RECT 54.720 21.520 57.070 22.000 ;
        RECT 58.120 21.520 60.980 22.000 ;
        RECT 62.045 21.520 64.390 22.000 ;
        RECT 70.430 21.970 72.770 22.000 ;
        RECT 73.580 21.970 75.920 22.000 ;
        RECT 70.430 21.550 72.775 21.970 ;
        RECT 73.575 21.550 75.920 21.970 ;
        RECT 70.430 21.520 72.770 21.550 ;
        RECT 73.580 21.520 75.920 21.550 ;
        RECT 84.220 21.520 86.570 22.000 ;
        RECT 87.620 21.520 90.480 22.000 ;
        RECT 91.545 21.520 93.890 22.000 ;
        RECT 99.930 21.970 102.270 22.000 ;
        RECT 103.080 21.970 105.420 22.000 ;
        RECT 99.930 21.550 102.275 21.970 ;
        RECT 103.075 21.550 105.420 21.970 ;
        RECT 99.930 21.520 102.270 21.550 ;
        RECT 103.080 21.520 105.420 21.550 ;
        RECT 113.720 21.520 116.070 22.000 ;
        RECT 117.120 21.520 119.980 22.000 ;
        RECT 121.045 21.520 123.390 22.000 ;
        RECT 129.430 21.970 131.770 22.000 ;
        RECT 132.580 21.970 134.920 22.000 ;
        RECT 129.430 21.550 131.775 21.970 ;
        RECT 132.575 21.550 134.920 21.970 ;
        RECT 129.430 21.520 131.770 21.550 ;
        RECT 132.580 21.520 134.920 21.550 ;
        RECT 143.220 21.520 145.570 22.000 ;
        RECT 146.620 21.520 149.480 22.000 ;
        RECT 150.545 21.520 152.890 22.000 ;
        RECT 158.930 21.970 161.270 22.000 ;
        RECT 162.080 21.970 164.420 22.000 ;
        RECT 158.930 21.550 161.275 21.970 ;
        RECT 162.075 21.550 164.420 21.970 ;
        RECT 158.930 21.520 161.270 21.550 ;
        RECT 162.080 21.520 164.420 21.550 ;
        RECT 2.970 16.530 5.310 16.560 ;
        RECT 6.120 16.530 8.460 16.560 ;
        RECT 2.970 16.110 5.315 16.530 ;
        RECT 6.115 16.110 8.460 16.530 ;
        RECT 2.970 16.080 5.310 16.110 ;
        RECT 6.120 16.080 8.460 16.110 ;
        RECT 14.500 16.080 16.845 16.560 ;
        RECT 17.910 16.080 20.770 16.560 ;
        RECT 21.820 16.080 24.170 16.560 ;
        RECT 32.470 16.530 34.810 16.560 ;
        RECT 35.620 16.530 37.960 16.560 ;
        RECT 32.470 16.110 34.815 16.530 ;
        RECT 35.615 16.110 37.960 16.530 ;
        RECT 32.470 16.080 34.810 16.110 ;
        RECT 35.620 16.080 37.960 16.110 ;
        RECT 44.000 16.080 46.345 16.560 ;
        RECT 47.410 16.080 50.270 16.560 ;
        RECT 51.320 16.080 53.670 16.560 ;
        RECT 61.970 16.530 64.310 16.560 ;
        RECT 65.120 16.530 67.460 16.560 ;
        RECT 61.970 16.110 64.315 16.530 ;
        RECT 65.115 16.110 67.460 16.530 ;
        RECT 61.970 16.080 64.310 16.110 ;
        RECT 65.120 16.080 67.460 16.110 ;
        RECT 73.500 16.080 75.845 16.560 ;
        RECT 76.910 16.080 79.770 16.560 ;
        RECT 80.820 16.080 83.170 16.560 ;
        RECT 91.470 16.530 93.810 16.560 ;
        RECT 94.620 16.530 96.960 16.560 ;
        RECT 91.470 16.110 93.815 16.530 ;
        RECT 94.615 16.110 96.960 16.530 ;
        RECT 91.470 16.080 93.810 16.110 ;
        RECT 94.620 16.080 96.960 16.110 ;
        RECT 103.000 16.080 105.345 16.560 ;
        RECT 106.410 16.080 109.270 16.560 ;
        RECT 110.320 16.080 112.670 16.560 ;
        RECT 120.970 16.530 123.310 16.560 ;
        RECT 124.120 16.530 126.460 16.560 ;
        RECT 120.970 16.110 123.315 16.530 ;
        RECT 124.115 16.110 126.460 16.530 ;
        RECT 120.970 16.080 123.310 16.110 ;
        RECT 124.120 16.080 126.460 16.110 ;
        RECT 132.500 16.080 134.845 16.560 ;
        RECT 135.910 16.080 138.770 16.560 ;
        RECT 139.820 16.080 142.170 16.560 ;
        RECT 150.470 16.530 152.810 16.560 ;
        RECT 153.620 16.530 155.960 16.560 ;
        RECT 150.470 16.110 152.815 16.530 ;
        RECT 153.615 16.110 155.960 16.530 ;
        RECT 150.470 16.080 152.810 16.110 ;
        RECT 153.620 16.080 155.960 16.110 ;
        RECT 162.000 16.080 164.345 16.560 ;
        RECT 165.410 16.080 168.270 16.560 ;
        RECT 169.320 16.080 171.670 16.560 ;
        RECT 3.480 11.735 3.770 16.080 ;
        RECT 3.770 9.820 4.950 10.100 ;
        RECT 3.270 9.220 4.950 9.820 ;
        RECT 3.770 9.020 4.950 9.220 ;
        RECT 2.970 2.960 3.140 7.375 ;
        RECT 3.480 2.960 3.770 7.370 ;
        RECT 5.570 7.185 5.865 15.775 ;
        RECT 7.660 11.735 7.950 16.080 ;
        RECT 10.750 13.810 12.845 13.840 ;
        RECT 10.595 13.650 12.845 13.810 ;
        RECT 9.445 13.480 12.845 13.650 ;
        RECT 7.435 8.730 7.935 9.880 ;
        RECT 9.445 9.445 9.615 13.480 ;
        RECT 10.595 13.390 12.845 13.480 ;
        RECT 10.750 13.360 12.845 13.390 ;
        RECT 9.950 8.730 10.245 12.995 ;
        RECT 12.045 9.290 12.335 13.360 ;
        RECT 12.675 9.435 12.845 13.360 ;
        RECT 15.010 11.495 15.300 16.080 ;
        RECT 15.070 11.270 15.240 11.495 ;
        RECT 17.100 10.460 17.390 15.790 ;
        RECT 19.190 11.495 19.480 16.080 ;
        RECT 19.250 11.270 19.420 11.495 ;
        RECT 21.280 10.460 21.570 15.790 ;
        RECT 23.370 11.495 23.660 16.080 ;
        RECT 25.330 13.810 27.675 13.840 ;
        RECT 25.150 13.655 27.675 13.810 ;
        RECT 28.475 13.655 30.820 13.840 ;
        RECT 25.150 13.485 30.820 13.655 ;
        RECT 25.150 13.390 27.675 13.485 ;
        RECT 25.330 13.360 27.675 13.390 ;
        RECT 28.475 13.360 30.820 13.485 ;
        RECT 23.430 11.485 23.625 11.495 ;
        RECT 23.430 11.250 23.600 11.485 ;
        RECT 15.300 9.880 16.500 10.460 ;
        RECT 17.100 10.170 21.570 10.460 ;
        RECT 14.500 9.760 16.500 9.880 ;
        RECT 14.500 9.160 18.500 9.760 ;
        RECT 19.530 8.730 20.030 10.170 ;
        RECT 7.435 8.230 20.030 8.730 ;
        RECT 25.330 8.505 25.500 13.360 ;
        RECT 25.840 8.510 26.130 13.360 ;
        RECT 5.355 6.405 6.095 7.185 ;
        RECT 5.570 3.330 5.865 6.405 ;
        RECT 2.970 2.930 5.065 2.960 ;
        RECT 2.970 2.845 5.220 2.930 ;
        RECT 6.200 2.845 6.370 5.820 ;
        RECT 2.970 2.675 6.370 2.845 ;
        RECT 2.970 2.510 5.220 2.675 ;
        RECT 2.970 2.480 5.065 2.510 ;
        RECT 7.865 0.240 8.155 4.590 ;
        RECT 9.955 0.550 10.250 8.230 ;
        RECT 10.900 7.120 12.100 7.320 ;
        RECT 10.900 6.500 12.600 7.120 ;
        RECT 10.900 6.190 12.100 6.500 ;
        RECT 12.045 0.240 12.335 4.590 ;
        RECT 14.500 2.960 14.670 7.560 ;
        RECT 15.010 2.960 15.300 7.790 ;
        RECT 17.100 3.230 17.390 8.230 ;
        RECT 19.190 2.960 19.480 7.790 ;
        RECT 19.820 2.960 19.990 7.620 ;
        RECT 27.930 7.100 28.220 13.050 ;
        RECT 30.020 8.510 30.310 13.360 ;
        RECT 30.650 8.505 30.820 13.360 ;
        RECT 32.980 11.735 33.270 16.080 ;
        RECT 33.270 9.820 34.450 10.100 ;
        RECT 32.770 9.220 34.450 9.820 ;
        RECT 33.270 9.020 34.450 9.220 ;
        RECT 23.220 6.600 28.220 7.100 ;
        RECT 23.220 6.500 24.040 6.600 ;
        RECT 21.720 4.845 21.890 5.080 ;
        RECT 21.695 4.835 21.890 4.845 ;
        RECT 14.500 2.795 16.845 2.960 ;
        RECT 17.645 2.795 19.990 2.960 ;
        RECT 14.500 2.625 19.990 2.795 ;
        RECT 14.500 2.480 16.845 2.625 ;
        RECT 17.645 2.480 19.990 2.625 ;
        RECT 21.660 0.240 21.950 4.835 ;
        RECT 23.750 0.540 24.040 6.500 ;
        RECT 25.900 4.835 26.070 5.080 ;
        RECT 25.840 0.240 26.130 4.835 ;
        RECT 27.930 0.540 28.220 6.600 ;
        RECT 28.970 6.290 30.100 7.290 ;
        RECT 30.080 4.835 30.250 5.080 ;
        RECT 30.020 0.240 30.310 4.835 ;
        RECT 32.470 2.960 32.640 7.375 ;
        RECT 32.980 2.960 33.270 7.370 ;
        RECT 35.070 7.185 35.365 15.775 ;
        RECT 37.160 11.735 37.450 16.080 ;
        RECT 40.250 13.810 42.345 13.840 ;
        RECT 40.095 13.650 42.345 13.810 ;
        RECT 38.945 13.480 42.345 13.650 ;
        RECT 36.935 8.730 37.435 9.880 ;
        RECT 38.945 9.445 39.115 13.480 ;
        RECT 40.095 13.390 42.345 13.480 ;
        RECT 40.250 13.360 42.345 13.390 ;
        RECT 39.450 8.730 39.745 12.995 ;
        RECT 41.545 9.290 41.835 13.360 ;
        RECT 42.175 9.435 42.345 13.360 ;
        RECT 44.510 11.495 44.800 16.080 ;
        RECT 44.570 11.270 44.740 11.495 ;
        RECT 46.600 10.460 46.890 15.790 ;
        RECT 48.690 11.495 48.980 16.080 ;
        RECT 48.750 11.270 48.920 11.495 ;
        RECT 50.780 10.460 51.070 15.790 ;
        RECT 52.870 11.495 53.160 16.080 ;
        RECT 54.830 13.810 57.175 13.840 ;
        RECT 54.650 13.655 57.175 13.810 ;
        RECT 57.975 13.655 60.320 13.840 ;
        RECT 54.650 13.485 60.320 13.655 ;
        RECT 54.650 13.390 57.175 13.485 ;
        RECT 54.830 13.360 57.175 13.390 ;
        RECT 57.975 13.360 60.320 13.485 ;
        RECT 52.930 11.485 53.125 11.495 ;
        RECT 52.930 11.250 53.100 11.485 ;
        RECT 44.800 9.880 46.000 10.460 ;
        RECT 46.600 10.170 51.070 10.460 ;
        RECT 44.000 9.760 46.000 9.880 ;
        RECT 44.000 9.160 48.000 9.760 ;
        RECT 49.030 8.730 49.530 10.170 ;
        RECT 36.935 8.230 49.530 8.730 ;
        RECT 54.830 8.505 55.000 13.360 ;
        RECT 55.340 8.510 55.630 13.360 ;
        RECT 34.855 6.405 35.595 7.185 ;
        RECT 35.070 3.330 35.365 6.405 ;
        RECT 32.470 2.930 34.565 2.960 ;
        RECT 32.470 2.845 34.720 2.930 ;
        RECT 35.700 2.845 35.870 5.820 ;
        RECT 32.470 2.675 35.870 2.845 ;
        RECT 32.470 2.510 34.720 2.675 ;
        RECT 32.470 2.480 34.565 2.510 ;
        RECT 37.365 0.240 37.655 4.590 ;
        RECT 39.455 0.550 39.750 8.230 ;
        RECT 40.400 7.120 41.600 7.320 ;
        RECT 40.400 6.500 42.100 7.120 ;
        RECT 40.400 6.190 41.600 6.500 ;
        RECT 41.545 0.240 41.835 4.590 ;
        RECT 44.000 2.960 44.170 7.560 ;
        RECT 44.510 2.960 44.800 7.790 ;
        RECT 46.600 3.230 46.890 8.230 ;
        RECT 48.690 2.960 48.980 7.790 ;
        RECT 49.320 2.960 49.490 7.620 ;
        RECT 57.430 7.100 57.720 13.050 ;
        RECT 59.520 8.510 59.810 13.360 ;
        RECT 60.150 8.505 60.320 13.360 ;
        RECT 62.480 11.735 62.770 16.080 ;
        RECT 62.770 9.820 63.950 10.100 ;
        RECT 62.270 9.220 63.950 9.820 ;
        RECT 62.770 9.020 63.950 9.220 ;
        RECT 52.720 6.600 57.720 7.100 ;
        RECT 52.720 6.500 53.540 6.600 ;
        RECT 51.220 4.845 51.390 5.080 ;
        RECT 51.195 4.835 51.390 4.845 ;
        RECT 44.000 2.795 46.345 2.960 ;
        RECT 47.145 2.795 49.490 2.960 ;
        RECT 44.000 2.625 49.490 2.795 ;
        RECT 44.000 2.480 46.345 2.625 ;
        RECT 47.145 2.480 49.490 2.625 ;
        RECT 51.160 0.240 51.450 4.835 ;
        RECT 53.250 0.540 53.540 6.500 ;
        RECT 55.400 4.835 55.570 5.080 ;
        RECT 55.340 0.240 55.630 4.835 ;
        RECT 57.430 0.540 57.720 6.600 ;
        RECT 58.470 6.290 59.600 7.290 ;
        RECT 59.580 4.835 59.750 5.080 ;
        RECT 59.520 0.240 59.810 4.835 ;
        RECT 61.970 2.960 62.140 7.375 ;
        RECT 62.480 2.960 62.770 7.370 ;
        RECT 64.570 7.185 64.865 15.775 ;
        RECT 66.660 11.735 66.950 16.080 ;
        RECT 69.750 13.810 71.845 13.840 ;
        RECT 69.595 13.650 71.845 13.810 ;
        RECT 68.445 13.480 71.845 13.650 ;
        RECT 66.435 8.730 66.935 9.880 ;
        RECT 68.445 9.445 68.615 13.480 ;
        RECT 69.595 13.390 71.845 13.480 ;
        RECT 69.750 13.360 71.845 13.390 ;
        RECT 68.950 8.730 69.245 12.995 ;
        RECT 71.045 9.290 71.335 13.360 ;
        RECT 71.675 9.435 71.845 13.360 ;
        RECT 74.010 11.495 74.300 16.080 ;
        RECT 74.070 11.270 74.240 11.495 ;
        RECT 76.100 10.460 76.390 15.790 ;
        RECT 78.190 11.495 78.480 16.080 ;
        RECT 78.250 11.270 78.420 11.495 ;
        RECT 80.280 10.460 80.570 15.790 ;
        RECT 82.370 11.495 82.660 16.080 ;
        RECT 84.330 13.810 86.675 13.840 ;
        RECT 84.150 13.655 86.675 13.810 ;
        RECT 87.475 13.655 89.820 13.840 ;
        RECT 84.150 13.485 89.820 13.655 ;
        RECT 84.150 13.390 86.675 13.485 ;
        RECT 84.330 13.360 86.675 13.390 ;
        RECT 87.475 13.360 89.820 13.485 ;
        RECT 82.430 11.485 82.625 11.495 ;
        RECT 82.430 11.250 82.600 11.485 ;
        RECT 74.300 9.880 75.500 10.460 ;
        RECT 76.100 10.170 80.570 10.460 ;
        RECT 73.500 9.760 75.500 9.880 ;
        RECT 73.500 9.160 77.500 9.760 ;
        RECT 78.530 8.730 79.030 10.170 ;
        RECT 66.435 8.230 79.030 8.730 ;
        RECT 84.330 8.505 84.500 13.360 ;
        RECT 84.840 8.510 85.130 13.360 ;
        RECT 64.355 6.405 65.095 7.185 ;
        RECT 64.570 3.330 64.865 6.405 ;
        RECT 61.970 2.930 64.065 2.960 ;
        RECT 61.970 2.845 64.220 2.930 ;
        RECT 65.200 2.845 65.370 5.820 ;
        RECT 61.970 2.675 65.370 2.845 ;
        RECT 61.970 2.510 64.220 2.675 ;
        RECT 61.970 2.480 64.065 2.510 ;
        RECT 66.865 0.240 67.155 4.590 ;
        RECT 68.955 0.550 69.250 8.230 ;
        RECT 69.900 7.120 71.100 7.320 ;
        RECT 69.900 6.500 71.600 7.120 ;
        RECT 69.900 6.190 71.100 6.500 ;
        RECT 71.045 0.240 71.335 4.590 ;
        RECT 73.500 2.960 73.670 7.560 ;
        RECT 74.010 2.960 74.300 7.790 ;
        RECT 76.100 3.230 76.390 8.230 ;
        RECT 78.190 2.960 78.480 7.790 ;
        RECT 78.820 2.960 78.990 7.620 ;
        RECT 86.930 7.100 87.220 13.050 ;
        RECT 89.020 8.510 89.310 13.360 ;
        RECT 89.650 8.505 89.820 13.360 ;
        RECT 91.980 11.735 92.270 16.080 ;
        RECT 92.270 9.820 93.450 10.100 ;
        RECT 91.770 9.220 93.450 9.820 ;
        RECT 92.270 9.020 93.450 9.220 ;
        RECT 82.220 6.600 87.220 7.100 ;
        RECT 82.220 6.500 83.040 6.600 ;
        RECT 80.720 4.845 80.890 5.080 ;
        RECT 80.695 4.835 80.890 4.845 ;
        RECT 73.500 2.795 75.845 2.960 ;
        RECT 76.645 2.795 78.990 2.960 ;
        RECT 73.500 2.625 78.990 2.795 ;
        RECT 73.500 2.480 75.845 2.625 ;
        RECT 76.645 2.480 78.990 2.625 ;
        RECT 80.660 0.240 80.950 4.835 ;
        RECT 82.750 0.540 83.040 6.500 ;
        RECT 84.900 4.835 85.070 5.080 ;
        RECT 84.840 0.240 85.130 4.835 ;
        RECT 86.930 0.540 87.220 6.600 ;
        RECT 87.970 6.290 89.100 7.290 ;
        RECT 89.080 4.835 89.250 5.080 ;
        RECT 89.020 0.240 89.310 4.835 ;
        RECT 91.470 2.960 91.640 7.375 ;
        RECT 91.980 2.960 92.270 7.370 ;
        RECT 94.070 7.185 94.365 15.775 ;
        RECT 96.160 11.735 96.450 16.080 ;
        RECT 99.250 13.810 101.345 13.840 ;
        RECT 99.095 13.650 101.345 13.810 ;
        RECT 97.945 13.480 101.345 13.650 ;
        RECT 95.935 8.730 96.435 9.880 ;
        RECT 97.945 9.445 98.115 13.480 ;
        RECT 99.095 13.390 101.345 13.480 ;
        RECT 99.250 13.360 101.345 13.390 ;
        RECT 98.450 8.730 98.745 12.995 ;
        RECT 100.545 9.290 100.835 13.360 ;
        RECT 101.175 9.435 101.345 13.360 ;
        RECT 103.510 11.495 103.800 16.080 ;
        RECT 103.570 11.270 103.740 11.495 ;
        RECT 105.600 10.460 105.890 15.790 ;
        RECT 107.690 11.495 107.980 16.080 ;
        RECT 107.750 11.270 107.920 11.495 ;
        RECT 109.780 10.460 110.070 15.790 ;
        RECT 111.870 11.495 112.160 16.080 ;
        RECT 113.830 13.810 116.175 13.840 ;
        RECT 113.650 13.655 116.175 13.810 ;
        RECT 116.975 13.655 119.320 13.840 ;
        RECT 113.650 13.485 119.320 13.655 ;
        RECT 113.650 13.390 116.175 13.485 ;
        RECT 113.830 13.360 116.175 13.390 ;
        RECT 116.975 13.360 119.320 13.485 ;
        RECT 111.930 11.485 112.125 11.495 ;
        RECT 111.930 11.250 112.100 11.485 ;
        RECT 103.800 9.880 105.000 10.460 ;
        RECT 105.600 10.170 110.070 10.460 ;
        RECT 103.000 9.760 105.000 9.880 ;
        RECT 103.000 9.160 107.000 9.760 ;
        RECT 108.030 8.730 108.530 10.170 ;
        RECT 95.935 8.230 108.530 8.730 ;
        RECT 113.830 8.505 114.000 13.360 ;
        RECT 114.340 8.510 114.630 13.360 ;
        RECT 93.855 6.405 94.595 7.185 ;
        RECT 94.070 3.330 94.365 6.405 ;
        RECT 91.470 2.930 93.565 2.960 ;
        RECT 91.470 2.845 93.720 2.930 ;
        RECT 94.700 2.845 94.870 5.820 ;
        RECT 91.470 2.675 94.870 2.845 ;
        RECT 91.470 2.510 93.720 2.675 ;
        RECT 91.470 2.480 93.565 2.510 ;
        RECT 96.365 0.240 96.655 4.590 ;
        RECT 98.455 0.550 98.750 8.230 ;
        RECT 99.400 7.120 100.600 7.320 ;
        RECT 99.400 6.500 101.100 7.120 ;
        RECT 99.400 6.190 100.600 6.500 ;
        RECT 100.545 0.240 100.835 4.590 ;
        RECT 103.000 2.960 103.170 7.560 ;
        RECT 103.510 2.960 103.800 7.790 ;
        RECT 105.600 3.230 105.890 8.230 ;
        RECT 107.690 2.960 107.980 7.790 ;
        RECT 108.320 2.960 108.490 7.620 ;
        RECT 116.430 7.100 116.720 13.050 ;
        RECT 118.520 8.510 118.810 13.360 ;
        RECT 119.150 8.505 119.320 13.360 ;
        RECT 121.480 11.735 121.770 16.080 ;
        RECT 121.770 9.820 122.950 10.100 ;
        RECT 121.270 9.220 122.950 9.820 ;
        RECT 121.770 9.020 122.950 9.220 ;
        RECT 111.720 6.600 116.720 7.100 ;
        RECT 111.720 6.500 112.540 6.600 ;
        RECT 110.220 4.845 110.390 5.080 ;
        RECT 110.195 4.835 110.390 4.845 ;
        RECT 103.000 2.795 105.345 2.960 ;
        RECT 106.145 2.795 108.490 2.960 ;
        RECT 103.000 2.625 108.490 2.795 ;
        RECT 103.000 2.480 105.345 2.625 ;
        RECT 106.145 2.480 108.490 2.625 ;
        RECT 110.160 0.240 110.450 4.835 ;
        RECT 112.250 0.540 112.540 6.500 ;
        RECT 114.400 4.835 114.570 5.080 ;
        RECT 114.340 0.240 114.630 4.835 ;
        RECT 116.430 0.540 116.720 6.600 ;
        RECT 117.470 6.290 118.600 7.290 ;
        RECT 118.580 4.835 118.750 5.080 ;
        RECT 118.520 0.240 118.810 4.835 ;
        RECT 120.970 2.960 121.140 7.375 ;
        RECT 121.480 2.960 121.770 7.370 ;
        RECT 123.570 7.185 123.865 15.775 ;
        RECT 125.660 11.735 125.950 16.080 ;
        RECT 128.750 13.810 130.845 13.840 ;
        RECT 128.595 13.650 130.845 13.810 ;
        RECT 127.445 13.480 130.845 13.650 ;
        RECT 125.435 8.730 125.935 9.880 ;
        RECT 127.445 9.445 127.615 13.480 ;
        RECT 128.595 13.390 130.845 13.480 ;
        RECT 128.750 13.360 130.845 13.390 ;
        RECT 127.950 8.730 128.245 12.995 ;
        RECT 130.045 9.290 130.335 13.360 ;
        RECT 130.675 9.435 130.845 13.360 ;
        RECT 133.010 11.495 133.300 16.080 ;
        RECT 133.070 11.270 133.240 11.495 ;
        RECT 135.100 10.460 135.390 15.790 ;
        RECT 137.190 11.495 137.480 16.080 ;
        RECT 137.250 11.270 137.420 11.495 ;
        RECT 139.280 10.460 139.570 15.790 ;
        RECT 141.370 11.495 141.660 16.080 ;
        RECT 143.330 13.810 145.675 13.840 ;
        RECT 143.150 13.655 145.675 13.810 ;
        RECT 146.475 13.655 148.820 13.840 ;
        RECT 143.150 13.485 148.820 13.655 ;
        RECT 143.150 13.390 145.675 13.485 ;
        RECT 143.330 13.360 145.675 13.390 ;
        RECT 146.475 13.360 148.820 13.485 ;
        RECT 141.430 11.485 141.625 11.495 ;
        RECT 141.430 11.250 141.600 11.485 ;
        RECT 133.300 9.880 134.500 10.460 ;
        RECT 135.100 10.170 139.570 10.460 ;
        RECT 132.500 9.760 134.500 9.880 ;
        RECT 132.500 9.160 136.500 9.760 ;
        RECT 137.530 8.730 138.030 10.170 ;
        RECT 125.435 8.230 138.030 8.730 ;
        RECT 143.330 8.505 143.500 13.360 ;
        RECT 143.840 8.510 144.130 13.360 ;
        RECT 123.355 6.405 124.095 7.185 ;
        RECT 123.570 3.330 123.865 6.405 ;
        RECT 120.970 2.930 123.065 2.960 ;
        RECT 120.970 2.845 123.220 2.930 ;
        RECT 124.200 2.845 124.370 5.820 ;
        RECT 120.970 2.675 124.370 2.845 ;
        RECT 120.970 2.510 123.220 2.675 ;
        RECT 120.970 2.480 123.065 2.510 ;
        RECT 125.865 0.240 126.155 4.590 ;
        RECT 127.955 0.550 128.250 8.230 ;
        RECT 128.900 7.120 130.100 7.320 ;
        RECT 128.900 6.500 130.600 7.120 ;
        RECT 128.900 6.190 130.100 6.500 ;
        RECT 130.045 0.240 130.335 4.590 ;
        RECT 132.500 2.960 132.670 7.560 ;
        RECT 133.010 2.960 133.300 7.790 ;
        RECT 135.100 3.230 135.390 8.230 ;
        RECT 137.190 2.960 137.480 7.790 ;
        RECT 137.820 2.960 137.990 7.620 ;
        RECT 145.930 7.100 146.220 13.050 ;
        RECT 148.020 8.510 148.310 13.360 ;
        RECT 148.650 8.505 148.820 13.360 ;
        RECT 150.980 11.735 151.270 16.080 ;
        RECT 151.270 9.820 152.450 10.100 ;
        RECT 150.770 9.220 152.450 9.820 ;
        RECT 151.270 9.020 152.450 9.220 ;
        RECT 141.220 6.600 146.220 7.100 ;
        RECT 141.220 6.500 142.040 6.600 ;
        RECT 139.720 4.845 139.890 5.080 ;
        RECT 139.695 4.835 139.890 4.845 ;
        RECT 132.500 2.795 134.845 2.960 ;
        RECT 135.645 2.795 137.990 2.960 ;
        RECT 132.500 2.625 137.990 2.795 ;
        RECT 132.500 2.480 134.845 2.625 ;
        RECT 135.645 2.480 137.990 2.625 ;
        RECT 139.660 0.240 139.950 4.835 ;
        RECT 141.750 0.540 142.040 6.500 ;
        RECT 143.900 4.835 144.070 5.080 ;
        RECT 143.840 0.240 144.130 4.835 ;
        RECT 145.930 0.540 146.220 6.600 ;
        RECT 146.970 6.290 148.100 7.290 ;
        RECT 148.080 4.835 148.250 5.080 ;
        RECT 148.020 0.240 148.310 4.835 ;
        RECT 150.470 2.960 150.640 7.375 ;
        RECT 150.980 2.960 151.270 7.370 ;
        RECT 153.070 7.185 153.365 15.775 ;
        RECT 155.160 11.735 155.450 16.080 ;
        RECT 158.250 13.810 160.345 13.840 ;
        RECT 158.095 13.650 160.345 13.810 ;
        RECT 156.945 13.480 160.345 13.650 ;
        RECT 154.935 8.730 155.435 9.880 ;
        RECT 156.945 9.445 157.115 13.480 ;
        RECT 158.095 13.390 160.345 13.480 ;
        RECT 158.250 13.360 160.345 13.390 ;
        RECT 157.450 8.730 157.745 12.995 ;
        RECT 159.545 9.290 159.835 13.360 ;
        RECT 160.175 9.435 160.345 13.360 ;
        RECT 162.510 11.495 162.800 16.080 ;
        RECT 162.570 11.270 162.740 11.495 ;
        RECT 164.600 10.460 164.890 15.790 ;
        RECT 166.690 11.495 166.980 16.080 ;
        RECT 166.750 11.270 166.920 11.495 ;
        RECT 168.780 10.460 169.070 15.790 ;
        RECT 170.870 11.495 171.160 16.080 ;
        RECT 172.830 13.810 175.175 13.840 ;
        RECT 172.650 13.655 175.175 13.810 ;
        RECT 175.975 13.655 178.320 13.840 ;
        RECT 172.650 13.485 178.320 13.655 ;
        RECT 172.650 13.390 175.175 13.485 ;
        RECT 172.830 13.360 175.175 13.390 ;
        RECT 175.975 13.360 178.320 13.485 ;
        RECT 170.930 11.485 171.125 11.495 ;
        RECT 170.930 11.250 171.100 11.485 ;
        RECT 162.800 9.880 164.000 10.460 ;
        RECT 164.600 10.170 169.070 10.460 ;
        RECT 162.000 9.760 164.000 9.880 ;
        RECT 162.000 9.160 166.000 9.760 ;
        RECT 167.030 8.730 167.530 10.170 ;
        RECT 154.935 8.230 167.530 8.730 ;
        RECT 172.830 8.505 173.000 13.360 ;
        RECT 173.340 8.510 173.630 13.360 ;
        RECT 152.855 6.405 153.595 7.185 ;
        RECT 153.070 3.330 153.365 6.405 ;
        RECT 150.470 2.930 152.565 2.960 ;
        RECT 150.470 2.845 152.720 2.930 ;
        RECT 153.700 2.845 153.870 5.820 ;
        RECT 150.470 2.675 153.870 2.845 ;
        RECT 150.470 2.510 152.720 2.675 ;
        RECT 150.470 2.480 152.565 2.510 ;
        RECT 155.365 0.240 155.655 4.590 ;
        RECT 157.455 0.550 157.750 8.230 ;
        RECT 158.400 7.120 159.600 7.320 ;
        RECT 158.400 6.500 160.100 7.120 ;
        RECT 158.400 6.190 159.600 6.500 ;
        RECT 159.545 0.240 159.835 4.590 ;
        RECT 162.000 2.960 162.170 7.560 ;
        RECT 162.510 2.960 162.800 7.790 ;
        RECT 164.600 3.230 164.890 8.230 ;
        RECT 166.690 2.960 166.980 7.790 ;
        RECT 167.320 2.960 167.490 7.620 ;
        RECT 175.430 7.100 175.720 13.050 ;
        RECT 177.520 8.510 177.810 13.360 ;
        RECT 178.150 8.505 178.320 13.360 ;
        RECT 170.720 6.600 175.720 7.100 ;
        RECT 170.720 6.500 171.540 6.600 ;
        RECT 169.220 4.845 169.390 5.080 ;
        RECT 169.195 4.835 169.390 4.845 ;
        RECT 162.000 2.795 164.345 2.960 ;
        RECT 165.145 2.795 167.490 2.960 ;
        RECT 162.000 2.625 167.490 2.795 ;
        RECT 162.000 2.480 164.345 2.625 ;
        RECT 165.145 2.480 167.490 2.625 ;
        RECT 169.160 0.240 169.450 4.835 ;
        RECT 171.250 0.540 171.540 6.500 ;
        RECT 173.400 4.835 173.570 5.080 ;
        RECT 173.340 0.240 173.630 4.835 ;
        RECT 175.430 0.540 175.720 6.600 ;
        RECT 176.470 6.290 177.600 7.290 ;
        RECT 177.580 4.835 177.750 5.080 ;
        RECT 177.520 0.240 177.810 4.835 ;
        RECT 7.355 -0.240 9.700 0.240 ;
        RECT 10.500 -0.240 12.845 0.240 ;
        RECT 21.150 -0.240 23.495 0.240 ;
        RECT 24.550 -0.240 27.410 0.240 ;
        RECT 28.475 -0.240 30.820 0.240 ;
        RECT 36.855 -0.240 39.200 0.240 ;
        RECT 40.000 -0.240 42.345 0.240 ;
        RECT 50.650 -0.240 52.995 0.240 ;
        RECT 54.050 -0.240 56.910 0.240 ;
        RECT 57.975 -0.240 60.320 0.240 ;
        RECT 66.355 -0.240 68.700 0.240 ;
        RECT 69.500 -0.240 71.845 0.240 ;
        RECT 80.150 -0.240 82.495 0.240 ;
        RECT 83.550 -0.240 86.410 0.240 ;
        RECT 87.475 -0.240 89.820 0.240 ;
        RECT 95.855 -0.240 98.200 0.240 ;
        RECT 99.000 -0.240 101.345 0.240 ;
        RECT 109.650 -0.240 111.995 0.240 ;
        RECT 113.050 -0.240 115.910 0.240 ;
        RECT 116.975 -0.240 119.320 0.240 ;
        RECT 125.355 -0.240 127.700 0.240 ;
        RECT 128.500 -0.240 130.845 0.240 ;
        RECT 139.150 -0.240 141.495 0.240 ;
        RECT 142.550 -0.240 145.410 0.240 ;
        RECT 146.475 -0.240 148.820 0.240 ;
        RECT 154.855 -0.240 157.200 0.240 ;
        RECT 158.000 -0.240 160.345 0.240 ;
        RECT 168.650 -0.240 170.995 0.240 ;
        RECT 172.050 -0.240 174.910 0.240 ;
        RECT 175.975 -0.240 178.320 0.240 ;
      LAYER mcon ;
        RECT 18.570 37.870 19.085 38.290 ;
        RECT 19.275 37.870 19.695 38.290 ;
        RECT 19.885 37.870 20.305 38.290 ;
        RECT 20.495 37.870 20.915 38.290 ;
        RECT 21.980 37.870 22.400 38.290 ;
        RECT 22.590 37.870 23.010 38.290 ;
        RECT 23.200 37.870 23.620 38.290 ;
        RECT 23.810 37.870 24.230 38.290 ;
        RECT 24.420 37.870 24.840 38.290 ;
        RECT 25.895 37.870 26.315 38.290 ;
        RECT 26.505 37.870 26.925 38.290 ;
        RECT 27.115 37.870 27.535 38.290 ;
        RECT 27.725 37.870 28.240 38.290 ;
        RECT 36.545 37.870 36.965 38.290 ;
        RECT 37.155 37.870 37.575 38.290 ;
        RECT 37.765 37.870 38.185 38.290 ;
        RECT 38.375 37.870 38.890 38.290 ;
        RECT 39.690 37.870 40.205 38.290 ;
        RECT 40.395 37.870 40.815 38.290 ;
        RECT 41.005 37.870 41.425 38.290 ;
        RECT 41.615 37.870 42.035 38.290 ;
        RECT 48.070 37.870 48.585 38.290 ;
        RECT 48.775 37.870 49.195 38.290 ;
        RECT 49.385 37.870 49.805 38.290 ;
        RECT 49.995 37.870 50.415 38.290 ;
        RECT 51.480 37.870 51.900 38.290 ;
        RECT 52.090 37.870 52.510 38.290 ;
        RECT 52.700 37.870 53.120 38.290 ;
        RECT 53.310 37.870 53.730 38.290 ;
        RECT 53.920 37.870 54.340 38.290 ;
        RECT 55.395 37.870 55.815 38.290 ;
        RECT 56.005 37.870 56.425 38.290 ;
        RECT 56.615 37.870 57.035 38.290 ;
        RECT 57.225 37.870 57.740 38.290 ;
        RECT 66.045 37.870 66.465 38.290 ;
        RECT 66.655 37.870 67.075 38.290 ;
        RECT 67.265 37.870 67.685 38.290 ;
        RECT 67.875 37.870 68.390 38.290 ;
        RECT 69.190 37.870 69.705 38.290 ;
        RECT 69.895 37.870 70.315 38.290 ;
        RECT 70.505 37.870 70.925 38.290 ;
        RECT 71.115 37.870 71.535 38.290 ;
        RECT 77.570 37.870 78.085 38.290 ;
        RECT 78.275 37.870 78.695 38.290 ;
        RECT 78.885 37.870 79.305 38.290 ;
        RECT 79.495 37.870 79.915 38.290 ;
        RECT 80.980 37.870 81.400 38.290 ;
        RECT 81.590 37.870 82.010 38.290 ;
        RECT 82.200 37.870 82.620 38.290 ;
        RECT 82.810 37.870 83.230 38.290 ;
        RECT 83.420 37.870 83.840 38.290 ;
        RECT 84.895 37.870 85.315 38.290 ;
        RECT 85.505 37.870 85.925 38.290 ;
        RECT 86.115 37.870 86.535 38.290 ;
        RECT 86.725 37.870 87.240 38.290 ;
        RECT 95.545 37.870 95.965 38.290 ;
        RECT 96.155 37.870 96.575 38.290 ;
        RECT 96.765 37.870 97.185 38.290 ;
        RECT 97.375 37.870 97.890 38.290 ;
        RECT 98.690 37.870 99.205 38.290 ;
        RECT 99.395 37.870 99.815 38.290 ;
        RECT 100.005 37.870 100.425 38.290 ;
        RECT 100.615 37.870 101.035 38.290 ;
        RECT 107.070 37.870 107.585 38.290 ;
        RECT 107.775 37.870 108.195 38.290 ;
        RECT 108.385 37.870 108.805 38.290 ;
        RECT 108.995 37.870 109.415 38.290 ;
        RECT 110.480 37.870 110.900 38.290 ;
        RECT 111.090 37.870 111.510 38.290 ;
        RECT 111.700 37.870 112.120 38.290 ;
        RECT 112.310 37.870 112.730 38.290 ;
        RECT 112.920 37.870 113.340 38.290 ;
        RECT 114.395 37.870 114.815 38.290 ;
        RECT 115.005 37.870 115.425 38.290 ;
        RECT 115.615 37.870 116.035 38.290 ;
        RECT 116.225 37.870 116.740 38.290 ;
        RECT 125.045 37.870 125.465 38.290 ;
        RECT 125.655 37.870 126.075 38.290 ;
        RECT 126.265 37.870 126.685 38.290 ;
        RECT 126.875 37.870 127.390 38.290 ;
        RECT 128.190 37.870 128.705 38.290 ;
        RECT 128.895 37.870 129.315 38.290 ;
        RECT 129.505 37.870 129.925 38.290 ;
        RECT 130.115 37.870 130.535 38.290 ;
        RECT 136.570 37.870 137.085 38.290 ;
        RECT 137.275 37.870 137.695 38.290 ;
        RECT 137.885 37.870 138.305 38.290 ;
        RECT 138.495 37.870 138.915 38.290 ;
        RECT 139.980 37.870 140.400 38.290 ;
        RECT 140.590 37.870 141.010 38.290 ;
        RECT 141.200 37.870 141.620 38.290 ;
        RECT 141.810 37.870 142.230 38.290 ;
        RECT 142.420 37.870 142.840 38.290 ;
        RECT 143.895 37.870 144.315 38.290 ;
        RECT 144.505 37.870 144.925 38.290 ;
        RECT 145.115 37.870 145.535 38.290 ;
        RECT 145.725 37.870 146.240 38.290 ;
        RECT 154.545 37.870 154.965 38.290 ;
        RECT 155.155 37.870 155.575 38.290 ;
        RECT 155.765 37.870 156.185 38.290 ;
        RECT 156.375 37.870 156.890 38.290 ;
        RECT 157.690 37.870 158.205 38.290 ;
        RECT 158.395 37.870 158.815 38.290 ;
        RECT 159.005 37.870 159.425 38.290 ;
        RECT 159.615 37.870 160.035 38.290 ;
        RECT 19.320 30.820 20.330 31.760 ;
        RECT 29.400 35.150 29.915 35.570 ;
        RECT 30.105 35.150 30.525 35.570 ;
        RECT 30.715 35.150 31.135 35.570 ;
        RECT 31.325 35.150 31.745 35.570 ;
        RECT 32.545 35.150 32.965 35.570 ;
        RECT 33.155 35.150 33.575 35.570 ;
        RECT 33.765 35.150 34.185 35.570 ;
        RECT 34.375 35.150 34.890 35.570 ;
        RECT 25.350 30.980 26.170 31.580 ;
        RECT 3.965 29.835 4.135 30.005 ;
        RECT 4.425 29.835 4.595 30.005 ;
        RECT 4.885 29.835 5.055 30.005 ;
        RECT 5.345 29.835 5.515 30.005 ;
        RECT 5.805 29.835 5.975 30.005 ;
        RECT 8.135 29.835 8.305 30.005 ;
        RECT 8.595 29.835 8.765 30.005 ;
        RECT 9.055 29.835 9.225 30.005 ;
        RECT 6.925 28.475 7.095 28.645 ;
        RECT 3.965 27.115 4.135 27.285 ;
        RECT 4.425 27.115 4.595 27.285 ;
        RECT 4.885 27.115 5.055 27.285 ;
        RECT 5.345 27.115 5.515 27.285 ;
        RECT 5.805 27.115 5.975 27.285 ;
        RECT 8.135 27.115 8.305 27.285 ;
        RECT 8.595 27.115 8.765 27.285 ;
        RECT 9.055 27.115 9.225 27.285 ;
        RECT 36.820 30.990 37.270 31.580 ;
        RECT 37.460 30.990 38.490 31.580 ;
        RECT 44.780 35.150 45.200 35.570 ;
        RECT 45.390 35.150 45.810 35.570 ;
        RECT 46.000 35.150 46.420 35.570 ;
        RECT 43.355 30.925 43.975 31.645 ;
        RECT 30.890 28.320 31.490 28.920 ;
        RECT 31.690 28.320 32.290 28.920 ;
        RECT 32.490 28.320 33.090 28.920 ;
        RECT 33.290 28.230 33.990 28.920 ;
        RECT 34.190 28.230 34.830 28.860 ;
        RECT 18.570 24.270 19.085 24.690 ;
        RECT 19.275 24.270 19.695 24.690 ;
        RECT 19.885 24.270 20.305 24.690 ;
        RECT 20.495 24.270 20.915 24.690 ;
        RECT 21.895 24.270 22.315 24.690 ;
        RECT 22.505 24.270 22.925 24.690 ;
        RECT 23.115 24.270 23.535 24.690 ;
        RECT 23.725 24.270 24.240 24.690 ;
        RECT 37.155 24.270 37.575 24.690 ;
        RECT 37.765 24.270 38.185 24.690 ;
        RECT 38.375 24.270 38.795 24.690 ;
        RECT 41.455 28.260 41.955 28.860 ;
        RECT 48.820 30.820 49.830 31.760 ;
        RECT 58.900 35.150 59.415 35.570 ;
        RECT 59.605 35.150 60.025 35.570 ;
        RECT 60.215 35.150 60.635 35.570 ;
        RECT 60.825 35.150 61.245 35.570 ;
        RECT 62.045 35.150 62.465 35.570 ;
        RECT 62.655 35.150 63.075 35.570 ;
        RECT 63.265 35.150 63.685 35.570 ;
        RECT 63.875 35.150 64.390 35.570 ;
        RECT 54.850 30.980 55.670 31.580 ;
        RECT 44.520 28.310 45.470 28.810 ;
        RECT 45.670 28.310 46.070 28.810 ;
        RECT 66.320 30.990 66.770 31.580 ;
        RECT 66.960 30.990 67.990 31.580 ;
        RECT 74.280 35.150 74.700 35.570 ;
        RECT 74.890 35.150 75.310 35.570 ;
        RECT 75.500 35.150 75.920 35.570 ;
        RECT 72.855 30.925 73.475 31.645 ;
        RECT 60.390 28.320 60.990 28.920 ;
        RECT 61.190 28.320 61.790 28.920 ;
        RECT 61.990 28.320 62.590 28.920 ;
        RECT 62.790 28.230 63.490 28.920 ;
        RECT 63.690 28.230 64.330 28.860 ;
        RECT 48.070 24.270 48.585 24.690 ;
        RECT 48.775 24.270 49.195 24.690 ;
        RECT 49.385 24.270 49.805 24.690 ;
        RECT 49.995 24.270 50.415 24.690 ;
        RECT 51.395 24.270 51.815 24.690 ;
        RECT 52.005 24.270 52.425 24.690 ;
        RECT 52.615 24.270 53.035 24.690 ;
        RECT 53.225 24.270 53.740 24.690 ;
        RECT 66.655 24.270 67.075 24.690 ;
        RECT 67.265 24.270 67.685 24.690 ;
        RECT 67.875 24.270 68.295 24.690 ;
        RECT 70.955 28.260 71.455 28.860 ;
        RECT 78.320 30.820 79.330 31.760 ;
        RECT 88.400 35.150 88.915 35.570 ;
        RECT 89.105 35.150 89.525 35.570 ;
        RECT 89.715 35.150 90.135 35.570 ;
        RECT 90.325 35.150 90.745 35.570 ;
        RECT 91.545 35.150 91.965 35.570 ;
        RECT 92.155 35.150 92.575 35.570 ;
        RECT 92.765 35.150 93.185 35.570 ;
        RECT 93.375 35.150 93.890 35.570 ;
        RECT 84.350 30.980 85.170 31.580 ;
        RECT 74.020 28.310 74.970 28.810 ;
        RECT 75.170 28.310 75.570 28.810 ;
        RECT 95.820 30.990 96.270 31.580 ;
        RECT 96.460 30.990 97.490 31.580 ;
        RECT 103.780 35.150 104.200 35.570 ;
        RECT 104.390 35.150 104.810 35.570 ;
        RECT 105.000 35.150 105.420 35.570 ;
        RECT 102.355 30.925 102.975 31.645 ;
        RECT 89.890 28.320 90.490 28.920 ;
        RECT 90.690 28.320 91.290 28.920 ;
        RECT 91.490 28.320 92.090 28.920 ;
        RECT 92.290 28.230 92.990 28.920 ;
        RECT 93.190 28.230 93.830 28.860 ;
        RECT 77.570 24.270 78.085 24.690 ;
        RECT 78.275 24.270 78.695 24.690 ;
        RECT 78.885 24.270 79.305 24.690 ;
        RECT 79.495 24.270 79.915 24.690 ;
        RECT 80.895 24.270 81.315 24.690 ;
        RECT 81.505 24.270 81.925 24.690 ;
        RECT 82.115 24.270 82.535 24.690 ;
        RECT 82.725 24.270 83.240 24.690 ;
        RECT 96.155 24.270 96.575 24.690 ;
        RECT 96.765 24.270 97.185 24.690 ;
        RECT 97.375 24.270 97.795 24.690 ;
        RECT 100.455 28.260 100.955 28.860 ;
        RECT 107.820 30.820 108.830 31.760 ;
        RECT 117.900 35.150 118.415 35.570 ;
        RECT 118.605 35.150 119.025 35.570 ;
        RECT 119.215 35.150 119.635 35.570 ;
        RECT 119.825 35.150 120.245 35.570 ;
        RECT 121.045 35.150 121.465 35.570 ;
        RECT 121.655 35.150 122.075 35.570 ;
        RECT 122.265 35.150 122.685 35.570 ;
        RECT 122.875 35.150 123.390 35.570 ;
        RECT 113.850 30.980 114.670 31.580 ;
        RECT 103.520 28.310 104.470 28.810 ;
        RECT 104.670 28.310 105.070 28.810 ;
        RECT 125.320 30.990 125.770 31.580 ;
        RECT 125.960 30.990 126.990 31.580 ;
        RECT 133.280 35.150 133.700 35.570 ;
        RECT 133.890 35.150 134.310 35.570 ;
        RECT 134.500 35.150 134.920 35.570 ;
        RECT 131.855 30.925 132.475 31.645 ;
        RECT 119.390 28.320 119.990 28.920 ;
        RECT 120.190 28.320 120.790 28.920 ;
        RECT 120.990 28.320 121.590 28.920 ;
        RECT 121.790 28.230 122.490 28.920 ;
        RECT 122.690 28.230 123.330 28.860 ;
        RECT 107.070 24.270 107.585 24.690 ;
        RECT 107.775 24.270 108.195 24.690 ;
        RECT 108.385 24.270 108.805 24.690 ;
        RECT 108.995 24.270 109.415 24.690 ;
        RECT 110.395 24.270 110.815 24.690 ;
        RECT 111.005 24.270 111.425 24.690 ;
        RECT 111.615 24.270 112.035 24.690 ;
        RECT 112.225 24.270 112.740 24.690 ;
        RECT 125.655 24.270 126.075 24.690 ;
        RECT 126.265 24.270 126.685 24.690 ;
        RECT 126.875 24.270 127.295 24.690 ;
        RECT 129.955 28.260 130.455 28.860 ;
        RECT 137.320 30.820 138.330 31.760 ;
        RECT 147.400 35.150 147.915 35.570 ;
        RECT 148.105 35.150 148.525 35.570 ;
        RECT 148.715 35.150 149.135 35.570 ;
        RECT 149.325 35.150 149.745 35.570 ;
        RECT 150.545 35.150 150.965 35.570 ;
        RECT 151.155 35.150 151.575 35.570 ;
        RECT 151.765 35.150 152.185 35.570 ;
        RECT 152.375 35.150 152.890 35.570 ;
        RECT 143.350 30.980 144.170 31.580 ;
        RECT 133.020 28.310 133.970 28.810 ;
        RECT 134.170 28.310 134.570 28.810 ;
        RECT 154.820 30.990 155.270 31.580 ;
        RECT 155.460 30.990 156.490 31.580 ;
        RECT 162.780 35.150 163.200 35.570 ;
        RECT 163.390 35.150 163.810 35.570 ;
        RECT 164.000 35.150 164.420 35.570 ;
        RECT 161.355 30.925 161.975 31.645 ;
        RECT 148.890 28.320 149.490 28.920 ;
        RECT 149.690 28.320 150.290 28.920 ;
        RECT 150.490 28.320 151.090 28.920 ;
        RECT 151.290 28.230 151.990 28.920 ;
        RECT 152.190 28.230 152.830 28.860 ;
        RECT 136.570 24.270 137.085 24.690 ;
        RECT 137.275 24.270 137.695 24.690 ;
        RECT 137.885 24.270 138.305 24.690 ;
        RECT 138.495 24.270 138.915 24.690 ;
        RECT 139.895 24.270 140.315 24.690 ;
        RECT 140.505 24.270 140.925 24.690 ;
        RECT 141.115 24.270 141.535 24.690 ;
        RECT 141.725 24.270 142.240 24.690 ;
        RECT 155.155 24.270 155.575 24.690 ;
        RECT 155.765 24.270 156.185 24.690 ;
        RECT 156.375 24.270 156.795 24.690 ;
        RECT 159.455 28.260 159.955 28.860 ;
        RECT 162.520 28.310 163.470 28.810 ;
        RECT 163.670 28.310 164.070 28.810 ;
        RECT 25.220 21.550 25.735 21.970 ;
        RECT 25.925 21.550 26.345 21.970 ;
        RECT 26.535 21.550 26.955 21.970 ;
        RECT 27.145 21.550 27.565 21.970 ;
        RECT 28.620 21.550 29.040 21.970 ;
        RECT 29.230 21.550 29.650 21.970 ;
        RECT 29.840 21.550 30.260 21.970 ;
        RECT 30.450 21.550 30.870 21.970 ;
        RECT 31.060 21.550 31.480 21.970 ;
        RECT 32.545 21.550 32.965 21.970 ;
        RECT 33.155 21.550 33.575 21.970 ;
        RECT 33.765 21.550 34.185 21.970 ;
        RECT 34.375 21.550 34.890 21.970 ;
        RECT 41.640 21.550 42.050 21.970 ;
        RECT 42.250 21.550 42.660 21.970 ;
        RECT 42.860 21.550 43.275 21.970 ;
        RECT 44.685 21.550 45.105 21.970 ;
        RECT 45.295 21.550 45.715 21.970 ;
        RECT 45.905 21.550 46.420 21.970 ;
        RECT 54.720 21.550 55.235 21.970 ;
        RECT 55.425 21.550 55.845 21.970 ;
        RECT 56.035 21.550 56.455 21.970 ;
        RECT 56.645 21.550 57.065 21.970 ;
        RECT 58.120 21.550 58.540 21.970 ;
        RECT 58.730 21.550 59.150 21.970 ;
        RECT 59.340 21.550 59.760 21.970 ;
        RECT 59.950 21.550 60.370 21.970 ;
        RECT 60.560 21.550 60.980 21.970 ;
        RECT 62.045 21.550 62.465 21.970 ;
        RECT 62.655 21.550 63.075 21.970 ;
        RECT 63.265 21.550 63.685 21.970 ;
        RECT 63.875 21.550 64.390 21.970 ;
        RECT 71.140 21.550 71.550 21.970 ;
        RECT 71.750 21.550 72.160 21.970 ;
        RECT 72.360 21.550 72.775 21.970 ;
        RECT 74.185 21.550 74.605 21.970 ;
        RECT 74.795 21.550 75.215 21.970 ;
        RECT 75.405 21.550 75.920 21.970 ;
        RECT 84.220 21.550 84.735 21.970 ;
        RECT 84.925 21.550 85.345 21.970 ;
        RECT 85.535 21.550 85.955 21.970 ;
        RECT 86.145 21.550 86.565 21.970 ;
        RECT 87.620 21.550 88.040 21.970 ;
        RECT 88.230 21.550 88.650 21.970 ;
        RECT 88.840 21.550 89.260 21.970 ;
        RECT 89.450 21.550 89.870 21.970 ;
        RECT 90.060 21.550 90.480 21.970 ;
        RECT 91.545 21.550 91.965 21.970 ;
        RECT 92.155 21.550 92.575 21.970 ;
        RECT 92.765 21.550 93.185 21.970 ;
        RECT 93.375 21.550 93.890 21.970 ;
        RECT 100.640 21.550 101.050 21.970 ;
        RECT 101.250 21.550 101.660 21.970 ;
        RECT 101.860 21.550 102.275 21.970 ;
        RECT 103.685 21.550 104.105 21.970 ;
        RECT 104.295 21.550 104.715 21.970 ;
        RECT 104.905 21.550 105.420 21.970 ;
        RECT 113.720 21.550 114.235 21.970 ;
        RECT 114.425 21.550 114.845 21.970 ;
        RECT 115.035 21.550 115.455 21.970 ;
        RECT 115.645 21.550 116.065 21.970 ;
        RECT 117.120 21.550 117.540 21.970 ;
        RECT 117.730 21.550 118.150 21.970 ;
        RECT 118.340 21.550 118.760 21.970 ;
        RECT 118.950 21.550 119.370 21.970 ;
        RECT 119.560 21.550 119.980 21.970 ;
        RECT 121.045 21.550 121.465 21.970 ;
        RECT 121.655 21.550 122.075 21.970 ;
        RECT 122.265 21.550 122.685 21.970 ;
        RECT 122.875 21.550 123.390 21.970 ;
        RECT 130.140 21.550 130.550 21.970 ;
        RECT 130.750 21.550 131.160 21.970 ;
        RECT 131.360 21.550 131.775 21.970 ;
        RECT 133.185 21.550 133.605 21.970 ;
        RECT 133.795 21.550 134.215 21.970 ;
        RECT 134.405 21.550 134.920 21.970 ;
        RECT 143.220 21.550 143.735 21.970 ;
        RECT 143.925 21.550 144.345 21.970 ;
        RECT 144.535 21.550 144.955 21.970 ;
        RECT 145.145 21.550 145.565 21.970 ;
        RECT 146.620 21.550 147.040 21.970 ;
        RECT 147.230 21.550 147.650 21.970 ;
        RECT 147.840 21.550 148.260 21.970 ;
        RECT 148.450 21.550 148.870 21.970 ;
        RECT 149.060 21.550 149.480 21.970 ;
        RECT 150.545 21.550 150.965 21.970 ;
        RECT 151.155 21.550 151.575 21.970 ;
        RECT 151.765 21.550 152.185 21.970 ;
        RECT 152.375 21.550 152.890 21.970 ;
        RECT 159.640 21.550 160.050 21.970 ;
        RECT 160.250 21.550 160.660 21.970 ;
        RECT 160.860 21.550 161.275 21.970 ;
        RECT 162.685 21.550 163.105 21.970 ;
        RECT 163.295 21.550 163.715 21.970 ;
        RECT 163.905 21.550 164.420 21.970 ;
        RECT 3.675 16.110 4.095 16.530 ;
        RECT 4.285 16.110 4.705 16.530 ;
        RECT 4.895 16.110 5.315 16.530 ;
        RECT 6.730 16.110 7.140 16.530 ;
        RECT 7.340 16.110 7.750 16.530 ;
        RECT 7.950 16.110 8.460 16.530 ;
        RECT 14.500 16.110 15.015 16.530 ;
        RECT 15.205 16.110 15.625 16.530 ;
        RECT 15.815 16.110 16.235 16.530 ;
        RECT 16.425 16.110 16.845 16.530 ;
        RECT 17.910 16.110 18.330 16.530 ;
        RECT 18.520 16.110 18.940 16.530 ;
        RECT 19.130 16.110 19.550 16.530 ;
        RECT 19.740 16.110 20.160 16.530 ;
        RECT 20.350 16.110 20.770 16.530 ;
        RECT 21.825 16.110 22.245 16.530 ;
        RECT 22.435 16.110 22.855 16.530 ;
        RECT 23.045 16.110 23.465 16.530 ;
        RECT 23.655 16.110 24.170 16.530 ;
        RECT 33.175 16.110 33.595 16.530 ;
        RECT 33.785 16.110 34.205 16.530 ;
        RECT 34.395 16.110 34.815 16.530 ;
        RECT 36.230 16.110 36.640 16.530 ;
        RECT 36.840 16.110 37.250 16.530 ;
        RECT 37.450 16.110 37.960 16.530 ;
        RECT 44.000 16.110 44.515 16.530 ;
        RECT 44.705 16.110 45.125 16.530 ;
        RECT 45.315 16.110 45.735 16.530 ;
        RECT 45.925 16.110 46.345 16.530 ;
        RECT 47.410 16.110 47.830 16.530 ;
        RECT 48.020 16.110 48.440 16.530 ;
        RECT 48.630 16.110 49.050 16.530 ;
        RECT 49.240 16.110 49.660 16.530 ;
        RECT 49.850 16.110 50.270 16.530 ;
        RECT 51.325 16.110 51.745 16.530 ;
        RECT 51.935 16.110 52.355 16.530 ;
        RECT 52.545 16.110 52.965 16.530 ;
        RECT 53.155 16.110 53.670 16.530 ;
        RECT 62.675 16.110 63.095 16.530 ;
        RECT 63.285 16.110 63.705 16.530 ;
        RECT 63.895 16.110 64.315 16.530 ;
        RECT 65.730 16.110 66.140 16.530 ;
        RECT 66.340 16.110 66.750 16.530 ;
        RECT 66.950 16.110 67.460 16.530 ;
        RECT 73.500 16.110 74.015 16.530 ;
        RECT 74.205 16.110 74.625 16.530 ;
        RECT 74.815 16.110 75.235 16.530 ;
        RECT 75.425 16.110 75.845 16.530 ;
        RECT 76.910 16.110 77.330 16.530 ;
        RECT 77.520 16.110 77.940 16.530 ;
        RECT 78.130 16.110 78.550 16.530 ;
        RECT 78.740 16.110 79.160 16.530 ;
        RECT 79.350 16.110 79.770 16.530 ;
        RECT 80.825 16.110 81.245 16.530 ;
        RECT 81.435 16.110 81.855 16.530 ;
        RECT 82.045 16.110 82.465 16.530 ;
        RECT 82.655 16.110 83.170 16.530 ;
        RECT 92.175 16.110 92.595 16.530 ;
        RECT 92.785 16.110 93.205 16.530 ;
        RECT 93.395 16.110 93.815 16.530 ;
        RECT 95.230 16.110 95.640 16.530 ;
        RECT 95.840 16.110 96.250 16.530 ;
        RECT 96.450 16.110 96.960 16.530 ;
        RECT 103.000 16.110 103.515 16.530 ;
        RECT 103.705 16.110 104.125 16.530 ;
        RECT 104.315 16.110 104.735 16.530 ;
        RECT 104.925 16.110 105.345 16.530 ;
        RECT 106.410 16.110 106.830 16.530 ;
        RECT 107.020 16.110 107.440 16.530 ;
        RECT 107.630 16.110 108.050 16.530 ;
        RECT 108.240 16.110 108.660 16.530 ;
        RECT 108.850 16.110 109.270 16.530 ;
        RECT 110.325 16.110 110.745 16.530 ;
        RECT 110.935 16.110 111.355 16.530 ;
        RECT 111.545 16.110 111.965 16.530 ;
        RECT 112.155 16.110 112.670 16.530 ;
        RECT 121.675 16.110 122.095 16.530 ;
        RECT 122.285 16.110 122.705 16.530 ;
        RECT 122.895 16.110 123.315 16.530 ;
        RECT 124.730 16.110 125.140 16.530 ;
        RECT 125.340 16.110 125.750 16.530 ;
        RECT 125.950 16.110 126.460 16.530 ;
        RECT 132.500 16.110 133.015 16.530 ;
        RECT 133.205 16.110 133.625 16.530 ;
        RECT 133.815 16.110 134.235 16.530 ;
        RECT 134.425 16.110 134.845 16.530 ;
        RECT 135.910 16.110 136.330 16.530 ;
        RECT 136.520 16.110 136.940 16.530 ;
        RECT 137.130 16.110 137.550 16.530 ;
        RECT 137.740 16.110 138.160 16.530 ;
        RECT 138.350 16.110 138.770 16.530 ;
        RECT 139.825 16.110 140.245 16.530 ;
        RECT 140.435 16.110 140.855 16.530 ;
        RECT 141.045 16.110 141.465 16.530 ;
        RECT 141.655 16.110 142.170 16.530 ;
        RECT 151.175 16.110 151.595 16.530 ;
        RECT 151.785 16.110 152.205 16.530 ;
        RECT 152.395 16.110 152.815 16.530 ;
        RECT 154.230 16.110 154.640 16.530 ;
        RECT 154.840 16.110 155.250 16.530 ;
        RECT 155.450 16.110 155.960 16.530 ;
        RECT 162.000 16.110 162.515 16.530 ;
        RECT 162.705 16.110 163.125 16.530 ;
        RECT 163.315 16.110 163.735 16.530 ;
        RECT 163.925 16.110 164.345 16.530 ;
        RECT 165.410 16.110 165.830 16.530 ;
        RECT 166.020 16.110 166.440 16.530 ;
        RECT 166.630 16.110 167.050 16.530 ;
        RECT 167.240 16.110 167.660 16.530 ;
        RECT 167.850 16.110 168.270 16.530 ;
        RECT 169.325 16.110 169.745 16.530 ;
        RECT 169.935 16.110 170.355 16.530 ;
        RECT 170.545 16.110 170.965 16.530 ;
        RECT 171.155 16.110 171.670 16.530 ;
        RECT 3.320 9.270 3.720 9.770 ;
        RECT 3.920 9.270 4.870 9.770 ;
        RECT 7.435 9.220 7.935 9.820 ;
        RECT 11.205 13.390 11.625 13.810 ;
        RECT 11.815 13.390 12.235 13.810 ;
        RECT 12.425 13.390 12.845 13.810 ;
        RECT 25.855 13.390 26.275 13.810 ;
        RECT 26.465 13.390 26.885 13.810 ;
        RECT 27.075 13.390 27.495 13.810 ;
        RECT 28.475 13.390 28.895 13.810 ;
        RECT 29.085 13.390 29.505 13.810 ;
        RECT 29.695 13.390 30.115 13.810 ;
        RECT 30.305 13.390 30.820 13.810 ;
        RECT 14.560 9.220 15.200 9.850 ;
        RECT 15.400 9.160 16.100 9.850 ;
        RECT 16.300 9.160 16.900 9.760 ;
        RECT 17.100 9.160 17.700 9.760 ;
        RECT 17.900 9.160 18.500 9.760 ;
        RECT 5.415 6.435 6.035 7.155 ;
        RECT 3.580 2.510 4.000 2.930 ;
        RECT 4.190 2.510 4.610 2.930 ;
        RECT 4.800 2.510 5.220 2.930 ;
        RECT 10.900 6.500 11.930 7.090 ;
        RECT 12.120 6.500 12.570 7.090 ;
        RECT 32.820 9.270 33.220 9.770 ;
        RECT 33.420 9.270 34.370 9.770 ;
        RECT 14.500 2.510 15.015 2.930 ;
        RECT 15.205 2.510 15.625 2.930 ;
        RECT 15.815 2.510 16.235 2.930 ;
        RECT 16.425 2.510 16.845 2.930 ;
        RECT 17.645 2.510 18.065 2.930 ;
        RECT 18.255 2.510 18.675 2.930 ;
        RECT 18.865 2.510 19.285 2.930 ;
        RECT 19.475 2.510 19.990 2.930 ;
        RECT 29.060 6.320 30.070 7.260 ;
        RECT 36.935 9.220 37.435 9.820 ;
        RECT 40.705 13.390 41.125 13.810 ;
        RECT 41.315 13.390 41.735 13.810 ;
        RECT 41.925 13.390 42.345 13.810 ;
        RECT 55.355 13.390 55.775 13.810 ;
        RECT 55.965 13.390 56.385 13.810 ;
        RECT 56.575 13.390 56.995 13.810 ;
        RECT 57.975 13.390 58.395 13.810 ;
        RECT 58.585 13.390 59.005 13.810 ;
        RECT 59.195 13.390 59.615 13.810 ;
        RECT 59.805 13.390 60.320 13.810 ;
        RECT 44.060 9.220 44.700 9.850 ;
        RECT 44.900 9.160 45.600 9.850 ;
        RECT 45.800 9.160 46.400 9.760 ;
        RECT 46.600 9.160 47.200 9.760 ;
        RECT 47.400 9.160 48.000 9.760 ;
        RECT 34.915 6.435 35.535 7.155 ;
        RECT 33.080 2.510 33.500 2.930 ;
        RECT 33.690 2.510 34.110 2.930 ;
        RECT 34.300 2.510 34.720 2.930 ;
        RECT 40.400 6.500 41.430 7.090 ;
        RECT 41.620 6.500 42.070 7.090 ;
        RECT 62.320 9.270 62.720 9.770 ;
        RECT 62.920 9.270 63.870 9.770 ;
        RECT 44.000 2.510 44.515 2.930 ;
        RECT 44.705 2.510 45.125 2.930 ;
        RECT 45.315 2.510 45.735 2.930 ;
        RECT 45.925 2.510 46.345 2.930 ;
        RECT 47.145 2.510 47.565 2.930 ;
        RECT 47.755 2.510 48.175 2.930 ;
        RECT 48.365 2.510 48.785 2.930 ;
        RECT 48.975 2.510 49.490 2.930 ;
        RECT 58.560 6.320 59.570 7.260 ;
        RECT 66.435 9.220 66.935 9.820 ;
        RECT 70.205 13.390 70.625 13.810 ;
        RECT 70.815 13.390 71.235 13.810 ;
        RECT 71.425 13.390 71.845 13.810 ;
        RECT 84.855 13.390 85.275 13.810 ;
        RECT 85.465 13.390 85.885 13.810 ;
        RECT 86.075 13.390 86.495 13.810 ;
        RECT 87.475 13.390 87.895 13.810 ;
        RECT 88.085 13.390 88.505 13.810 ;
        RECT 88.695 13.390 89.115 13.810 ;
        RECT 89.305 13.390 89.820 13.810 ;
        RECT 73.560 9.220 74.200 9.850 ;
        RECT 74.400 9.160 75.100 9.850 ;
        RECT 75.300 9.160 75.900 9.760 ;
        RECT 76.100 9.160 76.700 9.760 ;
        RECT 76.900 9.160 77.500 9.760 ;
        RECT 64.415 6.435 65.035 7.155 ;
        RECT 62.580 2.510 63.000 2.930 ;
        RECT 63.190 2.510 63.610 2.930 ;
        RECT 63.800 2.510 64.220 2.930 ;
        RECT 69.900 6.500 70.930 7.090 ;
        RECT 71.120 6.500 71.570 7.090 ;
        RECT 91.820 9.270 92.220 9.770 ;
        RECT 92.420 9.270 93.370 9.770 ;
        RECT 73.500 2.510 74.015 2.930 ;
        RECT 74.205 2.510 74.625 2.930 ;
        RECT 74.815 2.510 75.235 2.930 ;
        RECT 75.425 2.510 75.845 2.930 ;
        RECT 76.645 2.510 77.065 2.930 ;
        RECT 77.255 2.510 77.675 2.930 ;
        RECT 77.865 2.510 78.285 2.930 ;
        RECT 78.475 2.510 78.990 2.930 ;
        RECT 88.060 6.320 89.070 7.260 ;
        RECT 95.935 9.220 96.435 9.820 ;
        RECT 99.705 13.390 100.125 13.810 ;
        RECT 100.315 13.390 100.735 13.810 ;
        RECT 100.925 13.390 101.345 13.810 ;
        RECT 114.355 13.390 114.775 13.810 ;
        RECT 114.965 13.390 115.385 13.810 ;
        RECT 115.575 13.390 115.995 13.810 ;
        RECT 116.975 13.390 117.395 13.810 ;
        RECT 117.585 13.390 118.005 13.810 ;
        RECT 118.195 13.390 118.615 13.810 ;
        RECT 118.805 13.390 119.320 13.810 ;
        RECT 103.060 9.220 103.700 9.850 ;
        RECT 103.900 9.160 104.600 9.850 ;
        RECT 104.800 9.160 105.400 9.760 ;
        RECT 105.600 9.160 106.200 9.760 ;
        RECT 106.400 9.160 107.000 9.760 ;
        RECT 93.915 6.435 94.535 7.155 ;
        RECT 92.080 2.510 92.500 2.930 ;
        RECT 92.690 2.510 93.110 2.930 ;
        RECT 93.300 2.510 93.720 2.930 ;
        RECT 99.400 6.500 100.430 7.090 ;
        RECT 100.620 6.500 101.070 7.090 ;
        RECT 121.320 9.270 121.720 9.770 ;
        RECT 121.920 9.270 122.870 9.770 ;
        RECT 103.000 2.510 103.515 2.930 ;
        RECT 103.705 2.510 104.125 2.930 ;
        RECT 104.315 2.510 104.735 2.930 ;
        RECT 104.925 2.510 105.345 2.930 ;
        RECT 106.145 2.510 106.565 2.930 ;
        RECT 106.755 2.510 107.175 2.930 ;
        RECT 107.365 2.510 107.785 2.930 ;
        RECT 107.975 2.510 108.490 2.930 ;
        RECT 117.560 6.320 118.570 7.260 ;
        RECT 125.435 9.220 125.935 9.820 ;
        RECT 129.205 13.390 129.625 13.810 ;
        RECT 129.815 13.390 130.235 13.810 ;
        RECT 130.425 13.390 130.845 13.810 ;
        RECT 143.855 13.390 144.275 13.810 ;
        RECT 144.465 13.390 144.885 13.810 ;
        RECT 145.075 13.390 145.495 13.810 ;
        RECT 146.475 13.390 146.895 13.810 ;
        RECT 147.085 13.390 147.505 13.810 ;
        RECT 147.695 13.390 148.115 13.810 ;
        RECT 148.305 13.390 148.820 13.810 ;
        RECT 132.560 9.220 133.200 9.850 ;
        RECT 133.400 9.160 134.100 9.850 ;
        RECT 134.300 9.160 134.900 9.760 ;
        RECT 135.100 9.160 135.700 9.760 ;
        RECT 135.900 9.160 136.500 9.760 ;
        RECT 123.415 6.435 124.035 7.155 ;
        RECT 121.580 2.510 122.000 2.930 ;
        RECT 122.190 2.510 122.610 2.930 ;
        RECT 122.800 2.510 123.220 2.930 ;
        RECT 128.900 6.500 129.930 7.090 ;
        RECT 130.120 6.500 130.570 7.090 ;
        RECT 150.820 9.270 151.220 9.770 ;
        RECT 151.420 9.270 152.370 9.770 ;
        RECT 132.500 2.510 133.015 2.930 ;
        RECT 133.205 2.510 133.625 2.930 ;
        RECT 133.815 2.510 134.235 2.930 ;
        RECT 134.425 2.510 134.845 2.930 ;
        RECT 135.645 2.510 136.065 2.930 ;
        RECT 136.255 2.510 136.675 2.930 ;
        RECT 136.865 2.510 137.285 2.930 ;
        RECT 137.475 2.510 137.990 2.930 ;
        RECT 147.060 6.320 148.070 7.260 ;
        RECT 154.935 9.220 155.435 9.820 ;
        RECT 158.705 13.390 159.125 13.810 ;
        RECT 159.315 13.390 159.735 13.810 ;
        RECT 159.925 13.390 160.345 13.810 ;
        RECT 173.355 13.390 173.775 13.810 ;
        RECT 173.965 13.390 174.385 13.810 ;
        RECT 174.575 13.390 174.995 13.810 ;
        RECT 175.975 13.390 176.395 13.810 ;
        RECT 176.585 13.390 177.005 13.810 ;
        RECT 177.195 13.390 177.615 13.810 ;
        RECT 177.805 13.390 178.320 13.810 ;
        RECT 162.060 9.220 162.700 9.850 ;
        RECT 162.900 9.160 163.600 9.850 ;
        RECT 163.800 9.160 164.400 9.760 ;
        RECT 164.600 9.160 165.200 9.760 ;
        RECT 165.400 9.160 166.000 9.760 ;
        RECT 152.915 6.435 153.535 7.155 ;
        RECT 151.080 2.510 151.500 2.930 ;
        RECT 151.690 2.510 152.110 2.930 ;
        RECT 152.300 2.510 152.720 2.930 ;
        RECT 158.400 6.500 159.430 7.090 ;
        RECT 159.620 6.500 160.070 7.090 ;
        RECT 162.000 2.510 162.515 2.930 ;
        RECT 162.705 2.510 163.125 2.930 ;
        RECT 163.315 2.510 163.735 2.930 ;
        RECT 163.925 2.510 164.345 2.930 ;
        RECT 165.145 2.510 165.565 2.930 ;
        RECT 165.755 2.510 166.175 2.930 ;
        RECT 166.365 2.510 166.785 2.930 ;
        RECT 166.975 2.510 167.490 2.930 ;
        RECT 176.560 6.320 177.570 7.260 ;
        RECT 7.355 -0.210 7.775 0.210 ;
        RECT 7.965 -0.210 8.385 0.210 ;
        RECT 8.575 -0.210 8.995 0.210 ;
        RECT 9.185 -0.210 9.700 0.210 ;
        RECT 10.500 -0.210 11.015 0.210 ;
        RECT 11.205 -0.210 11.625 0.210 ;
        RECT 11.815 -0.210 12.235 0.210 ;
        RECT 12.425 -0.210 12.845 0.210 ;
        RECT 21.150 -0.210 21.665 0.210 ;
        RECT 21.855 -0.210 22.275 0.210 ;
        RECT 22.465 -0.210 22.885 0.210 ;
        RECT 23.075 -0.210 23.495 0.210 ;
        RECT 24.550 -0.210 24.970 0.210 ;
        RECT 25.160 -0.210 25.580 0.210 ;
        RECT 25.770 -0.210 26.190 0.210 ;
        RECT 26.380 -0.210 26.800 0.210 ;
        RECT 26.990 -0.210 27.410 0.210 ;
        RECT 28.475 -0.210 28.895 0.210 ;
        RECT 29.085 -0.210 29.505 0.210 ;
        RECT 29.695 -0.210 30.115 0.210 ;
        RECT 30.305 -0.210 30.820 0.210 ;
        RECT 36.855 -0.210 37.275 0.210 ;
        RECT 37.465 -0.210 37.885 0.210 ;
        RECT 38.075 -0.210 38.495 0.210 ;
        RECT 38.685 -0.210 39.200 0.210 ;
        RECT 40.000 -0.210 40.515 0.210 ;
        RECT 40.705 -0.210 41.125 0.210 ;
        RECT 41.315 -0.210 41.735 0.210 ;
        RECT 41.925 -0.210 42.345 0.210 ;
        RECT 50.650 -0.210 51.165 0.210 ;
        RECT 51.355 -0.210 51.775 0.210 ;
        RECT 51.965 -0.210 52.385 0.210 ;
        RECT 52.575 -0.210 52.995 0.210 ;
        RECT 54.050 -0.210 54.470 0.210 ;
        RECT 54.660 -0.210 55.080 0.210 ;
        RECT 55.270 -0.210 55.690 0.210 ;
        RECT 55.880 -0.210 56.300 0.210 ;
        RECT 56.490 -0.210 56.910 0.210 ;
        RECT 57.975 -0.210 58.395 0.210 ;
        RECT 58.585 -0.210 59.005 0.210 ;
        RECT 59.195 -0.210 59.615 0.210 ;
        RECT 59.805 -0.210 60.320 0.210 ;
        RECT 66.355 -0.210 66.775 0.210 ;
        RECT 66.965 -0.210 67.385 0.210 ;
        RECT 67.575 -0.210 67.995 0.210 ;
        RECT 68.185 -0.210 68.700 0.210 ;
        RECT 69.500 -0.210 70.015 0.210 ;
        RECT 70.205 -0.210 70.625 0.210 ;
        RECT 70.815 -0.210 71.235 0.210 ;
        RECT 71.425 -0.210 71.845 0.210 ;
        RECT 80.150 -0.210 80.665 0.210 ;
        RECT 80.855 -0.210 81.275 0.210 ;
        RECT 81.465 -0.210 81.885 0.210 ;
        RECT 82.075 -0.210 82.495 0.210 ;
        RECT 83.550 -0.210 83.970 0.210 ;
        RECT 84.160 -0.210 84.580 0.210 ;
        RECT 84.770 -0.210 85.190 0.210 ;
        RECT 85.380 -0.210 85.800 0.210 ;
        RECT 85.990 -0.210 86.410 0.210 ;
        RECT 87.475 -0.210 87.895 0.210 ;
        RECT 88.085 -0.210 88.505 0.210 ;
        RECT 88.695 -0.210 89.115 0.210 ;
        RECT 89.305 -0.210 89.820 0.210 ;
        RECT 95.855 -0.210 96.275 0.210 ;
        RECT 96.465 -0.210 96.885 0.210 ;
        RECT 97.075 -0.210 97.495 0.210 ;
        RECT 97.685 -0.210 98.200 0.210 ;
        RECT 99.000 -0.210 99.515 0.210 ;
        RECT 99.705 -0.210 100.125 0.210 ;
        RECT 100.315 -0.210 100.735 0.210 ;
        RECT 100.925 -0.210 101.345 0.210 ;
        RECT 109.650 -0.210 110.165 0.210 ;
        RECT 110.355 -0.210 110.775 0.210 ;
        RECT 110.965 -0.210 111.385 0.210 ;
        RECT 111.575 -0.210 111.995 0.210 ;
        RECT 113.050 -0.210 113.470 0.210 ;
        RECT 113.660 -0.210 114.080 0.210 ;
        RECT 114.270 -0.210 114.690 0.210 ;
        RECT 114.880 -0.210 115.300 0.210 ;
        RECT 115.490 -0.210 115.910 0.210 ;
        RECT 116.975 -0.210 117.395 0.210 ;
        RECT 117.585 -0.210 118.005 0.210 ;
        RECT 118.195 -0.210 118.615 0.210 ;
        RECT 118.805 -0.210 119.320 0.210 ;
        RECT 125.355 -0.210 125.775 0.210 ;
        RECT 125.965 -0.210 126.385 0.210 ;
        RECT 126.575 -0.210 126.995 0.210 ;
        RECT 127.185 -0.210 127.700 0.210 ;
        RECT 128.500 -0.210 129.015 0.210 ;
        RECT 129.205 -0.210 129.625 0.210 ;
        RECT 129.815 -0.210 130.235 0.210 ;
        RECT 130.425 -0.210 130.845 0.210 ;
        RECT 139.150 -0.210 139.665 0.210 ;
        RECT 139.855 -0.210 140.275 0.210 ;
        RECT 140.465 -0.210 140.885 0.210 ;
        RECT 141.075 -0.210 141.495 0.210 ;
        RECT 142.550 -0.210 142.970 0.210 ;
        RECT 143.160 -0.210 143.580 0.210 ;
        RECT 143.770 -0.210 144.190 0.210 ;
        RECT 144.380 -0.210 144.800 0.210 ;
        RECT 144.990 -0.210 145.410 0.210 ;
        RECT 146.475 -0.210 146.895 0.210 ;
        RECT 147.085 -0.210 147.505 0.210 ;
        RECT 147.695 -0.210 148.115 0.210 ;
        RECT 148.305 -0.210 148.820 0.210 ;
        RECT 154.855 -0.210 155.275 0.210 ;
        RECT 155.465 -0.210 155.885 0.210 ;
        RECT 156.075 -0.210 156.495 0.210 ;
        RECT 156.685 -0.210 157.200 0.210 ;
        RECT 158.000 -0.210 158.515 0.210 ;
        RECT 158.705 -0.210 159.125 0.210 ;
        RECT 159.315 -0.210 159.735 0.210 ;
        RECT 159.925 -0.210 160.345 0.210 ;
        RECT 168.650 -0.210 169.165 0.210 ;
        RECT 169.355 -0.210 169.775 0.210 ;
        RECT 169.965 -0.210 170.385 0.210 ;
        RECT 170.575 -0.210 170.995 0.210 ;
        RECT 172.050 -0.210 172.470 0.210 ;
        RECT 172.660 -0.210 173.080 0.210 ;
        RECT 173.270 -0.210 173.690 0.210 ;
        RECT 173.880 -0.210 174.300 0.210 ;
        RECT 174.490 -0.210 174.910 0.210 ;
        RECT 175.975 -0.210 176.395 0.210 ;
        RECT 176.585 -0.210 177.005 0.210 ;
        RECT 177.195 -0.210 177.615 0.210 ;
        RECT 177.805 -0.210 178.320 0.210 ;
      LAYER met1 ;
        RECT 16.280 37.840 173.490 38.320 ;
        RECT 16.000 35.120 165.390 35.600 ;
        RECT 19.290 31.615 20.420 31.840 ;
        RECT 43.295 31.615 44.035 31.675 ;
        RECT 48.790 31.615 49.920 31.840 ;
        RECT 72.795 31.615 73.535 31.675 ;
        RECT 78.290 31.615 79.420 31.840 ;
        RECT 102.295 31.615 103.035 31.675 ;
        RECT 107.790 31.615 108.920 31.840 ;
        RECT 131.795 31.615 132.535 31.675 ;
        RECT 137.290 31.615 138.420 31.840 ;
        RECT 161.295 31.615 162.035 31.675 ;
        RECT 17.840 30.955 20.420 31.615 ;
        RECT 35.060 31.610 49.920 31.615 ;
        RECT 64.560 31.610 79.420 31.615 ;
        RECT 94.060 31.610 108.920 31.615 ;
        RECT 123.560 31.610 138.420 31.615 ;
        RECT 153.060 31.610 165.440 31.615 ;
        RECT 19.290 30.740 20.420 30.955 ;
        RECT 25.290 30.955 49.920 31.610 ;
        RECT 25.290 30.950 38.550 30.955 ;
        RECT 43.295 30.895 44.035 30.955 ;
        RECT 48.790 30.740 49.920 30.955 ;
        RECT 54.790 30.955 79.420 31.610 ;
        RECT 54.790 30.950 68.050 30.955 ;
        RECT 72.795 30.895 73.535 30.955 ;
        RECT 78.290 30.740 79.420 30.955 ;
        RECT 84.290 30.955 108.920 31.610 ;
        RECT 84.290 30.950 97.550 30.955 ;
        RECT 102.295 30.895 103.035 30.955 ;
        RECT 107.790 30.740 108.920 30.955 ;
        RECT 113.790 30.955 138.420 31.610 ;
        RECT 113.790 30.950 127.050 30.955 ;
        RECT 131.795 30.895 132.535 30.955 ;
        RECT 137.290 30.740 138.420 30.955 ;
        RECT 143.290 30.955 165.440 31.610 ;
        RECT 143.290 30.950 156.550 30.955 ;
        RECT 161.295 30.895 162.035 30.955 ;
        RECT 3.820 29.680 20.290 30.160 ;
        RECT 30.790 28.920 34.090 28.950 ;
        RECT 60.290 28.920 63.590 28.950 ;
        RECT 89.790 28.920 93.090 28.950 ;
        RECT 119.290 28.920 122.590 28.950 ;
        RECT 148.790 28.920 152.090 28.950 ;
        RECT 30.790 28.860 34.890 28.920 ;
        RECT 6.800 28.710 7.220 28.740 ;
        RECT 17.000 28.710 34.890 28.860 ;
        RECT 6.800 28.410 34.890 28.710 ;
        RECT 6.800 28.380 7.220 28.410 ;
        RECT 17.000 28.260 34.890 28.410 ;
        RECT 30.790 28.200 34.890 28.260 ;
        RECT 41.425 28.860 41.985 28.920 ;
        RECT 60.290 28.860 64.390 28.920 ;
        RECT 41.425 28.260 64.390 28.860 ;
        RECT 41.425 28.200 41.985 28.260 ;
        RECT 60.290 28.200 64.390 28.260 ;
        RECT 70.925 28.860 71.485 28.920 ;
        RECT 89.790 28.860 93.890 28.920 ;
        RECT 70.925 28.260 93.890 28.860 ;
        RECT 70.925 28.200 71.485 28.260 ;
        RECT 89.790 28.200 93.890 28.260 ;
        RECT 100.425 28.860 100.985 28.920 ;
        RECT 119.290 28.860 123.390 28.920 ;
        RECT 100.425 28.260 123.390 28.860 ;
        RECT 100.425 28.200 100.985 28.260 ;
        RECT 119.290 28.200 123.390 28.260 ;
        RECT 129.925 28.860 130.485 28.920 ;
        RECT 148.790 28.860 152.890 28.920 ;
        RECT 129.925 28.260 152.890 28.860 ;
        RECT 129.925 28.200 130.485 28.260 ;
        RECT 148.790 28.200 152.890 28.260 ;
        RECT 159.425 28.860 159.985 28.920 ;
        RECT 159.425 28.260 165.440 28.860 ;
        RECT 159.425 28.200 159.985 28.260 ;
        RECT 0.500 26.960 9.965 27.440 ;
        RECT 15.005 24.240 172.440 24.720 ;
        RECT 17.890 21.990 165.390 22.000 ;
        RECT 17.000 21.510 177.530 21.990 ;
        RECT 2.000 16.080 180.440 16.560 ;
        RECT 0.500 13.360 179.440 13.840 ;
        RECT 7.405 9.820 7.965 9.880 ;
        RECT 2.000 9.220 7.965 9.820 ;
        RECT 7.405 9.160 7.965 9.220 ;
        RECT 14.500 9.820 18.600 9.880 ;
        RECT 36.905 9.820 37.465 9.880 ;
        RECT 14.500 9.220 37.465 9.820 ;
        RECT 14.500 9.160 18.600 9.220 ;
        RECT 36.905 9.160 37.465 9.220 ;
        RECT 44.000 9.820 48.100 9.880 ;
        RECT 66.405 9.820 66.965 9.880 ;
        RECT 44.000 9.220 66.965 9.820 ;
        RECT 44.000 9.160 48.100 9.220 ;
        RECT 66.405 9.160 66.965 9.220 ;
        RECT 73.500 9.820 77.600 9.880 ;
        RECT 95.905 9.820 96.465 9.880 ;
        RECT 73.500 9.220 96.465 9.820 ;
        RECT 73.500 9.160 77.600 9.220 ;
        RECT 95.905 9.160 96.465 9.220 ;
        RECT 103.000 9.820 107.100 9.880 ;
        RECT 125.405 9.820 125.965 9.880 ;
        RECT 103.000 9.220 125.965 9.820 ;
        RECT 103.000 9.160 107.100 9.220 ;
        RECT 125.405 9.160 125.965 9.220 ;
        RECT 132.500 9.820 136.600 9.880 ;
        RECT 154.905 9.820 155.465 9.880 ;
        RECT 132.500 9.220 155.465 9.820 ;
        RECT 132.500 9.160 136.600 9.220 ;
        RECT 154.905 9.160 155.465 9.220 ;
        RECT 162.000 9.820 166.100 9.880 ;
        RECT 162.000 9.220 179.000 9.820 ;
        RECT 162.000 9.160 166.100 9.220 ;
        RECT 15.300 9.130 18.600 9.160 ;
        RECT 44.800 9.130 48.100 9.160 ;
        RECT 74.300 9.130 77.600 9.160 ;
        RECT 103.800 9.130 107.100 9.160 ;
        RECT 133.300 9.130 136.600 9.160 ;
        RECT 162.800 9.130 166.100 9.160 ;
        RECT 5.355 7.125 6.095 7.185 ;
        RECT 10.840 7.125 24.100 7.130 ;
        RECT 2.000 6.470 24.100 7.125 ;
        RECT 28.970 7.125 30.100 7.340 ;
        RECT 34.855 7.125 35.595 7.185 ;
        RECT 40.340 7.125 53.600 7.130 ;
        RECT 28.970 6.470 53.600 7.125 ;
        RECT 58.470 7.125 59.600 7.340 ;
        RECT 64.355 7.125 65.095 7.185 ;
        RECT 69.840 7.125 83.100 7.130 ;
        RECT 58.470 6.470 83.100 7.125 ;
        RECT 87.970 7.125 89.100 7.340 ;
        RECT 93.855 7.125 94.595 7.185 ;
        RECT 99.340 7.125 112.600 7.130 ;
        RECT 87.970 6.470 112.600 7.125 ;
        RECT 117.470 7.125 118.600 7.340 ;
        RECT 123.355 7.125 124.095 7.185 ;
        RECT 128.840 7.125 142.100 7.130 ;
        RECT 117.470 6.470 142.100 7.125 ;
        RECT 146.970 7.125 148.100 7.340 ;
        RECT 152.855 7.125 153.595 7.185 ;
        RECT 158.340 7.125 171.600 7.130 ;
        RECT 146.970 6.470 171.600 7.125 ;
        RECT 176.470 7.125 177.600 7.340 ;
        RECT 176.470 7.095 179.000 7.125 ;
        RECT 172.640 6.495 179.000 7.095 ;
        RECT 2.000 6.465 14.330 6.470 ;
        RECT 28.970 6.465 43.830 6.470 ;
        RECT 58.470 6.465 73.330 6.470 ;
        RECT 87.970 6.465 102.830 6.470 ;
        RECT 117.470 6.465 132.330 6.470 ;
        RECT 146.970 6.465 161.830 6.470 ;
        RECT 176.470 6.465 179.000 6.495 ;
        RECT 5.355 6.405 6.095 6.465 ;
        RECT 28.970 6.240 30.100 6.465 ;
        RECT 34.855 6.405 35.595 6.465 ;
        RECT 58.470 6.240 59.600 6.465 ;
        RECT 64.355 6.405 65.095 6.465 ;
        RECT 87.970 6.240 89.100 6.465 ;
        RECT 93.855 6.405 94.595 6.465 ;
        RECT 117.470 6.240 118.600 6.465 ;
        RECT 123.355 6.405 124.095 6.465 ;
        RECT 146.970 6.240 148.100 6.465 ;
        RECT 152.855 6.405 153.595 6.465 ;
        RECT 176.470 6.240 177.600 6.465 ;
        RECT 0.500 2.480 179.440 2.960 ;
        RECT 2.000 -0.240 180.440 0.240 ;
      LAYER via ;
        RECT 39.000 37.940 39.260 38.200 ;
        RECT 39.370 37.940 39.630 38.200 ;
        RECT 39.740 37.940 40.000 38.200 ;
        RECT 70.000 37.940 70.260 38.200 ;
        RECT 70.370 37.940 70.630 38.200 ;
        RECT 70.740 37.940 71.000 38.200 ;
        RECT 112.000 37.940 112.260 38.200 ;
        RECT 112.370 37.940 112.630 38.200 ;
        RECT 112.740 37.940 113.000 38.200 ;
        RECT 143.000 37.940 143.260 38.200 ;
        RECT 143.370 37.940 143.630 38.200 ;
        RECT 143.740 37.940 144.000 38.200 ;
        RECT 172.490 37.950 172.750 38.210 ;
        RECT 172.810 37.950 173.070 38.210 ;
        RECT 173.130 37.950 173.390 38.210 ;
        RECT 18.045 30.995 18.625 31.575 ;
        RECT 164.480 30.995 165.380 31.575 ;
        RECT 17.925 28.270 18.825 28.850 ;
        RECT 164.470 28.270 165.370 28.850 ;
        RECT 39.000 21.620 39.260 21.880 ;
        RECT 39.370 21.620 39.630 21.880 ;
        RECT 39.740 21.620 40.000 21.880 ;
        RECT 70.000 21.620 70.260 21.880 ;
        RECT 70.370 21.620 70.630 21.880 ;
        RECT 70.740 21.620 71.000 21.880 ;
        RECT 112.000 21.620 112.260 21.880 ;
        RECT 112.370 21.620 112.630 21.880 ;
        RECT 112.740 21.620 113.000 21.880 ;
        RECT 143.000 21.620 143.260 21.880 ;
        RECT 143.370 21.620 143.630 21.880 ;
        RECT 143.740 21.620 144.000 21.880 ;
        RECT 173.155 21.650 173.415 21.910 ;
        RECT 173.530 21.650 173.790 21.910 ;
        RECT 173.910 21.650 174.170 21.910 ;
        RECT 174.285 21.650 174.545 21.910 ;
        RECT 174.660 21.650 174.920 21.910 ;
        RECT 175.035 21.650 175.295 21.910 ;
        RECT 175.415 21.650 175.675 21.910 ;
        RECT 175.790 21.650 176.050 21.910 ;
        RECT 176.165 21.650 176.425 21.910 ;
        RECT 176.535 21.650 176.795 21.910 ;
        RECT 176.915 21.650 177.175 21.910 ;
        RECT 39.000 16.180 39.260 16.440 ;
        RECT 39.370 16.180 39.630 16.440 ;
        RECT 39.740 16.180 40.000 16.440 ;
        RECT 70.000 16.180 70.260 16.440 ;
        RECT 70.370 16.180 70.630 16.440 ;
        RECT 70.740 16.180 71.000 16.440 ;
        RECT 112.000 16.180 112.260 16.440 ;
        RECT 112.370 16.180 112.630 16.440 ;
        RECT 112.740 16.180 113.000 16.440 ;
        RECT 143.000 16.180 143.260 16.440 ;
        RECT 143.370 16.180 143.630 16.440 ;
        RECT 143.740 16.180 144.000 16.440 ;
        RECT 179.465 16.190 179.725 16.450 ;
        RECT 179.785 16.190 180.045 16.450 ;
        RECT 180.105 16.190 180.365 16.450 ;
        RECT 6.765 9.230 7.345 9.810 ;
        RECT 166.150 9.230 166.730 9.810 ;
        RECT 166.870 9.230 167.450 9.810 ;
        RECT 4.055 6.505 4.635 7.085 ;
        RECT 172.760 6.505 173.340 7.085 ;
        RECT 39.000 -0.140 39.260 0.120 ;
        RECT 39.370 -0.140 39.630 0.120 ;
        RECT 39.740 -0.140 40.000 0.120 ;
        RECT 70.000 -0.140 70.260 0.120 ;
        RECT 70.370 -0.140 70.630 0.120 ;
        RECT 70.740 -0.140 71.000 0.120 ;
        RECT 112.000 -0.140 112.260 0.120 ;
        RECT 112.370 -0.140 112.630 0.120 ;
        RECT 112.740 -0.140 113.000 0.120 ;
        RECT 143.000 -0.140 143.260 0.120 ;
        RECT 143.370 -0.140 143.630 0.120 ;
        RECT 143.740 -0.140 144.000 0.120 ;
        RECT 179.475 -0.130 179.735 0.130 ;
        RECT 179.795 -0.130 180.055 0.130 ;
        RECT 180.115 -0.130 180.375 0.130 ;
      LAYER met2 ;
        RECT 39.000 37.870 40.000 38.270 ;
        RECT 70.000 37.870 71.000 38.270 ;
        RECT 112.000 37.870 113.000 38.270 ;
        RECT 143.000 37.870 144.000 38.270 ;
        RECT 17.890 31.635 18.785 31.665 ;
        RECT 14.420 30.935 18.785 31.635 ;
        RECT 14.420 20.050 15.120 30.935 ;
        RECT 17.890 30.905 18.785 30.935 ;
        RECT 164.470 31.635 165.390 31.665 ;
        RECT 164.470 30.935 169.490 31.635 ;
        RECT 164.470 30.905 165.390 30.935 ;
        RECT 4.000 19.350 15.120 20.050 ;
        RECT 17.120 28.210 18.865 28.910 ;
        RECT 164.450 28.210 166.790 28.910 ;
        RECT 4.000 18.535 4.700 19.350 ;
        RECT 3.995 12.965 4.700 18.535 ;
        RECT 17.120 17.350 17.820 28.210 ;
        RECT 39.000 21.550 40.000 21.950 ;
        RECT 70.000 21.550 71.000 21.950 ;
        RECT 112.000 21.550 113.000 21.950 ;
        RECT 143.000 21.550 144.000 21.950 ;
        RECT 6.705 16.650 17.820 17.350 ;
        RECT 3.995 6.415 4.695 12.965 ;
        RECT 6.705 9.170 7.405 16.650 ;
        RECT 13.270 16.630 14.070 16.650 ;
        RECT 39.000 16.110 40.000 16.510 ;
        RECT 70.000 16.110 71.000 16.510 ;
        RECT 112.000 16.110 113.000 16.510 ;
        RECT 143.000 16.110 144.000 16.510 ;
        RECT 166.090 9.870 166.790 28.210 ;
        RECT 168.790 17.635 169.490 30.935 ;
        RECT 172.440 22.240 173.440 38.370 ;
        RECT 172.440 21.440 183.500 22.240 ;
        RECT 172.440 21.240 180.440 21.440 ;
        RECT 179.440 20.700 180.435 21.240 ;
        RECT 168.790 16.935 173.400 17.635 ;
        RECT 166.090 9.140 167.460 9.870 ;
        RECT 172.700 6.445 173.400 16.935 ;
        RECT 39.000 -0.210 40.000 0.190 ;
        RECT 70.000 -0.210 71.000 0.190 ;
        RECT 112.000 -0.210 113.000 0.190 ;
        RECT 143.000 -0.210 144.000 0.190 ;
        RECT 179.440 -0.290 180.440 20.700 ;
      LAYER via2 ;
        RECT 39.100 37.920 39.400 38.220 ;
        RECT 39.600 37.920 39.900 38.220 ;
        RECT 70.100 37.920 70.400 38.220 ;
        RECT 70.600 37.920 70.900 38.220 ;
        RECT 112.100 37.920 112.400 38.220 ;
        RECT 112.600 37.920 112.900 38.220 ;
        RECT 143.100 37.920 143.400 38.220 ;
        RECT 143.600 37.920 143.900 38.220 ;
        RECT 39.100 21.600 39.400 21.900 ;
        RECT 39.600 21.600 39.900 21.900 ;
        RECT 70.100 21.600 70.400 21.900 ;
        RECT 70.600 21.600 70.900 21.900 ;
        RECT 112.100 21.600 112.400 21.900 ;
        RECT 112.600 21.600 112.900 21.900 ;
        RECT 143.100 21.600 143.400 21.900 ;
        RECT 143.600 21.600 143.900 21.900 ;
        RECT 39.100 16.160 39.400 16.460 ;
        RECT 39.600 16.160 39.900 16.460 ;
        RECT 70.100 16.160 70.400 16.460 ;
        RECT 70.600 16.160 70.900 16.460 ;
        RECT 112.100 16.160 112.400 16.460 ;
        RECT 112.600 16.160 112.900 16.460 ;
        RECT 143.100 16.160 143.400 16.460 ;
        RECT 143.600 16.160 143.900 16.460 ;
        RECT 179.750 19.100 180.150 19.500 ;
        RECT 179.750 18.570 180.150 18.970 ;
        RECT 39.100 -0.160 39.400 0.140 ;
        RECT 39.600 -0.160 39.900 0.140 ;
        RECT 70.100 -0.160 70.400 0.140 ;
        RECT 70.600 -0.160 70.900 0.140 ;
        RECT 112.100 -0.160 112.400 0.140 ;
        RECT 112.600 -0.160 112.900 0.140 ;
        RECT 143.100 -0.160 143.400 0.140 ;
        RECT 143.600 -0.160 143.900 0.140 ;
      LAYER met3 ;
        RECT 39.000 19.610 40.000 38.320 ;
        RECT 70.000 19.610 71.000 38.320 ;
        RECT 112.000 19.610 113.000 38.320 ;
        RECT 143.000 19.610 144.000 38.320 ;
        RECT 39.000 18.460 180.440 19.610 ;
        RECT 39.000 -0.240 40.000 18.460 ;
        RECT 70.000 -0.240 71.000 18.460 ;
        RECT 112.000 -0.240 113.000 18.460 ;
        RECT 143.000 -0.240 144.000 18.460 ;
  END
END ring_osc
MACRO power_ring_2_2
  CLASS BLOCK ;
  FOREIGN power_ring_2_2 ;
  ORIGIN -135.000 -16.000 ;
  SIZE 182.000 BY 105.000 ;
  OBS
      LAYER met3 ;
        RECT 140.000 119.000 312.000 121.000 ;
        RECT 135.000 115.000 317.000 117.000 ;
        RECT 135.000 20.000 317.000 22.000 ;
        RECT 140.000 16.000 312.000 18.000 ;
      LAYER via3 ;
        RECT 140.200 120.400 140.600 120.800 ;
        RECT 140.800 120.400 141.200 120.800 ;
        RECT 141.400 120.400 141.800 120.800 ;
        RECT 153.200 120.400 153.600 120.800 ;
        RECT 153.800 120.400 154.200 120.800 ;
        RECT 154.400 120.400 154.800 120.800 ;
        RECT 189.200 120.400 189.600 120.800 ;
        RECT 189.800 120.400 190.200 120.800 ;
        RECT 190.400 120.400 190.800 120.800 ;
        RECT 225.200 120.400 225.600 120.800 ;
        RECT 225.800 120.400 226.200 120.800 ;
        RECT 226.400 120.400 226.800 120.800 ;
        RECT 261.200 120.400 261.600 120.800 ;
        RECT 261.800 120.400 262.200 120.800 ;
        RECT 262.400 120.400 262.800 120.800 ;
        RECT 297.200 120.400 297.600 120.800 ;
        RECT 297.800 120.400 298.200 120.800 ;
        RECT 298.400 120.400 298.800 120.800 ;
        RECT 310.200 120.400 310.600 120.800 ;
        RECT 310.800 120.400 311.200 120.800 ;
        RECT 311.400 120.400 311.800 120.800 ;
        RECT 140.200 119.800 140.600 120.200 ;
        RECT 140.800 119.800 141.200 120.200 ;
        RECT 141.400 119.800 141.800 120.200 ;
        RECT 153.200 119.800 153.600 120.200 ;
        RECT 153.800 119.800 154.200 120.200 ;
        RECT 154.400 119.800 154.800 120.200 ;
        RECT 189.200 119.800 189.600 120.200 ;
        RECT 189.800 119.800 190.200 120.200 ;
        RECT 190.400 119.800 190.800 120.200 ;
        RECT 225.200 119.800 225.600 120.200 ;
        RECT 225.800 119.800 226.200 120.200 ;
        RECT 226.400 119.800 226.800 120.200 ;
        RECT 261.200 119.800 261.600 120.200 ;
        RECT 261.800 119.800 262.200 120.200 ;
        RECT 262.400 119.800 262.800 120.200 ;
        RECT 297.200 119.800 297.600 120.200 ;
        RECT 297.800 119.800 298.200 120.200 ;
        RECT 298.400 119.800 298.800 120.200 ;
        RECT 310.200 119.800 310.600 120.200 ;
        RECT 310.800 119.800 311.200 120.200 ;
        RECT 311.400 119.800 311.800 120.200 ;
        RECT 140.200 119.200 140.600 119.600 ;
        RECT 140.800 119.200 141.200 119.600 ;
        RECT 141.400 119.200 141.800 119.600 ;
        RECT 153.200 119.200 153.600 119.600 ;
        RECT 153.800 119.200 154.200 119.600 ;
        RECT 154.400 119.200 154.800 119.600 ;
        RECT 189.200 119.200 189.600 119.600 ;
        RECT 189.800 119.200 190.200 119.600 ;
        RECT 190.400 119.200 190.800 119.600 ;
        RECT 225.200 119.200 225.600 119.600 ;
        RECT 225.800 119.200 226.200 119.600 ;
        RECT 226.400 119.200 226.800 119.600 ;
        RECT 261.200 119.200 261.600 119.600 ;
        RECT 261.800 119.200 262.200 119.600 ;
        RECT 262.400 119.200 262.800 119.600 ;
        RECT 297.200 119.200 297.600 119.600 ;
        RECT 297.800 119.200 298.200 119.600 ;
        RECT 298.400 119.200 298.800 119.600 ;
        RECT 310.200 119.200 310.600 119.600 ;
        RECT 310.800 119.200 311.200 119.600 ;
        RECT 311.400 119.200 311.800 119.600 ;
        RECT 135.200 116.400 135.600 116.800 ;
        RECT 135.800 116.400 136.200 116.800 ;
        RECT 136.400 116.400 136.800 116.800 ;
        RECT 171.200 116.400 171.600 116.800 ;
        RECT 171.800 116.400 172.200 116.800 ;
        RECT 172.400 116.400 172.800 116.800 ;
        RECT 207.200 116.400 207.600 116.800 ;
        RECT 207.800 116.400 208.200 116.800 ;
        RECT 208.400 116.400 208.800 116.800 ;
        RECT 243.200 116.400 243.600 116.800 ;
        RECT 243.800 116.400 244.200 116.800 ;
        RECT 244.400 116.400 244.800 116.800 ;
        RECT 279.200 116.400 279.600 116.800 ;
        RECT 279.800 116.400 280.200 116.800 ;
        RECT 280.400 116.400 280.800 116.800 ;
        RECT 315.200 116.400 315.600 116.800 ;
        RECT 315.800 116.400 316.200 116.800 ;
        RECT 316.400 116.400 316.800 116.800 ;
        RECT 135.200 115.800 135.600 116.200 ;
        RECT 135.800 115.800 136.200 116.200 ;
        RECT 136.400 115.800 136.800 116.200 ;
        RECT 171.200 115.800 171.600 116.200 ;
        RECT 171.800 115.800 172.200 116.200 ;
        RECT 172.400 115.800 172.800 116.200 ;
        RECT 207.200 115.800 207.600 116.200 ;
        RECT 207.800 115.800 208.200 116.200 ;
        RECT 208.400 115.800 208.800 116.200 ;
        RECT 243.200 115.800 243.600 116.200 ;
        RECT 243.800 115.800 244.200 116.200 ;
        RECT 244.400 115.800 244.800 116.200 ;
        RECT 279.200 115.800 279.600 116.200 ;
        RECT 279.800 115.800 280.200 116.200 ;
        RECT 280.400 115.800 280.800 116.200 ;
        RECT 315.200 115.800 315.600 116.200 ;
        RECT 315.800 115.800 316.200 116.200 ;
        RECT 316.400 115.800 316.800 116.200 ;
        RECT 135.200 115.200 135.600 115.600 ;
        RECT 135.800 115.200 136.200 115.600 ;
        RECT 136.400 115.200 136.800 115.600 ;
        RECT 171.200 115.200 171.600 115.600 ;
        RECT 171.800 115.200 172.200 115.600 ;
        RECT 172.400 115.200 172.800 115.600 ;
        RECT 207.200 115.200 207.600 115.600 ;
        RECT 207.800 115.200 208.200 115.600 ;
        RECT 208.400 115.200 208.800 115.600 ;
        RECT 243.200 115.200 243.600 115.600 ;
        RECT 243.800 115.200 244.200 115.600 ;
        RECT 244.400 115.200 244.800 115.600 ;
        RECT 279.200 115.200 279.600 115.600 ;
        RECT 279.800 115.200 280.200 115.600 ;
        RECT 280.400 115.200 280.800 115.600 ;
        RECT 315.200 115.200 315.600 115.600 ;
        RECT 315.800 115.200 316.200 115.600 ;
        RECT 316.400 115.200 316.800 115.600 ;
        RECT 135.200 21.400 135.600 21.800 ;
        RECT 135.800 21.400 136.200 21.800 ;
        RECT 136.400 21.400 136.800 21.800 ;
        RECT 171.200 21.400 171.600 21.800 ;
        RECT 171.800 21.400 172.200 21.800 ;
        RECT 172.400 21.400 172.800 21.800 ;
        RECT 207.200 21.400 207.600 21.800 ;
        RECT 207.800 21.400 208.200 21.800 ;
        RECT 208.400 21.400 208.800 21.800 ;
        RECT 243.200 21.400 243.600 21.800 ;
        RECT 243.800 21.400 244.200 21.800 ;
        RECT 244.400 21.400 244.800 21.800 ;
        RECT 279.200 21.400 279.600 21.800 ;
        RECT 279.800 21.400 280.200 21.800 ;
        RECT 280.400 21.400 280.800 21.800 ;
        RECT 315.200 21.400 315.600 21.800 ;
        RECT 315.800 21.400 316.200 21.800 ;
        RECT 316.400 21.400 316.800 21.800 ;
        RECT 135.200 20.800 135.600 21.200 ;
        RECT 135.800 20.800 136.200 21.200 ;
        RECT 136.400 20.800 136.800 21.200 ;
        RECT 171.200 20.800 171.600 21.200 ;
        RECT 171.800 20.800 172.200 21.200 ;
        RECT 172.400 20.800 172.800 21.200 ;
        RECT 207.200 20.800 207.600 21.200 ;
        RECT 207.800 20.800 208.200 21.200 ;
        RECT 208.400 20.800 208.800 21.200 ;
        RECT 243.200 20.800 243.600 21.200 ;
        RECT 243.800 20.800 244.200 21.200 ;
        RECT 244.400 20.800 244.800 21.200 ;
        RECT 279.200 20.800 279.600 21.200 ;
        RECT 279.800 20.800 280.200 21.200 ;
        RECT 280.400 20.800 280.800 21.200 ;
        RECT 315.200 20.800 315.600 21.200 ;
        RECT 315.800 20.800 316.200 21.200 ;
        RECT 316.400 20.800 316.800 21.200 ;
        RECT 135.200 20.200 135.600 20.600 ;
        RECT 135.800 20.200 136.200 20.600 ;
        RECT 136.400 20.200 136.800 20.600 ;
        RECT 171.200 20.200 171.600 20.600 ;
        RECT 171.800 20.200 172.200 20.600 ;
        RECT 172.400 20.200 172.800 20.600 ;
        RECT 207.200 20.200 207.600 20.600 ;
        RECT 207.800 20.200 208.200 20.600 ;
        RECT 208.400 20.200 208.800 20.600 ;
        RECT 243.200 20.200 243.600 20.600 ;
        RECT 243.800 20.200 244.200 20.600 ;
        RECT 244.400 20.200 244.800 20.600 ;
        RECT 279.200 20.200 279.600 20.600 ;
        RECT 279.800 20.200 280.200 20.600 ;
        RECT 280.400 20.200 280.800 20.600 ;
        RECT 315.200 20.200 315.600 20.600 ;
        RECT 315.800 20.200 316.200 20.600 ;
        RECT 316.400 20.200 316.800 20.600 ;
        RECT 140.200 17.400 140.600 17.800 ;
        RECT 140.800 17.400 141.200 17.800 ;
        RECT 141.400 17.400 141.800 17.800 ;
        RECT 153.200 17.400 153.600 17.800 ;
        RECT 153.800 17.400 154.200 17.800 ;
        RECT 154.400 17.400 154.800 17.800 ;
        RECT 189.200 17.400 189.600 17.800 ;
        RECT 189.800 17.400 190.200 17.800 ;
        RECT 190.400 17.400 190.800 17.800 ;
        RECT 225.200 17.400 225.600 17.800 ;
        RECT 225.800 17.400 226.200 17.800 ;
        RECT 226.400 17.400 226.800 17.800 ;
        RECT 261.200 17.400 261.600 17.800 ;
        RECT 261.800 17.400 262.200 17.800 ;
        RECT 262.400 17.400 262.800 17.800 ;
        RECT 297.200 17.400 297.600 17.800 ;
        RECT 297.800 17.400 298.200 17.800 ;
        RECT 298.400 17.400 298.800 17.800 ;
        RECT 310.200 17.400 310.600 17.800 ;
        RECT 310.800 17.400 311.200 17.800 ;
        RECT 311.400 17.400 311.800 17.800 ;
        RECT 140.200 16.800 140.600 17.200 ;
        RECT 140.800 16.800 141.200 17.200 ;
        RECT 141.400 16.800 141.800 17.200 ;
        RECT 153.200 16.800 153.600 17.200 ;
        RECT 153.800 16.800 154.200 17.200 ;
        RECT 154.400 16.800 154.800 17.200 ;
        RECT 189.200 16.800 189.600 17.200 ;
        RECT 189.800 16.800 190.200 17.200 ;
        RECT 190.400 16.800 190.800 17.200 ;
        RECT 225.200 16.800 225.600 17.200 ;
        RECT 225.800 16.800 226.200 17.200 ;
        RECT 226.400 16.800 226.800 17.200 ;
        RECT 261.200 16.800 261.600 17.200 ;
        RECT 261.800 16.800 262.200 17.200 ;
        RECT 262.400 16.800 262.800 17.200 ;
        RECT 297.200 16.800 297.600 17.200 ;
        RECT 297.800 16.800 298.200 17.200 ;
        RECT 298.400 16.800 298.800 17.200 ;
        RECT 310.200 16.800 310.600 17.200 ;
        RECT 310.800 16.800 311.200 17.200 ;
        RECT 311.400 16.800 311.800 17.200 ;
        RECT 140.200 16.200 140.600 16.600 ;
        RECT 140.800 16.200 141.200 16.600 ;
        RECT 141.400 16.200 141.800 16.600 ;
        RECT 153.200 16.200 153.600 16.600 ;
        RECT 153.800 16.200 154.200 16.600 ;
        RECT 154.400 16.200 154.800 16.600 ;
        RECT 189.200 16.200 189.600 16.600 ;
        RECT 189.800 16.200 190.200 16.600 ;
        RECT 190.400 16.200 190.800 16.600 ;
        RECT 225.200 16.200 225.600 16.600 ;
        RECT 225.800 16.200 226.200 16.600 ;
        RECT 226.400 16.200 226.800 16.600 ;
        RECT 261.200 16.200 261.600 16.600 ;
        RECT 261.800 16.200 262.200 16.600 ;
        RECT 262.400 16.200 262.800 16.600 ;
        RECT 297.200 16.200 297.600 16.600 ;
        RECT 297.800 16.200 298.200 16.600 ;
        RECT 298.400 16.200 298.800 16.600 ;
        RECT 310.200 16.200 310.600 16.600 ;
        RECT 310.800 16.200 311.200 16.600 ;
        RECT 311.400 16.200 311.800 16.600 ;
      LAYER met4 ;
        RECT 135.000 20.000 137.000 117.000 ;
        RECT 140.000 16.000 142.000 121.000 ;
        RECT 153.000 16.000 155.000 121.000 ;
        RECT 171.000 20.000 173.000 117.000 ;
        RECT 189.000 16.000 191.000 121.000 ;
        RECT 207.000 20.000 209.000 117.000 ;
        RECT 225.000 16.000 227.000 121.000 ;
        RECT 243.000 20.000 245.000 117.000 ;
        RECT 261.000 16.000 263.000 121.000 ;
        RECT 279.000 20.000 281.000 117.000 ;
        RECT 297.000 16.000 299.000 121.000 ;
        RECT 310.000 16.000 312.000 121.000 ;
        RECT 315.000 20.000 317.000 117.000 ;
  END
END power_ring_2_2
MACRO pwell_co_ring
  CLASS BLOCK ;
  FOREIGN pwell_co_ring ;
  ORIGIN -0.880 -30.000 ;
  SIZE 179.740 BY 42.500 ;
  OBS
      LAYER li1 ;
        RECT 15.920 72.000 166.580 72.500 ;
        RECT 16.000 52.500 16.500 72.000 ;
        RECT 166.000 52.500 166.500 72.000 ;
        RECT 15.920 52.000 166.580 52.500 ;
        RECT 0.920 50.000 180.580 50.500 ;
        RECT 1.000 30.500 1.500 50.000 ;
        RECT 180.000 30.500 180.500 50.000 ;
        RECT 0.920 30.000 180.580 30.500 ;
  END
END pwell_co_ring
MACRO vco
  CLASS BLOCK ;
  FOREIGN vco ;
  ORIGIN 0.000 0.000 ;
  SIZE 183.010 BY 105.000 ;
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.680500 ;
    PORT
      LAYER met2 ;
        RECT 16.630 61.510 18.375 62.210 ;
        RECT 16.630 50.650 17.330 61.510 ;
        RECT 6.215 49.950 17.330 50.650 ;
        RECT 6.215 43.010 6.915 49.950 ;
        RECT 12.780 49.930 13.580 49.950 ;
        RECT 6.140 42.550 7.060 43.010 ;
        RECT 6.215 42.470 6.915 42.550 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 31.050 42.550 31.970 43.010 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 46.690 61.640 47.610 62.100 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 60.490 42.550 61.410 43.010 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 75.670 61.620 76.590 62.080 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 89.930 42.550 90.850 43.010 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 105.110 61.630 106.030 62.090 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 119.830 42.550 120.750 43.010 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 135.010 61.620 135.930 62.080 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 149.270 42.550 150.190 43.010 ;
    END
  END p[9]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 163.960 61.510 166.300 62.210 ;
        RECT 165.600 43.170 166.300 61.510 ;
        RECT 165.600 42.440 166.970 43.170 ;
    END
  END p[10]
  PIN input_analog
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 137.169998 ;
    PORT
      LAYER met3 ;
        RECT 38.510 52.910 39.510 71.620 ;
        RECT 69.510 52.910 70.510 71.620 ;
        RECT 111.510 52.910 112.510 71.620 ;
        RECT 142.510 52.910 143.510 71.620 ;
        RECT 181.980 54.740 183.010 55.540 ;
        RECT 38.510 51.760 179.950 52.910 ;
        RECT 38.510 33.060 39.510 51.760 ;
        RECT 69.510 33.060 70.510 51.760 ;
        RECT 111.510 33.060 112.510 51.760 ;
        RECT 142.510 33.060 143.510 51.760 ;
    END
  END input_analog
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 3.140 61.805 5.820 63.640 ;
        RECT 7.310 61.805 9.070 63.640 ;
        RECT 17.900 57.545 23.750 63.420 ;
        RECT 28.730 63.080 34.580 68.935 ;
        RECT 42.350 63.610 46.110 68.885 ;
        RECT 35.875 57.550 39.635 62.860 ;
        RECT 47.400 57.545 53.250 63.420 ;
        RECT 58.230 63.080 64.080 68.935 ;
        RECT 71.850 63.610 75.610 68.885 ;
        RECT 65.375 57.550 69.135 62.860 ;
        RECT 76.900 57.545 82.750 63.420 ;
        RECT 87.730 63.080 93.580 68.935 ;
        RECT 101.350 63.610 105.110 68.885 ;
        RECT 94.875 57.550 98.635 62.860 ;
        RECT 106.400 57.545 112.250 63.420 ;
        RECT 117.230 63.080 123.080 68.935 ;
        RECT 130.850 63.610 134.610 68.885 ;
        RECT 124.375 57.550 128.135 62.860 ;
        RECT 135.900 57.545 141.750 63.420 ;
        RECT 146.730 63.080 152.580 68.935 ;
        RECT 160.350 63.610 164.110 68.885 ;
        RECT 153.875 57.550 157.635 62.860 ;
        RECT 8.775 41.820 12.535 47.130 ;
        RECT 2.300 35.795 6.060 41.070 ;
        RECT 13.830 35.745 19.680 41.600 ;
        RECT 24.660 41.260 30.510 47.135 ;
        RECT 38.275 41.820 42.035 47.130 ;
        RECT 31.800 35.795 35.560 41.070 ;
        RECT 43.330 35.745 49.180 41.600 ;
        RECT 54.160 41.260 60.010 47.135 ;
        RECT 67.775 41.820 71.535 47.130 ;
        RECT 61.300 35.795 65.060 41.070 ;
        RECT 72.830 35.745 78.680 41.600 ;
        RECT 83.660 41.260 89.510 47.135 ;
        RECT 97.275 41.820 101.035 47.130 ;
        RECT 90.800 35.795 94.560 41.070 ;
        RECT 102.330 35.745 108.180 41.600 ;
        RECT 113.160 41.260 119.010 47.135 ;
        RECT 126.775 41.820 130.535 47.130 ;
        RECT 120.300 35.795 124.060 41.070 ;
        RECT 131.830 35.745 137.680 41.600 ;
        RECT 142.660 41.260 148.510 47.135 ;
        RECT 156.275 41.820 160.035 47.130 ;
        RECT 149.800 35.795 153.560 41.070 ;
        RECT 161.330 35.745 167.180 41.600 ;
        RECT 172.160 41.260 178.010 47.135 ;
      LAYER met4 ;
        RECT 5.000 0.000 7.000 105.000 ;
        RECT 18.000 0.000 20.000 105.000 ;
        RECT 54.000 0.000 56.000 105.000 ;
        RECT 90.000 0.000 92.000 105.000 ;
        RECT 126.000 0.000 128.000 105.000 ;
        RECT 162.000 0.000 164.000 105.000 ;
        RECT 175.000 0.000 177.000 105.000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 0.000 4.000 2.000 101.000 ;
        RECT 36.000 4.000 38.000 101.000 ;
        RECT 72.000 4.000 74.000 101.000 ;
        RECT 108.000 4.000 110.000 101.000 ;
        RECT 144.000 4.000 146.000 101.000 ;
        RECT 180.000 4.000 182.000 101.000 ;
    END
  END vssd2
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER met3 ;
        RECT 2.370 61.760 2.730 65.200 ;
    END
  END enb
  OBS
      LAYER pwell ;
        RECT 17.900 65.610 27.930 71.670 ;
        RECT 35.875 65.570 41.725 71.670 ;
        RECT 47.400 65.610 57.430 71.670 ;
        RECT 65.375 65.570 71.225 71.670 ;
        RECT 76.900 65.610 86.930 71.670 ;
        RECT 94.875 65.570 100.725 71.670 ;
        RECT 106.400 65.610 116.430 71.670 ;
        RECT 124.375 65.570 130.225 71.670 ;
        RECT 135.900 65.610 145.930 71.670 ;
        RECT 153.875 65.570 159.725 71.670 ;
        RECT 3.820 61.285 5.625 61.515 ;
        RECT 3.335 60.605 5.625 61.285 ;
        RECT 3.480 60.415 3.650 60.605 ;
        RECT 7.645 60.415 7.815 60.585 ;
        RECT 24.550 54.760 34.580 61.160 ;
        RECT 40.255 59.925 46.105 60.865 ;
        RECT 40.255 59.875 46.110 59.925 ;
        RECT 40.260 54.765 46.110 59.875 ;
        RECT 54.050 54.760 64.080 61.160 ;
        RECT 69.755 59.925 75.605 60.865 ;
        RECT 69.755 59.875 75.610 59.925 ;
        RECT 69.760 54.765 75.610 59.875 ;
        RECT 83.550 54.760 93.580 61.160 ;
        RECT 99.255 59.925 105.105 60.865 ;
        RECT 99.255 59.875 105.110 59.925 ;
        RECT 99.260 54.765 105.110 59.875 ;
        RECT 113.050 54.760 123.080 61.160 ;
        RECT 128.755 59.925 134.605 60.865 ;
        RECT 128.755 59.875 134.610 59.925 ;
        RECT 128.760 54.765 134.610 59.875 ;
        RECT 142.550 54.760 152.580 61.160 ;
        RECT 158.255 59.925 164.105 60.865 ;
        RECT 158.255 59.875 164.110 59.925 ;
        RECT 158.260 54.765 164.110 59.875 ;
        RECT 2.300 44.805 8.150 49.915 ;
        RECT 2.300 44.755 8.155 44.805 ;
        RECT 2.305 43.815 8.155 44.755 ;
        RECT 13.830 43.520 23.860 49.920 ;
        RECT 31.800 44.805 37.650 49.915 ;
        RECT 31.800 44.755 37.655 44.805 ;
        RECT 31.805 43.815 37.655 44.755 ;
        RECT 43.330 43.520 53.360 49.920 ;
        RECT 61.300 44.805 67.150 49.915 ;
        RECT 61.300 44.755 67.155 44.805 ;
        RECT 61.305 43.815 67.155 44.755 ;
        RECT 72.830 43.520 82.860 49.920 ;
        RECT 90.800 44.805 96.650 49.915 ;
        RECT 90.800 44.755 96.655 44.805 ;
        RECT 90.805 43.815 96.655 44.755 ;
        RECT 102.330 43.520 112.360 49.920 ;
        RECT 120.300 44.805 126.150 49.915 ;
        RECT 120.300 44.755 126.155 44.805 ;
        RECT 120.305 43.815 126.155 44.755 ;
        RECT 131.830 43.520 141.860 49.920 ;
        RECT 149.800 44.805 155.650 49.915 ;
        RECT 149.800 44.755 155.655 44.805 ;
        RECT 149.805 43.815 155.655 44.755 ;
        RECT 161.330 43.520 171.360 49.920 ;
        RECT 6.685 33.010 12.535 39.110 ;
        RECT 20.480 33.010 30.510 39.070 ;
        RECT 36.185 33.010 42.035 39.110 ;
        RECT 49.980 33.010 60.010 39.070 ;
        RECT 65.685 33.010 71.535 39.110 ;
        RECT 79.480 33.010 89.510 39.070 ;
        RECT 95.185 33.010 101.035 39.110 ;
        RECT 108.980 33.010 119.010 39.070 ;
        RECT 124.685 33.010 130.535 39.110 ;
        RECT 138.480 33.010 148.510 39.070 ;
        RECT 154.185 33.010 160.035 39.110 ;
        RECT 167.980 33.010 178.010 39.070 ;
      LAYER li1 ;
        RECT 15.430 73.000 166.090 73.500 ;
        RECT 3.850 63.305 4.820 63.460 ;
        RECT 7.850 63.305 8.820 63.460 ;
        RECT 3.330 63.135 5.630 63.305 ;
        RECT 7.500 63.135 8.880 63.305 ;
        RECT 3.415 62.565 3.675 62.965 ;
        RECT 3.845 62.735 4.780 63.135 ;
        RECT 4.950 62.625 5.545 62.965 ;
        RECT 3.415 62.395 4.780 62.565 ;
        RECT 3.415 62.100 3.875 62.225 ;
        RECT 2.400 61.800 3.875 62.100 ;
        RECT 3.415 61.495 3.875 61.800 ;
        RECT 4.045 61.325 4.780 62.395 ;
        RECT 3.415 61.155 4.780 61.325 ;
        RECT 4.950 61.305 5.125 62.625 ;
        RECT 5.840 62.455 7.290 62.675 ;
        RECT 5.305 62.375 7.290 62.455 ;
        RECT 7.775 62.410 8.105 63.135 ;
        RECT 5.305 62.155 6.140 62.375 ;
        RECT 6.990 62.240 7.290 62.375 ;
        RECT 5.305 61.475 5.545 62.155 ;
        RECT 4.950 61.175 5.545 61.305 ;
        RECT 6.370 61.175 6.670 62.010 ;
        RECT 6.990 61.940 8.105 62.240 ;
        RECT 3.415 60.755 3.675 61.155 ;
        RECT 3.845 60.585 4.780 60.985 ;
        RECT 4.950 60.875 6.670 61.175 ;
        RECT 4.950 60.755 5.545 60.875 ;
        RECT 7.585 60.755 8.105 61.940 ;
        RECT 8.275 61.415 8.795 62.965 ;
        RECT 8.275 60.585 8.615 61.245 ;
        RECT 3.330 60.415 5.630 60.585 ;
        RECT 7.500 60.415 8.880 60.585 ;
        RECT 15.510 53.500 16.010 73.000 ;
        RECT 18.080 71.140 20.425 71.620 ;
        RECT 21.490 71.140 24.350 71.620 ;
        RECT 25.405 71.140 27.750 71.620 ;
        RECT 36.055 71.140 38.400 71.620 ;
        RECT 39.200 71.140 41.545 71.620 ;
        RECT 47.580 71.140 49.925 71.620 ;
        RECT 50.990 71.140 53.850 71.620 ;
        RECT 54.905 71.140 57.250 71.620 ;
        RECT 65.555 71.140 67.900 71.620 ;
        RECT 68.700 71.140 71.045 71.620 ;
        RECT 77.080 71.140 79.425 71.620 ;
        RECT 80.490 71.140 83.350 71.620 ;
        RECT 84.405 71.140 86.750 71.620 ;
        RECT 95.055 71.140 97.400 71.620 ;
        RECT 98.200 71.140 100.545 71.620 ;
        RECT 106.580 71.140 108.925 71.620 ;
        RECT 109.990 71.140 112.850 71.620 ;
        RECT 113.905 71.140 116.250 71.620 ;
        RECT 124.555 71.140 126.900 71.620 ;
        RECT 127.700 71.140 130.045 71.620 ;
        RECT 136.080 71.140 138.425 71.620 ;
        RECT 139.490 71.140 142.350 71.620 ;
        RECT 143.405 71.140 145.750 71.620 ;
        RECT 154.055 71.140 156.400 71.620 ;
        RECT 157.200 71.140 159.545 71.620 ;
        RECT 18.590 66.545 18.880 71.140 ;
        RECT 18.650 66.300 18.820 66.545 ;
        RECT 18.800 64.090 19.930 65.090 ;
        RECT 20.680 64.780 20.970 70.840 ;
        RECT 22.770 66.545 23.060 71.140 ;
        RECT 22.830 66.300 23.000 66.545 ;
        RECT 24.860 64.880 25.150 70.840 ;
        RECT 26.950 66.545 27.240 71.140 ;
        RECT 28.910 68.755 31.255 68.900 ;
        RECT 32.055 68.755 34.400 68.900 ;
        RECT 28.910 68.585 34.400 68.755 ;
        RECT 28.910 68.420 31.255 68.585 ;
        RECT 32.055 68.420 34.400 68.585 ;
        RECT 27.010 66.535 27.205 66.545 ;
        RECT 27.010 66.300 27.180 66.535 ;
        RECT 24.860 64.780 25.680 64.880 ;
        RECT 20.680 64.280 25.680 64.780 ;
        RECT 18.080 58.020 18.250 62.875 ;
        RECT 18.590 58.020 18.880 62.870 ;
        RECT 20.680 58.330 20.970 64.280 ;
        RECT 28.910 63.760 29.080 68.420 ;
        RECT 29.420 63.590 29.710 68.420 ;
        RECT 31.510 63.150 31.800 68.150 ;
        RECT 33.600 63.590 33.890 68.420 ;
        RECT 34.230 63.820 34.400 68.420 ;
        RECT 36.565 66.790 36.855 71.140 ;
        RECT 36.800 64.880 38.000 65.190 ;
        RECT 36.300 64.260 38.000 64.880 ;
        RECT 36.800 64.060 38.000 64.260 ;
        RECT 38.650 63.150 38.945 70.830 ;
        RECT 40.745 66.790 41.035 71.140 ;
        RECT 43.835 68.870 45.930 68.900 ;
        RECT 43.680 68.705 45.930 68.870 ;
        RECT 42.530 68.535 45.930 68.705 ;
        RECT 42.530 65.560 42.700 68.535 ;
        RECT 43.680 68.450 45.930 68.535 ;
        RECT 43.835 68.420 45.930 68.450 ;
        RECT 43.035 64.975 43.330 68.050 ;
        RECT 42.805 64.195 43.545 64.975 ;
        RECT 22.770 58.020 23.060 62.870 ;
        RECT 23.400 58.020 23.570 62.875 ;
        RECT 28.870 62.650 41.465 63.150 ;
        RECT 28.870 61.210 29.370 62.650 ;
        RECT 30.400 61.620 34.400 62.220 ;
        RECT 32.400 61.500 34.400 61.620 ;
        RECT 27.330 60.920 31.800 61.210 ;
        RECT 32.400 60.920 33.600 61.500 ;
        RECT 25.300 59.895 25.470 60.130 ;
        RECT 25.275 59.885 25.470 59.895 ;
        RECT 18.080 57.895 20.425 58.020 ;
        RECT 21.225 57.990 23.570 58.020 ;
        RECT 21.225 57.895 23.750 57.990 ;
        RECT 18.080 57.725 23.750 57.895 ;
        RECT 18.080 57.540 20.425 57.725 ;
        RECT 21.225 57.570 23.750 57.725 ;
        RECT 21.225 57.540 23.570 57.570 ;
        RECT 25.240 55.300 25.530 59.885 ;
        RECT 27.330 55.590 27.620 60.920 ;
        RECT 29.480 59.885 29.650 60.110 ;
        RECT 29.420 55.300 29.710 59.885 ;
        RECT 31.510 55.590 31.800 60.920 ;
        RECT 33.660 59.885 33.830 60.110 ;
        RECT 33.600 55.300 33.890 59.885 ;
        RECT 36.055 58.020 36.225 61.945 ;
        RECT 36.565 58.020 36.855 62.090 ;
        RECT 38.655 58.385 38.950 62.650 ;
        RECT 36.055 57.990 38.150 58.020 ;
        RECT 36.055 57.900 38.305 57.990 ;
        RECT 39.285 57.900 39.455 61.935 ;
        RECT 40.965 61.500 41.465 62.650 ;
        RECT 36.055 57.730 39.455 57.900 ;
        RECT 36.055 57.570 38.305 57.730 ;
        RECT 36.055 57.540 38.150 57.570 ;
        RECT 40.950 55.300 41.240 59.645 ;
        RECT 43.035 55.605 43.330 64.195 ;
        RECT 45.130 64.010 45.420 68.420 ;
        RECT 45.760 64.005 45.930 68.420 ;
        RECT 48.090 66.545 48.380 71.140 ;
        RECT 48.150 66.300 48.320 66.545 ;
        RECT 48.300 64.090 49.430 65.090 ;
        RECT 50.180 64.780 50.470 70.840 ;
        RECT 52.270 66.545 52.560 71.140 ;
        RECT 52.330 66.300 52.500 66.545 ;
        RECT 54.360 64.880 54.650 70.840 ;
        RECT 56.450 66.545 56.740 71.140 ;
        RECT 58.410 68.755 60.755 68.900 ;
        RECT 61.555 68.755 63.900 68.900 ;
        RECT 58.410 68.585 63.900 68.755 ;
        RECT 58.410 68.420 60.755 68.585 ;
        RECT 61.555 68.420 63.900 68.585 ;
        RECT 56.510 66.535 56.705 66.545 ;
        RECT 56.510 66.300 56.680 66.535 ;
        RECT 54.360 64.780 55.180 64.880 ;
        RECT 50.180 64.280 55.180 64.780 ;
        RECT 43.950 62.160 45.130 62.360 ;
        RECT 43.950 61.560 45.630 62.160 ;
        RECT 43.950 61.280 45.130 61.560 ;
        RECT 45.130 55.300 45.420 59.645 ;
        RECT 47.580 58.020 47.750 62.875 ;
        RECT 48.090 58.020 48.380 62.870 ;
        RECT 50.180 58.330 50.470 64.280 ;
        RECT 58.410 63.760 58.580 68.420 ;
        RECT 58.920 63.590 59.210 68.420 ;
        RECT 61.010 63.150 61.300 68.150 ;
        RECT 63.100 63.590 63.390 68.420 ;
        RECT 63.730 63.820 63.900 68.420 ;
        RECT 66.065 66.790 66.355 71.140 ;
        RECT 66.300 64.880 67.500 65.190 ;
        RECT 65.800 64.260 67.500 64.880 ;
        RECT 66.300 64.060 67.500 64.260 ;
        RECT 68.150 63.150 68.445 70.830 ;
        RECT 70.245 66.790 70.535 71.140 ;
        RECT 73.335 68.870 75.430 68.900 ;
        RECT 73.180 68.705 75.430 68.870 ;
        RECT 72.030 68.535 75.430 68.705 ;
        RECT 72.030 65.560 72.200 68.535 ;
        RECT 73.180 68.450 75.430 68.535 ;
        RECT 73.335 68.420 75.430 68.450 ;
        RECT 72.535 64.975 72.830 68.050 ;
        RECT 72.305 64.195 73.045 64.975 ;
        RECT 52.270 58.020 52.560 62.870 ;
        RECT 52.900 58.020 53.070 62.875 ;
        RECT 58.370 62.650 70.965 63.150 ;
        RECT 58.370 61.210 58.870 62.650 ;
        RECT 59.900 61.620 63.900 62.220 ;
        RECT 61.900 61.500 63.900 61.620 ;
        RECT 56.830 60.920 61.300 61.210 ;
        RECT 61.900 60.920 63.100 61.500 ;
        RECT 54.800 59.895 54.970 60.130 ;
        RECT 54.775 59.885 54.970 59.895 ;
        RECT 47.580 57.895 49.925 58.020 ;
        RECT 50.725 57.990 53.070 58.020 ;
        RECT 50.725 57.895 53.250 57.990 ;
        RECT 47.580 57.725 53.250 57.895 ;
        RECT 47.580 57.540 49.925 57.725 ;
        RECT 50.725 57.570 53.250 57.725 ;
        RECT 50.725 57.540 53.070 57.570 ;
        RECT 54.740 55.300 55.030 59.885 ;
        RECT 56.830 55.590 57.120 60.920 ;
        RECT 58.980 59.885 59.150 60.110 ;
        RECT 58.920 55.300 59.210 59.885 ;
        RECT 61.010 55.590 61.300 60.920 ;
        RECT 63.160 59.885 63.330 60.110 ;
        RECT 63.100 55.300 63.390 59.885 ;
        RECT 65.555 58.020 65.725 61.945 ;
        RECT 66.065 58.020 66.355 62.090 ;
        RECT 68.155 58.385 68.450 62.650 ;
        RECT 65.555 57.990 67.650 58.020 ;
        RECT 65.555 57.900 67.805 57.990 ;
        RECT 68.785 57.900 68.955 61.935 ;
        RECT 70.465 61.500 70.965 62.650 ;
        RECT 65.555 57.730 68.955 57.900 ;
        RECT 65.555 57.570 67.805 57.730 ;
        RECT 65.555 57.540 67.650 57.570 ;
        RECT 70.450 55.300 70.740 59.645 ;
        RECT 72.535 55.605 72.830 64.195 ;
        RECT 74.630 64.010 74.920 68.420 ;
        RECT 75.260 64.005 75.430 68.420 ;
        RECT 77.590 66.545 77.880 71.140 ;
        RECT 77.650 66.300 77.820 66.545 ;
        RECT 77.800 64.090 78.930 65.090 ;
        RECT 79.680 64.780 79.970 70.840 ;
        RECT 81.770 66.545 82.060 71.140 ;
        RECT 81.830 66.300 82.000 66.545 ;
        RECT 83.860 64.880 84.150 70.840 ;
        RECT 85.950 66.545 86.240 71.140 ;
        RECT 87.910 68.755 90.255 68.900 ;
        RECT 91.055 68.755 93.400 68.900 ;
        RECT 87.910 68.585 93.400 68.755 ;
        RECT 87.910 68.420 90.255 68.585 ;
        RECT 91.055 68.420 93.400 68.585 ;
        RECT 86.010 66.535 86.205 66.545 ;
        RECT 86.010 66.300 86.180 66.535 ;
        RECT 83.860 64.780 84.680 64.880 ;
        RECT 79.680 64.280 84.680 64.780 ;
        RECT 73.450 62.160 74.630 62.360 ;
        RECT 73.450 61.560 75.130 62.160 ;
        RECT 73.450 61.280 74.630 61.560 ;
        RECT 74.630 55.300 74.920 59.645 ;
        RECT 77.080 58.020 77.250 62.875 ;
        RECT 77.590 58.020 77.880 62.870 ;
        RECT 79.680 58.330 79.970 64.280 ;
        RECT 87.910 63.760 88.080 68.420 ;
        RECT 88.420 63.590 88.710 68.420 ;
        RECT 90.510 63.150 90.800 68.150 ;
        RECT 92.600 63.590 92.890 68.420 ;
        RECT 93.230 63.820 93.400 68.420 ;
        RECT 95.565 66.790 95.855 71.140 ;
        RECT 95.800 64.880 97.000 65.190 ;
        RECT 95.300 64.260 97.000 64.880 ;
        RECT 95.800 64.060 97.000 64.260 ;
        RECT 97.650 63.150 97.945 70.830 ;
        RECT 99.745 66.790 100.035 71.140 ;
        RECT 102.835 68.870 104.930 68.900 ;
        RECT 102.680 68.705 104.930 68.870 ;
        RECT 101.530 68.535 104.930 68.705 ;
        RECT 101.530 65.560 101.700 68.535 ;
        RECT 102.680 68.450 104.930 68.535 ;
        RECT 102.835 68.420 104.930 68.450 ;
        RECT 102.035 64.975 102.330 68.050 ;
        RECT 101.805 64.195 102.545 64.975 ;
        RECT 81.770 58.020 82.060 62.870 ;
        RECT 82.400 58.020 82.570 62.875 ;
        RECT 87.870 62.650 100.465 63.150 ;
        RECT 87.870 61.210 88.370 62.650 ;
        RECT 89.400 61.620 93.400 62.220 ;
        RECT 91.400 61.500 93.400 61.620 ;
        RECT 86.330 60.920 90.800 61.210 ;
        RECT 91.400 60.920 92.600 61.500 ;
        RECT 84.300 59.895 84.470 60.130 ;
        RECT 84.275 59.885 84.470 59.895 ;
        RECT 77.080 57.895 79.425 58.020 ;
        RECT 80.225 57.990 82.570 58.020 ;
        RECT 80.225 57.895 82.750 57.990 ;
        RECT 77.080 57.725 82.750 57.895 ;
        RECT 77.080 57.540 79.425 57.725 ;
        RECT 80.225 57.570 82.750 57.725 ;
        RECT 80.225 57.540 82.570 57.570 ;
        RECT 84.240 55.300 84.530 59.885 ;
        RECT 86.330 55.590 86.620 60.920 ;
        RECT 88.480 59.885 88.650 60.110 ;
        RECT 88.420 55.300 88.710 59.885 ;
        RECT 90.510 55.590 90.800 60.920 ;
        RECT 92.660 59.885 92.830 60.110 ;
        RECT 92.600 55.300 92.890 59.885 ;
        RECT 95.055 58.020 95.225 61.945 ;
        RECT 95.565 58.020 95.855 62.090 ;
        RECT 97.655 58.385 97.950 62.650 ;
        RECT 95.055 57.990 97.150 58.020 ;
        RECT 95.055 57.900 97.305 57.990 ;
        RECT 98.285 57.900 98.455 61.935 ;
        RECT 99.965 61.500 100.465 62.650 ;
        RECT 95.055 57.730 98.455 57.900 ;
        RECT 95.055 57.570 97.305 57.730 ;
        RECT 95.055 57.540 97.150 57.570 ;
        RECT 99.950 55.300 100.240 59.645 ;
        RECT 102.035 55.605 102.330 64.195 ;
        RECT 104.130 64.010 104.420 68.420 ;
        RECT 104.760 64.005 104.930 68.420 ;
        RECT 107.090 66.545 107.380 71.140 ;
        RECT 107.150 66.300 107.320 66.545 ;
        RECT 107.300 64.090 108.430 65.090 ;
        RECT 109.180 64.780 109.470 70.840 ;
        RECT 111.270 66.545 111.560 71.140 ;
        RECT 111.330 66.300 111.500 66.545 ;
        RECT 113.360 64.880 113.650 70.840 ;
        RECT 115.450 66.545 115.740 71.140 ;
        RECT 117.410 68.755 119.755 68.900 ;
        RECT 120.555 68.755 122.900 68.900 ;
        RECT 117.410 68.585 122.900 68.755 ;
        RECT 117.410 68.420 119.755 68.585 ;
        RECT 120.555 68.420 122.900 68.585 ;
        RECT 115.510 66.535 115.705 66.545 ;
        RECT 115.510 66.300 115.680 66.535 ;
        RECT 113.360 64.780 114.180 64.880 ;
        RECT 109.180 64.280 114.180 64.780 ;
        RECT 102.950 62.160 104.130 62.360 ;
        RECT 102.950 61.560 104.630 62.160 ;
        RECT 102.950 61.280 104.130 61.560 ;
        RECT 104.130 55.300 104.420 59.645 ;
        RECT 106.580 58.020 106.750 62.875 ;
        RECT 107.090 58.020 107.380 62.870 ;
        RECT 109.180 58.330 109.470 64.280 ;
        RECT 117.410 63.760 117.580 68.420 ;
        RECT 117.920 63.590 118.210 68.420 ;
        RECT 120.010 63.150 120.300 68.150 ;
        RECT 122.100 63.590 122.390 68.420 ;
        RECT 122.730 63.820 122.900 68.420 ;
        RECT 125.065 66.790 125.355 71.140 ;
        RECT 125.300 64.880 126.500 65.190 ;
        RECT 124.800 64.260 126.500 64.880 ;
        RECT 125.300 64.060 126.500 64.260 ;
        RECT 127.150 63.150 127.445 70.830 ;
        RECT 129.245 66.790 129.535 71.140 ;
        RECT 132.335 68.870 134.430 68.900 ;
        RECT 132.180 68.705 134.430 68.870 ;
        RECT 131.030 68.535 134.430 68.705 ;
        RECT 131.030 65.560 131.200 68.535 ;
        RECT 132.180 68.450 134.430 68.535 ;
        RECT 132.335 68.420 134.430 68.450 ;
        RECT 131.535 64.975 131.830 68.050 ;
        RECT 131.305 64.195 132.045 64.975 ;
        RECT 111.270 58.020 111.560 62.870 ;
        RECT 111.900 58.020 112.070 62.875 ;
        RECT 117.370 62.650 129.965 63.150 ;
        RECT 117.370 61.210 117.870 62.650 ;
        RECT 118.900 61.620 122.900 62.220 ;
        RECT 120.900 61.500 122.900 61.620 ;
        RECT 115.830 60.920 120.300 61.210 ;
        RECT 120.900 60.920 122.100 61.500 ;
        RECT 113.800 59.895 113.970 60.130 ;
        RECT 113.775 59.885 113.970 59.895 ;
        RECT 106.580 57.895 108.925 58.020 ;
        RECT 109.725 57.990 112.070 58.020 ;
        RECT 109.725 57.895 112.250 57.990 ;
        RECT 106.580 57.725 112.250 57.895 ;
        RECT 106.580 57.540 108.925 57.725 ;
        RECT 109.725 57.570 112.250 57.725 ;
        RECT 109.725 57.540 112.070 57.570 ;
        RECT 113.740 55.300 114.030 59.885 ;
        RECT 115.830 55.590 116.120 60.920 ;
        RECT 117.980 59.885 118.150 60.110 ;
        RECT 117.920 55.300 118.210 59.885 ;
        RECT 120.010 55.590 120.300 60.920 ;
        RECT 122.160 59.885 122.330 60.110 ;
        RECT 122.100 55.300 122.390 59.885 ;
        RECT 124.555 58.020 124.725 61.945 ;
        RECT 125.065 58.020 125.355 62.090 ;
        RECT 127.155 58.385 127.450 62.650 ;
        RECT 124.555 57.990 126.650 58.020 ;
        RECT 124.555 57.900 126.805 57.990 ;
        RECT 127.785 57.900 127.955 61.935 ;
        RECT 129.465 61.500 129.965 62.650 ;
        RECT 124.555 57.730 127.955 57.900 ;
        RECT 124.555 57.570 126.805 57.730 ;
        RECT 124.555 57.540 126.650 57.570 ;
        RECT 129.450 55.300 129.740 59.645 ;
        RECT 131.535 55.605 131.830 64.195 ;
        RECT 133.630 64.010 133.920 68.420 ;
        RECT 134.260 64.005 134.430 68.420 ;
        RECT 136.590 66.545 136.880 71.140 ;
        RECT 136.650 66.300 136.820 66.545 ;
        RECT 136.800 64.090 137.930 65.090 ;
        RECT 138.680 64.780 138.970 70.840 ;
        RECT 140.770 66.545 141.060 71.140 ;
        RECT 140.830 66.300 141.000 66.545 ;
        RECT 142.860 64.880 143.150 70.840 ;
        RECT 144.950 66.545 145.240 71.140 ;
        RECT 146.910 68.755 149.255 68.900 ;
        RECT 150.055 68.755 152.400 68.900 ;
        RECT 146.910 68.585 152.400 68.755 ;
        RECT 146.910 68.420 149.255 68.585 ;
        RECT 150.055 68.420 152.400 68.585 ;
        RECT 145.010 66.535 145.205 66.545 ;
        RECT 145.010 66.300 145.180 66.535 ;
        RECT 142.860 64.780 143.680 64.880 ;
        RECT 138.680 64.280 143.680 64.780 ;
        RECT 132.450 62.160 133.630 62.360 ;
        RECT 132.450 61.560 134.130 62.160 ;
        RECT 132.450 61.280 133.630 61.560 ;
        RECT 133.630 55.300 133.920 59.645 ;
        RECT 136.080 58.020 136.250 62.875 ;
        RECT 136.590 58.020 136.880 62.870 ;
        RECT 138.680 58.330 138.970 64.280 ;
        RECT 146.910 63.760 147.080 68.420 ;
        RECT 147.420 63.590 147.710 68.420 ;
        RECT 149.510 63.150 149.800 68.150 ;
        RECT 151.600 63.590 151.890 68.420 ;
        RECT 152.230 63.820 152.400 68.420 ;
        RECT 154.565 66.790 154.855 71.140 ;
        RECT 154.800 64.880 156.000 65.190 ;
        RECT 154.300 64.260 156.000 64.880 ;
        RECT 154.800 64.060 156.000 64.260 ;
        RECT 156.650 63.150 156.945 70.830 ;
        RECT 158.745 66.790 159.035 71.140 ;
        RECT 161.835 68.870 163.930 68.900 ;
        RECT 161.680 68.705 163.930 68.870 ;
        RECT 160.530 68.535 163.930 68.705 ;
        RECT 160.530 65.560 160.700 68.535 ;
        RECT 161.680 68.450 163.930 68.535 ;
        RECT 161.835 68.420 163.930 68.450 ;
        RECT 161.035 64.975 161.330 68.050 ;
        RECT 160.805 64.195 161.545 64.975 ;
        RECT 140.770 58.020 141.060 62.870 ;
        RECT 141.400 58.020 141.570 62.875 ;
        RECT 146.870 62.650 159.465 63.150 ;
        RECT 146.870 61.210 147.370 62.650 ;
        RECT 148.400 61.620 152.400 62.220 ;
        RECT 150.400 61.500 152.400 61.620 ;
        RECT 145.330 60.920 149.800 61.210 ;
        RECT 150.400 60.920 151.600 61.500 ;
        RECT 143.300 59.895 143.470 60.130 ;
        RECT 143.275 59.885 143.470 59.895 ;
        RECT 136.080 57.895 138.425 58.020 ;
        RECT 139.225 57.990 141.570 58.020 ;
        RECT 139.225 57.895 141.750 57.990 ;
        RECT 136.080 57.725 141.750 57.895 ;
        RECT 136.080 57.540 138.425 57.725 ;
        RECT 139.225 57.570 141.750 57.725 ;
        RECT 139.225 57.540 141.570 57.570 ;
        RECT 143.240 55.300 143.530 59.885 ;
        RECT 145.330 55.590 145.620 60.920 ;
        RECT 147.480 59.885 147.650 60.110 ;
        RECT 147.420 55.300 147.710 59.885 ;
        RECT 149.510 55.590 149.800 60.920 ;
        RECT 151.660 59.885 151.830 60.110 ;
        RECT 151.600 55.300 151.890 59.885 ;
        RECT 154.055 58.020 154.225 61.945 ;
        RECT 154.565 58.020 154.855 62.090 ;
        RECT 156.655 58.385 156.950 62.650 ;
        RECT 154.055 57.990 156.150 58.020 ;
        RECT 154.055 57.900 156.305 57.990 ;
        RECT 157.285 57.900 157.455 61.935 ;
        RECT 158.965 61.500 159.465 62.650 ;
        RECT 154.055 57.730 157.455 57.900 ;
        RECT 154.055 57.570 156.305 57.730 ;
        RECT 154.055 57.540 156.150 57.570 ;
        RECT 158.950 55.300 159.240 59.645 ;
        RECT 161.035 55.605 161.330 64.195 ;
        RECT 163.130 64.010 163.420 68.420 ;
        RECT 163.760 64.005 163.930 68.420 ;
        RECT 161.950 62.160 163.130 62.360 ;
        RECT 161.950 61.560 163.630 62.160 ;
        RECT 161.950 61.280 163.130 61.560 ;
        RECT 163.130 55.300 163.420 59.645 ;
        RECT 24.730 54.820 27.080 55.300 ;
        RECT 28.130 54.820 30.990 55.300 ;
        RECT 32.055 54.820 34.400 55.300 ;
        RECT 40.440 55.270 42.780 55.300 ;
        RECT 43.590 55.270 45.930 55.300 ;
        RECT 40.440 54.850 42.785 55.270 ;
        RECT 43.585 54.850 45.930 55.270 ;
        RECT 40.440 54.820 42.780 54.850 ;
        RECT 43.590 54.820 45.930 54.850 ;
        RECT 54.230 54.820 56.580 55.300 ;
        RECT 57.630 54.820 60.490 55.300 ;
        RECT 61.555 54.820 63.900 55.300 ;
        RECT 69.940 55.270 72.280 55.300 ;
        RECT 73.090 55.270 75.430 55.300 ;
        RECT 69.940 54.850 72.285 55.270 ;
        RECT 73.085 54.850 75.430 55.270 ;
        RECT 69.940 54.820 72.280 54.850 ;
        RECT 73.090 54.820 75.430 54.850 ;
        RECT 83.730 54.820 86.080 55.300 ;
        RECT 87.130 54.820 89.990 55.300 ;
        RECT 91.055 54.820 93.400 55.300 ;
        RECT 99.440 55.270 101.780 55.300 ;
        RECT 102.590 55.270 104.930 55.300 ;
        RECT 99.440 54.850 101.785 55.270 ;
        RECT 102.585 54.850 104.930 55.270 ;
        RECT 99.440 54.820 101.780 54.850 ;
        RECT 102.590 54.820 104.930 54.850 ;
        RECT 113.230 54.820 115.580 55.300 ;
        RECT 116.630 54.820 119.490 55.300 ;
        RECT 120.555 54.820 122.900 55.300 ;
        RECT 128.940 55.270 131.280 55.300 ;
        RECT 132.090 55.270 134.430 55.300 ;
        RECT 128.940 54.850 131.285 55.270 ;
        RECT 132.085 54.850 134.430 55.270 ;
        RECT 128.940 54.820 131.280 54.850 ;
        RECT 132.090 54.820 134.430 54.850 ;
        RECT 142.730 54.820 145.080 55.300 ;
        RECT 146.130 54.820 148.990 55.300 ;
        RECT 150.055 54.820 152.400 55.300 ;
        RECT 158.440 55.270 160.780 55.300 ;
        RECT 161.590 55.270 163.930 55.300 ;
        RECT 158.440 54.850 160.785 55.270 ;
        RECT 161.585 54.850 163.930 55.270 ;
        RECT 158.440 54.820 160.780 54.850 ;
        RECT 161.590 54.820 163.930 54.850 ;
        RECT 165.510 53.500 166.010 73.000 ;
        RECT 15.430 53.000 166.090 53.500 ;
        RECT 0.430 51.000 180.090 51.500 ;
        RECT 0.510 31.500 1.010 51.000 ;
        RECT 2.480 49.830 4.820 49.860 ;
        RECT 5.630 49.830 7.970 49.860 ;
        RECT 2.480 49.410 4.825 49.830 ;
        RECT 5.625 49.410 7.970 49.830 ;
        RECT 2.480 49.380 4.820 49.410 ;
        RECT 5.630 49.380 7.970 49.410 ;
        RECT 14.010 49.380 16.355 49.860 ;
        RECT 17.420 49.380 20.280 49.860 ;
        RECT 21.330 49.380 23.680 49.860 ;
        RECT 31.980 49.830 34.320 49.860 ;
        RECT 35.130 49.830 37.470 49.860 ;
        RECT 31.980 49.410 34.325 49.830 ;
        RECT 35.125 49.410 37.470 49.830 ;
        RECT 31.980 49.380 34.320 49.410 ;
        RECT 35.130 49.380 37.470 49.410 ;
        RECT 43.510 49.380 45.855 49.860 ;
        RECT 46.920 49.380 49.780 49.860 ;
        RECT 50.830 49.380 53.180 49.860 ;
        RECT 61.480 49.830 63.820 49.860 ;
        RECT 64.630 49.830 66.970 49.860 ;
        RECT 61.480 49.410 63.825 49.830 ;
        RECT 64.625 49.410 66.970 49.830 ;
        RECT 61.480 49.380 63.820 49.410 ;
        RECT 64.630 49.380 66.970 49.410 ;
        RECT 73.010 49.380 75.355 49.860 ;
        RECT 76.420 49.380 79.280 49.860 ;
        RECT 80.330 49.380 82.680 49.860 ;
        RECT 90.980 49.830 93.320 49.860 ;
        RECT 94.130 49.830 96.470 49.860 ;
        RECT 90.980 49.410 93.325 49.830 ;
        RECT 94.125 49.410 96.470 49.830 ;
        RECT 90.980 49.380 93.320 49.410 ;
        RECT 94.130 49.380 96.470 49.410 ;
        RECT 102.510 49.380 104.855 49.860 ;
        RECT 105.920 49.380 108.780 49.860 ;
        RECT 109.830 49.380 112.180 49.860 ;
        RECT 120.480 49.830 122.820 49.860 ;
        RECT 123.630 49.830 125.970 49.860 ;
        RECT 120.480 49.410 122.825 49.830 ;
        RECT 123.625 49.410 125.970 49.830 ;
        RECT 120.480 49.380 122.820 49.410 ;
        RECT 123.630 49.380 125.970 49.410 ;
        RECT 132.010 49.380 134.355 49.860 ;
        RECT 135.420 49.380 138.280 49.860 ;
        RECT 139.330 49.380 141.680 49.860 ;
        RECT 149.980 49.830 152.320 49.860 ;
        RECT 153.130 49.830 155.470 49.860 ;
        RECT 149.980 49.410 152.325 49.830 ;
        RECT 153.125 49.410 155.470 49.830 ;
        RECT 149.980 49.380 152.320 49.410 ;
        RECT 153.130 49.380 155.470 49.410 ;
        RECT 161.510 49.380 163.855 49.860 ;
        RECT 164.920 49.380 167.780 49.860 ;
        RECT 168.830 49.380 171.180 49.860 ;
        RECT 2.990 45.035 3.280 49.380 ;
        RECT 3.280 43.120 4.460 43.400 ;
        RECT 2.780 42.520 4.460 43.120 ;
        RECT 3.280 42.320 4.460 42.520 ;
        RECT 2.480 36.260 2.650 40.675 ;
        RECT 2.990 36.260 3.280 40.670 ;
        RECT 5.080 40.485 5.375 49.075 ;
        RECT 7.170 45.035 7.460 49.380 ;
        RECT 10.260 47.110 12.355 47.140 ;
        RECT 10.105 46.950 12.355 47.110 ;
        RECT 8.955 46.780 12.355 46.950 ;
        RECT 6.945 42.030 7.445 43.180 ;
        RECT 8.955 42.745 9.125 46.780 ;
        RECT 10.105 46.690 12.355 46.780 ;
        RECT 10.260 46.660 12.355 46.690 ;
        RECT 9.460 42.030 9.755 46.295 ;
        RECT 11.555 42.590 11.845 46.660 ;
        RECT 12.185 42.735 12.355 46.660 ;
        RECT 14.520 44.795 14.810 49.380 ;
        RECT 14.580 44.570 14.750 44.795 ;
        RECT 16.610 43.760 16.900 49.090 ;
        RECT 18.700 44.795 18.990 49.380 ;
        RECT 18.760 44.570 18.930 44.795 ;
        RECT 20.790 43.760 21.080 49.090 ;
        RECT 22.880 44.795 23.170 49.380 ;
        RECT 24.840 47.110 27.185 47.140 ;
        RECT 24.660 46.955 27.185 47.110 ;
        RECT 27.985 46.955 30.330 47.140 ;
        RECT 24.660 46.785 30.330 46.955 ;
        RECT 24.660 46.690 27.185 46.785 ;
        RECT 24.840 46.660 27.185 46.690 ;
        RECT 27.985 46.660 30.330 46.785 ;
        RECT 22.940 44.785 23.135 44.795 ;
        RECT 22.940 44.550 23.110 44.785 ;
        RECT 14.810 43.180 16.010 43.760 ;
        RECT 16.610 43.470 21.080 43.760 ;
        RECT 14.010 43.060 16.010 43.180 ;
        RECT 14.010 42.460 18.010 43.060 ;
        RECT 19.040 42.030 19.540 43.470 ;
        RECT 6.945 41.530 19.540 42.030 ;
        RECT 24.840 41.805 25.010 46.660 ;
        RECT 25.350 41.810 25.640 46.660 ;
        RECT 4.865 39.705 5.605 40.485 ;
        RECT 5.080 36.630 5.375 39.705 ;
        RECT 2.480 36.230 4.575 36.260 ;
        RECT 2.480 36.145 4.730 36.230 ;
        RECT 5.710 36.145 5.880 39.120 ;
        RECT 2.480 35.975 5.880 36.145 ;
        RECT 2.480 35.810 4.730 35.975 ;
        RECT 2.480 35.780 4.575 35.810 ;
        RECT 7.375 33.540 7.665 37.890 ;
        RECT 9.465 33.850 9.760 41.530 ;
        RECT 10.410 40.420 11.610 40.620 ;
        RECT 10.410 39.800 12.110 40.420 ;
        RECT 10.410 39.490 11.610 39.800 ;
        RECT 11.555 33.540 11.845 37.890 ;
        RECT 14.010 36.260 14.180 40.860 ;
        RECT 14.520 36.260 14.810 41.090 ;
        RECT 16.610 36.530 16.900 41.530 ;
        RECT 18.700 36.260 18.990 41.090 ;
        RECT 19.330 36.260 19.500 40.920 ;
        RECT 27.440 40.400 27.730 46.350 ;
        RECT 29.530 41.810 29.820 46.660 ;
        RECT 30.160 41.805 30.330 46.660 ;
        RECT 32.490 45.035 32.780 49.380 ;
        RECT 32.780 43.120 33.960 43.400 ;
        RECT 32.280 42.520 33.960 43.120 ;
        RECT 32.780 42.320 33.960 42.520 ;
        RECT 22.730 39.900 27.730 40.400 ;
        RECT 22.730 39.800 23.550 39.900 ;
        RECT 21.230 38.145 21.400 38.380 ;
        RECT 21.205 38.135 21.400 38.145 ;
        RECT 14.010 36.095 16.355 36.260 ;
        RECT 17.155 36.095 19.500 36.260 ;
        RECT 14.010 35.925 19.500 36.095 ;
        RECT 14.010 35.780 16.355 35.925 ;
        RECT 17.155 35.780 19.500 35.925 ;
        RECT 21.170 33.540 21.460 38.135 ;
        RECT 23.260 33.840 23.550 39.800 ;
        RECT 25.410 38.135 25.580 38.380 ;
        RECT 25.350 33.540 25.640 38.135 ;
        RECT 27.440 33.840 27.730 39.900 ;
        RECT 28.480 39.590 29.610 40.590 ;
        RECT 29.590 38.135 29.760 38.380 ;
        RECT 29.530 33.540 29.820 38.135 ;
        RECT 31.980 36.260 32.150 40.675 ;
        RECT 32.490 36.260 32.780 40.670 ;
        RECT 34.580 40.485 34.875 49.075 ;
        RECT 36.670 45.035 36.960 49.380 ;
        RECT 39.760 47.110 41.855 47.140 ;
        RECT 39.605 46.950 41.855 47.110 ;
        RECT 38.455 46.780 41.855 46.950 ;
        RECT 36.445 42.030 36.945 43.180 ;
        RECT 38.455 42.745 38.625 46.780 ;
        RECT 39.605 46.690 41.855 46.780 ;
        RECT 39.760 46.660 41.855 46.690 ;
        RECT 38.960 42.030 39.255 46.295 ;
        RECT 41.055 42.590 41.345 46.660 ;
        RECT 41.685 42.735 41.855 46.660 ;
        RECT 44.020 44.795 44.310 49.380 ;
        RECT 44.080 44.570 44.250 44.795 ;
        RECT 46.110 43.760 46.400 49.090 ;
        RECT 48.200 44.795 48.490 49.380 ;
        RECT 48.260 44.570 48.430 44.795 ;
        RECT 50.290 43.760 50.580 49.090 ;
        RECT 52.380 44.795 52.670 49.380 ;
        RECT 54.340 47.110 56.685 47.140 ;
        RECT 54.160 46.955 56.685 47.110 ;
        RECT 57.485 46.955 59.830 47.140 ;
        RECT 54.160 46.785 59.830 46.955 ;
        RECT 54.160 46.690 56.685 46.785 ;
        RECT 54.340 46.660 56.685 46.690 ;
        RECT 57.485 46.660 59.830 46.785 ;
        RECT 52.440 44.785 52.635 44.795 ;
        RECT 52.440 44.550 52.610 44.785 ;
        RECT 44.310 43.180 45.510 43.760 ;
        RECT 46.110 43.470 50.580 43.760 ;
        RECT 43.510 43.060 45.510 43.180 ;
        RECT 43.510 42.460 47.510 43.060 ;
        RECT 48.540 42.030 49.040 43.470 ;
        RECT 36.445 41.530 49.040 42.030 ;
        RECT 54.340 41.805 54.510 46.660 ;
        RECT 54.850 41.810 55.140 46.660 ;
        RECT 34.365 39.705 35.105 40.485 ;
        RECT 34.580 36.630 34.875 39.705 ;
        RECT 31.980 36.230 34.075 36.260 ;
        RECT 31.980 36.145 34.230 36.230 ;
        RECT 35.210 36.145 35.380 39.120 ;
        RECT 31.980 35.975 35.380 36.145 ;
        RECT 31.980 35.810 34.230 35.975 ;
        RECT 31.980 35.780 34.075 35.810 ;
        RECT 36.875 33.540 37.165 37.890 ;
        RECT 38.965 33.850 39.260 41.530 ;
        RECT 39.910 40.420 41.110 40.620 ;
        RECT 39.910 39.800 41.610 40.420 ;
        RECT 39.910 39.490 41.110 39.800 ;
        RECT 41.055 33.540 41.345 37.890 ;
        RECT 43.510 36.260 43.680 40.860 ;
        RECT 44.020 36.260 44.310 41.090 ;
        RECT 46.110 36.530 46.400 41.530 ;
        RECT 48.200 36.260 48.490 41.090 ;
        RECT 48.830 36.260 49.000 40.920 ;
        RECT 56.940 40.400 57.230 46.350 ;
        RECT 59.030 41.810 59.320 46.660 ;
        RECT 59.660 41.805 59.830 46.660 ;
        RECT 61.990 45.035 62.280 49.380 ;
        RECT 62.280 43.120 63.460 43.400 ;
        RECT 61.780 42.520 63.460 43.120 ;
        RECT 62.280 42.320 63.460 42.520 ;
        RECT 52.230 39.900 57.230 40.400 ;
        RECT 52.230 39.800 53.050 39.900 ;
        RECT 50.730 38.145 50.900 38.380 ;
        RECT 50.705 38.135 50.900 38.145 ;
        RECT 43.510 36.095 45.855 36.260 ;
        RECT 46.655 36.095 49.000 36.260 ;
        RECT 43.510 35.925 49.000 36.095 ;
        RECT 43.510 35.780 45.855 35.925 ;
        RECT 46.655 35.780 49.000 35.925 ;
        RECT 50.670 33.540 50.960 38.135 ;
        RECT 52.760 33.840 53.050 39.800 ;
        RECT 54.910 38.135 55.080 38.380 ;
        RECT 54.850 33.540 55.140 38.135 ;
        RECT 56.940 33.840 57.230 39.900 ;
        RECT 57.980 39.590 59.110 40.590 ;
        RECT 59.090 38.135 59.260 38.380 ;
        RECT 59.030 33.540 59.320 38.135 ;
        RECT 61.480 36.260 61.650 40.675 ;
        RECT 61.990 36.260 62.280 40.670 ;
        RECT 64.080 40.485 64.375 49.075 ;
        RECT 66.170 45.035 66.460 49.380 ;
        RECT 69.260 47.110 71.355 47.140 ;
        RECT 69.105 46.950 71.355 47.110 ;
        RECT 67.955 46.780 71.355 46.950 ;
        RECT 65.945 42.030 66.445 43.180 ;
        RECT 67.955 42.745 68.125 46.780 ;
        RECT 69.105 46.690 71.355 46.780 ;
        RECT 69.260 46.660 71.355 46.690 ;
        RECT 68.460 42.030 68.755 46.295 ;
        RECT 70.555 42.590 70.845 46.660 ;
        RECT 71.185 42.735 71.355 46.660 ;
        RECT 73.520 44.795 73.810 49.380 ;
        RECT 73.580 44.570 73.750 44.795 ;
        RECT 75.610 43.760 75.900 49.090 ;
        RECT 77.700 44.795 77.990 49.380 ;
        RECT 77.760 44.570 77.930 44.795 ;
        RECT 79.790 43.760 80.080 49.090 ;
        RECT 81.880 44.795 82.170 49.380 ;
        RECT 83.840 47.110 86.185 47.140 ;
        RECT 83.660 46.955 86.185 47.110 ;
        RECT 86.985 46.955 89.330 47.140 ;
        RECT 83.660 46.785 89.330 46.955 ;
        RECT 83.660 46.690 86.185 46.785 ;
        RECT 83.840 46.660 86.185 46.690 ;
        RECT 86.985 46.660 89.330 46.785 ;
        RECT 81.940 44.785 82.135 44.795 ;
        RECT 81.940 44.550 82.110 44.785 ;
        RECT 73.810 43.180 75.010 43.760 ;
        RECT 75.610 43.470 80.080 43.760 ;
        RECT 73.010 43.060 75.010 43.180 ;
        RECT 73.010 42.460 77.010 43.060 ;
        RECT 78.040 42.030 78.540 43.470 ;
        RECT 65.945 41.530 78.540 42.030 ;
        RECT 83.840 41.805 84.010 46.660 ;
        RECT 84.350 41.810 84.640 46.660 ;
        RECT 63.865 39.705 64.605 40.485 ;
        RECT 64.080 36.630 64.375 39.705 ;
        RECT 61.480 36.230 63.575 36.260 ;
        RECT 61.480 36.145 63.730 36.230 ;
        RECT 64.710 36.145 64.880 39.120 ;
        RECT 61.480 35.975 64.880 36.145 ;
        RECT 61.480 35.810 63.730 35.975 ;
        RECT 61.480 35.780 63.575 35.810 ;
        RECT 66.375 33.540 66.665 37.890 ;
        RECT 68.465 33.850 68.760 41.530 ;
        RECT 69.410 40.420 70.610 40.620 ;
        RECT 69.410 39.800 71.110 40.420 ;
        RECT 69.410 39.490 70.610 39.800 ;
        RECT 70.555 33.540 70.845 37.890 ;
        RECT 73.010 36.260 73.180 40.860 ;
        RECT 73.520 36.260 73.810 41.090 ;
        RECT 75.610 36.530 75.900 41.530 ;
        RECT 77.700 36.260 77.990 41.090 ;
        RECT 78.330 36.260 78.500 40.920 ;
        RECT 86.440 40.400 86.730 46.350 ;
        RECT 88.530 41.810 88.820 46.660 ;
        RECT 89.160 41.805 89.330 46.660 ;
        RECT 91.490 45.035 91.780 49.380 ;
        RECT 91.780 43.120 92.960 43.400 ;
        RECT 91.280 42.520 92.960 43.120 ;
        RECT 91.780 42.320 92.960 42.520 ;
        RECT 81.730 39.900 86.730 40.400 ;
        RECT 81.730 39.800 82.550 39.900 ;
        RECT 80.230 38.145 80.400 38.380 ;
        RECT 80.205 38.135 80.400 38.145 ;
        RECT 73.010 36.095 75.355 36.260 ;
        RECT 76.155 36.095 78.500 36.260 ;
        RECT 73.010 35.925 78.500 36.095 ;
        RECT 73.010 35.780 75.355 35.925 ;
        RECT 76.155 35.780 78.500 35.925 ;
        RECT 80.170 33.540 80.460 38.135 ;
        RECT 82.260 33.840 82.550 39.800 ;
        RECT 84.410 38.135 84.580 38.380 ;
        RECT 84.350 33.540 84.640 38.135 ;
        RECT 86.440 33.840 86.730 39.900 ;
        RECT 87.480 39.590 88.610 40.590 ;
        RECT 88.590 38.135 88.760 38.380 ;
        RECT 88.530 33.540 88.820 38.135 ;
        RECT 90.980 36.260 91.150 40.675 ;
        RECT 91.490 36.260 91.780 40.670 ;
        RECT 93.580 40.485 93.875 49.075 ;
        RECT 95.670 45.035 95.960 49.380 ;
        RECT 98.760 47.110 100.855 47.140 ;
        RECT 98.605 46.950 100.855 47.110 ;
        RECT 97.455 46.780 100.855 46.950 ;
        RECT 95.445 42.030 95.945 43.180 ;
        RECT 97.455 42.745 97.625 46.780 ;
        RECT 98.605 46.690 100.855 46.780 ;
        RECT 98.760 46.660 100.855 46.690 ;
        RECT 97.960 42.030 98.255 46.295 ;
        RECT 100.055 42.590 100.345 46.660 ;
        RECT 100.685 42.735 100.855 46.660 ;
        RECT 103.020 44.795 103.310 49.380 ;
        RECT 103.080 44.570 103.250 44.795 ;
        RECT 105.110 43.760 105.400 49.090 ;
        RECT 107.200 44.795 107.490 49.380 ;
        RECT 107.260 44.570 107.430 44.795 ;
        RECT 109.290 43.760 109.580 49.090 ;
        RECT 111.380 44.795 111.670 49.380 ;
        RECT 113.340 47.110 115.685 47.140 ;
        RECT 113.160 46.955 115.685 47.110 ;
        RECT 116.485 46.955 118.830 47.140 ;
        RECT 113.160 46.785 118.830 46.955 ;
        RECT 113.160 46.690 115.685 46.785 ;
        RECT 113.340 46.660 115.685 46.690 ;
        RECT 116.485 46.660 118.830 46.785 ;
        RECT 111.440 44.785 111.635 44.795 ;
        RECT 111.440 44.550 111.610 44.785 ;
        RECT 103.310 43.180 104.510 43.760 ;
        RECT 105.110 43.470 109.580 43.760 ;
        RECT 102.510 43.060 104.510 43.180 ;
        RECT 102.510 42.460 106.510 43.060 ;
        RECT 107.540 42.030 108.040 43.470 ;
        RECT 95.445 41.530 108.040 42.030 ;
        RECT 113.340 41.805 113.510 46.660 ;
        RECT 113.850 41.810 114.140 46.660 ;
        RECT 93.365 39.705 94.105 40.485 ;
        RECT 93.580 36.630 93.875 39.705 ;
        RECT 90.980 36.230 93.075 36.260 ;
        RECT 90.980 36.145 93.230 36.230 ;
        RECT 94.210 36.145 94.380 39.120 ;
        RECT 90.980 35.975 94.380 36.145 ;
        RECT 90.980 35.810 93.230 35.975 ;
        RECT 90.980 35.780 93.075 35.810 ;
        RECT 95.875 33.540 96.165 37.890 ;
        RECT 97.965 33.850 98.260 41.530 ;
        RECT 98.910 40.420 100.110 40.620 ;
        RECT 98.910 39.800 100.610 40.420 ;
        RECT 98.910 39.490 100.110 39.800 ;
        RECT 100.055 33.540 100.345 37.890 ;
        RECT 102.510 36.260 102.680 40.860 ;
        RECT 103.020 36.260 103.310 41.090 ;
        RECT 105.110 36.530 105.400 41.530 ;
        RECT 107.200 36.260 107.490 41.090 ;
        RECT 107.830 36.260 108.000 40.920 ;
        RECT 115.940 40.400 116.230 46.350 ;
        RECT 118.030 41.810 118.320 46.660 ;
        RECT 118.660 41.805 118.830 46.660 ;
        RECT 120.990 45.035 121.280 49.380 ;
        RECT 121.280 43.120 122.460 43.400 ;
        RECT 120.780 42.520 122.460 43.120 ;
        RECT 121.280 42.320 122.460 42.520 ;
        RECT 111.230 39.900 116.230 40.400 ;
        RECT 111.230 39.800 112.050 39.900 ;
        RECT 109.730 38.145 109.900 38.380 ;
        RECT 109.705 38.135 109.900 38.145 ;
        RECT 102.510 36.095 104.855 36.260 ;
        RECT 105.655 36.095 108.000 36.260 ;
        RECT 102.510 35.925 108.000 36.095 ;
        RECT 102.510 35.780 104.855 35.925 ;
        RECT 105.655 35.780 108.000 35.925 ;
        RECT 109.670 33.540 109.960 38.135 ;
        RECT 111.760 33.840 112.050 39.800 ;
        RECT 113.910 38.135 114.080 38.380 ;
        RECT 113.850 33.540 114.140 38.135 ;
        RECT 115.940 33.840 116.230 39.900 ;
        RECT 116.980 39.590 118.110 40.590 ;
        RECT 118.090 38.135 118.260 38.380 ;
        RECT 118.030 33.540 118.320 38.135 ;
        RECT 120.480 36.260 120.650 40.675 ;
        RECT 120.990 36.260 121.280 40.670 ;
        RECT 123.080 40.485 123.375 49.075 ;
        RECT 125.170 45.035 125.460 49.380 ;
        RECT 128.260 47.110 130.355 47.140 ;
        RECT 128.105 46.950 130.355 47.110 ;
        RECT 126.955 46.780 130.355 46.950 ;
        RECT 124.945 42.030 125.445 43.180 ;
        RECT 126.955 42.745 127.125 46.780 ;
        RECT 128.105 46.690 130.355 46.780 ;
        RECT 128.260 46.660 130.355 46.690 ;
        RECT 127.460 42.030 127.755 46.295 ;
        RECT 129.555 42.590 129.845 46.660 ;
        RECT 130.185 42.735 130.355 46.660 ;
        RECT 132.520 44.795 132.810 49.380 ;
        RECT 132.580 44.570 132.750 44.795 ;
        RECT 134.610 43.760 134.900 49.090 ;
        RECT 136.700 44.795 136.990 49.380 ;
        RECT 136.760 44.570 136.930 44.795 ;
        RECT 138.790 43.760 139.080 49.090 ;
        RECT 140.880 44.795 141.170 49.380 ;
        RECT 142.840 47.110 145.185 47.140 ;
        RECT 142.660 46.955 145.185 47.110 ;
        RECT 145.985 46.955 148.330 47.140 ;
        RECT 142.660 46.785 148.330 46.955 ;
        RECT 142.660 46.690 145.185 46.785 ;
        RECT 142.840 46.660 145.185 46.690 ;
        RECT 145.985 46.660 148.330 46.785 ;
        RECT 140.940 44.785 141.135 44.795 ;
        RECT 140.940 44.550 141.110 44.785 ;
        RECT 132.810 43.180 134.010 43.760 ;
        RECT 134.610 43.470 139.080 43.760 ;
        RECT 132.010 43.060 134.010 43.180 ;
        RECT 132.010 42.460 136.010 43.060 ;
        RECT 137.040 42.030 137.540 43.470 ;
        RECT 124.945 41.530 137.540 42.030 ;
        RECT 142.840 41.805 143.010 46.660 ;
        RECT 143.350 41.810 143.640 46.660 ;
        RECT 122.865 39.705 123.605 40.485 ;
        RECT 123.080 36.630 123.375 39.705 ;
        RECT 120.480 36.230 122.575 36.260 ;
        RECT 120.480 36.145 122.730 36.230 ;
        RECT 123.710 36.145 123.880 39.120 ;
        RECT 120.480 35.975 123.880 36.145 ;
        RECT 120.480 35.810 122.730 35.975 ;
        RECT 120.480 35.780 122.575 35.810 ;
        RECT 125.375 33.540 125.665 37.890 ;
        RECT 127.465 33.850 127.760 41.530 ;
        RECT 128.410 40.420 129.610 40.620 ;
        RECT 128.410 39.800 130.110 40.420 ;
        RECT 128.410 39.490 129.610 39.800 ;
        RECT 129.555 33.540 129.845 37.890 ;
        RECT 132.010 36.260 132.180 40.860 ;
        RECT 132.520 36.260 132.810 41.090 ;
        RECT 134.610 36.530 134.900 41.530 ;
        RECT 136.700 36.260 136.990 41.090 ;
        RECT 137.330 36.260 137.500 40.920 ;
        RECT 145.440 40.400 145.730 46.350 ;
        RECT 147.530 41.810 147.820 46.660 ;
        RECT 148.160 41.805 148.330 46.660 ;
        RECT 150.490 45.035 150.780 49.380 ;
        RECT 150.780 43.120 151.960 43.400 ;
        RECT 150.280 42.520 151.960 43.120 ;
        RECT 150.780 42.320 151.960 42.520 ;
        RECT 140.730 39.900 145.730 40.400 ;
        RECT 140.730 39.800 141.550 39.900 ;
        RECT 139.230 38.145 139.400 38.380 ;
        RECT 139.205 38.135 139.400 38.145 ;
        RECT 132.010 36.095 134.355 36.260 ;
        RECT 135.155 36.095 137.500 36.260 ;
        RECT 132.010 35.925 137.500 36.095 ;
        RECT 132.010 35.780 134.355 35.925 ;
        RECT 135.155 35.780 137.500 35.925 ;
        RECT 139.170 33.540 139.460 38.135 ;
        RECT 141.260 33.840 141.550 39.800 ;
        RECT 143.410 38.135 143.580 38.380 ;
        RECT 143.350 33.540 143.640 38.135 ;
        RECT 145.440 33.840 145.730 39.900 ;
        RECT 146.480 39.590 147.610 40.590 ;
        RECT 147.590 38.135 147.760 38.380 ;
        RECT 147.530 33.540 147.820 38.135 ;
        RECT 149.980 36.260 150.150 40.675 ;
        RECT 150.490 36.260 150.780 40.670 ;
        RECT 152.580 40.485 152.875 49.075 ;
        RECT 154.670 45.035 154.960 49.380 ;
        RECT 157.760 47.110 159.855 47.140 ;
        RECT 157.605 46.950 159.855 47.110 ;
        RECT 156.455 46.780 159.855 46.950 ;
        RECT 154.445 42.030 154.945 43.180 ;
        RECT 156.455 42.745 156.625 46.780 ;
        RECT 157.605 46.690 159.855 46.780 ;
        RECT 157.760 46.660 159.855 46.690 ;
        RECT 156.960 42.030 157.255 46.295 ;
        RECT 159.055 42.590 159.345 46.660 ;
        RECT 159.685 42.735 159.855 46.660 ;
        RECT 162.020 44.795 162.310 49.380 ;
        RECT 162.080 44.570 162.250 44.795 ;
        RECT 164.110 43.760 164.400 49.090 ;
        RECT 166.200 44.795 166.490 49.380 ;
        RECT 166.260 44.570 166.430 44.795 ;
        RECT 168.290 43.760 168.580 49.090 ;
        RECT 170.380 44.795 170.670 49.380 ;
        RECT 172.340 47.110 174.685 47.140 ;
        RECT 172.160 46.955 174.685 47.110 ;
        RECT 175.485 46.955 177.830 47.140 ;
        RECT 172.160 46.785 177.830 46.955 ;
        RECT 172.160 46.690 174.685 46.785 ;
        RECT 172.340 46.660 174.685 46.690 ;
        RECT 175.485 46.660 177.830 46.785 ;
        RECT 170.440 44.785 170.635 44.795 ;
        RECT 170.440 44.550 170.610 44.785 ;
        RECT 162.310 43.180 163.510 43.760 ;
        RECT 164.110 43.470 168.580 43.760 ;
        RECT 161.510 43.060 163.510 43.180 ;
        RECT 161.510 42.460 165.510 43.060 ;
        RECT 166.540 42.030 167.040 43.470 ;
        RECT 154.445 41.530 167.040 42.030 ;
        RECT 172.340 41.805 172.510 46.660 ;
        RECT 172.850 41.810 173.140 46.660 ;
        RECT 152.365 39.705 153.105 40.485 ;
        RECT 152.580 36.630 152.875 39.705 ;
        RECT 149.980 36.230 152.075 36.260 ;
        RECT 149.980 36.145 152.230 36.230 ;
        RECT 153.210 36.145 153.380 39.120 ;
        RECT 149.980 35.975 153.380 36.145 ;
        RECT 149.980 35.810 152.230 35.975 ;
        RECT 149.980 35.780 152.075 35.810 ;
        RECT 154.875 33.540 155.165 37.890 ;
        RECT 156.965 33.850 157.260 41.530 ;
        RECT 157.910 40.420 159.110 40.620 ;
        RECT 157.910 39.800 159.610 40.420 ;
        RECT 157.910 39.490 159.110 39.800 ;
        RECT 159.055 33.540 159.345 37.890 ;
        RECT 161.510 36.260 161.680 40.860 ;
        RECT 162.020 36.260 162.310 41.090 ;
        RECT 164.110 36.530 164.400 41.530 ;
        RECT 166.200 36.260 166.490 41.090 ;
        RECT 166.830 36.260 167.000 40.920 ;
        RECT 174.940 40.400 175.230 46.350 ;
        RECT 177.030 41.810 177.320 46.660 ;
        RECT 177.660 41.805 177.830 46.660 ;
        RECT 170.230 39.900 175.230 40.400 ;
        RECT 170.230 39.800 171.050 39.900 ;
        RECT 168.730 38.145 168.900 38.380 ;
        RECT 168.705 38.135 168.900 38.145 ;
        RECT 161.510 36.095 163.855 36.260 ;
        RECT 164.655 36.095 167.000 36.260 ;
        RECT 161.510 35.925 167.000 36.095 ;
        RECT 161.510 35.780 163.855 35.925 ;
        RECT 164.655 35.780 167.000 35.925 ;
        RECT 168.670 33.540 168.960 38.135 ;
        RECT 170.760 33.840 171.050 39.800 ;
        RECT 172.910 38.135 173.080 38.380 ;
        RECT 172.850 33.540 173.140 38.135 ;
        RECT 174.940 33.840 175.230 39.900 ;
        RECT 175.980 39.590 177.110 40.590 ;
        RECT 177.090 38.135 177.260 38.380 ;
        RECT 177.030 33.540 177.320 38.135 ;
        RECT 6.865 33.060 9.210 33.540 ;
        RECT 10.010 33.060 12.355 33.540 ;
        RECT 20.660 33.060 23.005 33.540 ;
        RECT 24.060 33.060 26.920 33.540 ;
        RECT 27.985 33.060 30.330 33.540 ;
        RECT 36.365 33.060 38.710 33.540 ;
        RECT 39.510 33.060 41.855 33.540 ;
        RECT 50.160 33.060 52.505 33.540 ;
        RECT 53.560 33.060 56.420 33.540 ;
        RECT 57.485 33.060 59.830 33.540 ;
        RECT 65.865 33.060 68.210 33.540 ;
        RECT 69.010 33.060 71.355 33.540 ;
        RECT 79.660 33.060 82.005 33.540 ;
        RECT 83.060 33.060 85.920 33.540 ;
        RECT 86.985 33.060 89.330 33.540 ;
        RECT 95.365 33.060 97.710 33.540 ;
        RECT 98.510 33.060 100.855 33.540 ;
        RECT 109.160 33.060 111.505 33.540 ;
        RECT 112.560 33.060 115.420 33.540 ;
        RECT 116.485 33.060 118.830 33.540 ;
        RECT 124.865 33.060 127.210 33.540 ;
        RECT 128.010 33.060 130.355 33.540 ;
        RECT 138.660 33.060 141.005 33.540 ;
        RECT 142.060 33.060 144.920 33.540 ;
        RECT 145.985 33.060 148.330 33.540 ;
        RECT 154.365 33.060 156.710 33.540 ;
        RECT 157.510 33.060 159.855 33.540 ;
        RECT 168.160 33.060 170.505 33.540 ;
        RECT 171.560 33.060 174.420 33.540 ;
        RECT 175.485 33.060 177.830 33.540 ;
        RECT 179.510 31.500 180.010 51.000 ;
        RECT 0.430 31.000 180.090 31.500 ;
      LAYER mcon ;
        RECT 36.100 73.100 36.400 73.400 ;
        RECT 36.600 73.100 36.900 73.400 ;
        RECT 37.100 73.100 37.400 73.400 ;
        RECT 37.600 73.100 37.900 73.400 ;
        RECT 72.100 73.100 72.400 73.400 ;
        RECT 72.600 73.100 72.900 73.400 ;
        RECT 73.100 73.100 73.400 73.400 ;
        RECT 73.600 73.100 73.900 73.400 ;
        RECT 108.100 73.100 108.400 73.400 ;
        RECT 108.600 73.100 108.900 73.400 ;
        RECT 109.100 73.100 109.400 73.400 ;
        RECT 109.600 73.100 109.900 73.400 ;
        RECT 144.100 73.100 144.400 73.400 ;
        RECT 144.600 73.100 144.900 73.400 ;
        RECT 145.100 73.100 145.400 73.400 ;
        RECT 145.600 73.100 145.900 73.400 ;
        RECT 3.475 63.135 3.645 63.305 ;
        RECT 3.935 63.135 4.105 63.305 ;
        RECT 4.395 63.135 4.565 63.305 ;
        RECT 4.855 63.135 5.025 63.305 ;
        RECT 5.315 63.135 5.485 63.305 ;
        RECT 7.645 63.135 7.815 63.305 ;
        RECT 8.105 63.135 8.275 63.305 ;
        RECT 8.565 63.135 8.735 63.305 ;
        RECT 2.450 61.850 2.650 62.050 ;
        RECT 6.435 61.775 6.605 61.945 ;
        RECT 3.475 60.415 3.645 60.585 ;
        RECT 3.935 60.415 4.105 60.585 ;
        RECT 4.395 60.415 4.565 60.585 ;
        RECT 4.855 60.415 5.025 60.585 ;
        RECT 5.315 60.415 5.485 60.585 ;
        RECT 7.645 60.415 7.815 60.585 ;
        RECT 8.105 60.415 8.275 60.585 ;
        RECT 8.565 60.415 8.735 60.585 ;
        RECT 18.080 71.170 18.595 71.590 ;
        RECT 18.785 71.170 19.205 71.590 ;
        RECT 19.395 71.170 19.815 71.590 ;
        RECT 20.005 71.170 20.425 71.590 ;
        RECT 21.490 71.170 21.910 71.590 ;
        RECT 22.100 71.170 22.520 71.590 ;
        RECT 22.710 71.170 23.130 71.590 ;
        RECT 23.320 71.170 23.740 71.590 ;
        RECT 23.930 71.170 24.350 71.590 ;
        RECT 25.405 71.170 25.825 71.590 ;
        RECT 26.015 71.170 26.435 71.590 ;
        RECT 26.625 71.170 27.045 71.590 ;
        RECT 27.235 71.170 27.750 71.590 ;
        RECT 36.055 71.170 36.475 71.590 ;
        RECT 36.665 71.170 37.085 71.590 ;
        RECT 37.275 71.170 37.695 71.590 ;
        RECT 37.885 71.170 38.400 71.590 ;
        RECT 39.200 71.170 39.715 71.590 ;
        RECT 39.905 71.170 40.325 71.590 ;
        RECT 40.515 71.170 40.935 71.590 ;
        RECT 41.125 71.170 41.545 71.590 ;
        RECT 47.580 71.170 48.095 71.590 ;
        RECT 48.285 71.170 48.705 71.590 ;
        RECT 48.895 71.170 49.315 71.590 ;
        RECT 49.505 71.170 49.925 71.590 ;
        RECT 50.990 71.170 51.410 71.590 ;
        RECT 51.600 71.170 52.020 71.590 ;
        RECT 52.210 71.170 52.630 71.590 ;
        RECT 52.820 71.170 53.240 71.590 ;
        RECT 53.430 71.170 53.850 71.590 ;
        RECT 54.905 71.170 55.325 71.590 ;
        RECT 55.515 71.170 55.935 71.590 ;
        RECT 56.125 71.170 56.545 71.590 ;
        RECT 56.735 71.170 57.250 71.590 ;
        RECT 65.555 71.170 65.975 71.590 ;
        RECT 66.165 71.170 66.585 71.590 ;
        RECT 66.775 71.170 67.195 71.590 ;
        RECT 67.385 71.170 67.900 71.590 ;
        RECT 68.700 71.170 69.215 71.590 ;
        RECT 69.405 71.170 69.825 71.590 ;
        RECT 70.015 71.170 70.435 71.590 ;
        RECT 70.625 71.170 71.045 71.590 ;
        RECT 77.080 71.170 77.595 71.590 ;
        RECT 77.785 71.170 78.205 71.590 ;
        RECT 78.395 71.170 78.815 71.590 ;
        RECT 79.005 71.170 79.425 71.590 ;
        RECT 80.490 71.170 80.910 71.590 ;
        RECT 81.100 71.170 81.520 71.590 ;
        RECT 81.710 71.170 82.130 71.590 ;
        RECT 82.320 71.170 82.740 71.590 ;
        RECT 82.930 71.170 83.350 71.590 ;
        RECT 84.405 71.170 84.825 71.590 ;
        RECT 85.015 71.170 85.435 71.590 ;
        RECT 85.625 71.170 86.045 71.590 ;
        RECT 86.235 71.170 86.750 71.590 ;
        RECT 95.055 71.170 95.475 71.590 ;
        RECT 95.665 71.170 96.085 71.590 ;
        RECT 96.275 71.170 96.695 71.590 ;
        RECT 96.885 71.170 97.400 71.590 ;
        RECT 98.200 71.170 98.715 71.590 ;
        RECT 98.905 71.170 99.325 71.590 ;
        RECT 99.515 71.170 99.935 71.590 ;
        RECT 100.125 71.170 100.545 71.590 ;
        RECT 106.580 71.170 107.095 71.590 ;
        RECT 107.285 71.170 107.705 71.590 ;
        RECT 107.895 71.170 108.315 71.590 ;
        RECT 108.505 71.170 108.925 71.590 ;
        RECT 109.990 71.170 110.410 71.590 ;
        RECT 110.600 71.170 111.020 71.590 ;
        RECT 111.210 71.170 111.630 71.590 ;
        RECT 111.820 71.170 112.240 71.590 ;
        RECT 112.430 71.170 112.850 71.590 ;
        RECT 113.905 71.170 114.325 71.590 ;
        RECT 114.515 71.170 114.935 71.590 ;
        RECT 115.125 71.170 115.545 71.590 ;
        RECT 115.735 71.170 116.250 71.590 ;
        RECT 124.555 71.170 124.975 71.590 ;
        RECT 125.165 71.170 125.585 71.590 ;
        RECT 125.775 71.170 126.195 71.590 ;
        RECT 126.385 71.170 126.900 71.590 ;
        RECT 127.700 71.170 128.215 71.590 ;
        RECT 128.405 71.170 128.825 71.590 ;
        RECT 129.015 71.170 129.435 71.590 ;
        RECT 129.625 71.170 130.045 71.590 ;
        RECT 136.080 71.170 136.595 71.590 ;
        RECT 136.785 71.170 137.205 71.590 ;
        RECT 137.395 71.170 137.815 71.590 ;
        RECT 138.005 71.170 138.425 71.590 ;
        RECT 139.490 71.170 139.910 71.590 ;
        RECT 140.100 71.170 140.520 71.590 ;
        RECT 140.710 71.170 141.130 71.590 ;
        RECT 141.320 71.170 141.740 71.590 ;
        RECT 141.930 71.170 142.350 71.590 ;
        RECT 143.405 71.170 143.825 71.590 ;
        RECT 144.015 71.170 144.435 71.590 ;
        RECT 144.625 71.170 145.045 71.590 ;
        RECT 145.235 71.170 145.750 71.590 ;
        RECT 154.055 71.170 154.475 71.590 ;
        RECT 154.665 71.170 155.085 71.590 ;
        RECT 155.275 71.170 155.695 71.590 ;
        RECT 155.885 71.170 156.400 71.590 ;
        RECT 157.200 71.170 157.715 71.590 ;
        RECT 157.905 71.170 158.325 71.590 ;
        RECT 158.515 71.170 158.935 71.590 ;
        RECT 159.125 71.170 159.545 71.590 ;
        RECT 18.830 64.120 19.840 65.060 ;
        RECT 28.910 68.450 29.425 68.870 ;
        RECT 29.615 68.450 30.035 68.870 ;
        RECT 30.225 68.450 30.645 68.870 ;
        RECT 30.835 68.450 31.255 68.870 ;
        RECT 32.055 68.450 32.475 68.870 ;
        RECT 32.665 68.450 33.085 68.870 ;
        RECT 33.275 68.450 33.695 68.870 ;
        RECT 33.885 68.450 34.400 68.870 ;
        RECT 24.860 64.280 25.680 64.880 ;
        RECT 36.330 64.290 36.780 64.880 ;
        RECT 36.970 64.290 38.000 64.880 ;
        RECT 44.290 68.450 44.710 68.870 ;
        RECT 44.900 68.450 45.320 68.870 ;
        RECT 45.510 68.450 45.930 68.870 ;
        RECT 42.865 64.225 43.485 64.945 ;
        RECT 30.400 61.620 31.000 62.220 ;
        RECT 31.200 61.620 31.800 62.220 ;
        RECT 32.000 61.620 32.600 62.220 ;
        RECT 32.800 61.530 33.500 62.220 ;
        RECT 33.700 61.530 34.340 62.160 ;
        RECT 18.080 57.570 18.595 57.990 ;
        RECT 18.785 57.570 19.205 57.990 ;
        RECT 19.395 57.570 19.815 57.990 ;
        RECT 20.005 57.570 20.425 57.990 ;
        RECT 21.405 57.570 21.825 57.990 ;
        RECT 22.015 57.570 22.435 57.990 ;
        RECT 22.625 57.570 23.045 57.990 ;
        RECT 23.235 57.570 23.750 57.990 ;
        RECT 36.665 57.570 37.085 57.990 ;
        RECT 37.275 57.570 37.695 57.990 ;
        RECT 37.885 57.570 38.305 57.990 ;
        RECT 40.965 61.560 41.465 62.160 ;
        RECT 48.330 64.120 49.340 65.060 ;
        RECT 58.410 68.450 58.925 68.870 ;
        RECT 59.115 68.450 59.535 68.870 ;
        RECT 59.725 68.450 60.145 68.870 ;
        RECT 60.335 68.450 60.755 68.870 ;
        RECT 61.555 68.450 61.975 68.870 ;
        RECT 62.165 68.450 62.585 68.870 ;
        RECT 62.775 68.450 63.195 68.870 ;
        RECT 63.385 68.450 63.900 68.870 ;
        RECT 54.360 64.280 55.180 64.880 ;
        RECT 44.030 61.610 44.980 62.110 ;
        RECT 45.180 61.610 45.580 62.110 ;
        RECT 65.830 64.290 66.280 64.880 ;
        RECT 66.470 64.290 67.500 64.880 ;
        RECT 73.790 68.450 74.210 68.870 ;
        RECT 74.400 68.450 74.820 68.870 ;
        RECT 75.010 68.450 75.430 68.870 ;
        RECT 72.365 64.225 72.985 64.945 ;
        RECT 59.900 61.620 60.500 62.220 ;
        RECT 60.700 61.620 61.300 62.220 ;
        RECT 61.500 61.620 62.100 62.220 ;
        RECT 62.300 61.530 63.000 62.220 ;
        RECT 63.200 61.530 63.840 62.160 ;
        RECT 47.580 57.570 48.095 57.990 ;
        RECT 48.285 57.570 48.705 57.990 ;
        RECT 48.895 57.570 49.315 57.990 ;
        RECT 49.505 57.570 49.925 57.990 ;
        RECT 50.905 57.570 51.325 57.990 ;
        RECT 51.515 57.570 51.935 57.990 ;
        RECT 52.125 57.570 52.545 57.990 ;
        RECT 52.735 57.570 53.250 57.990 ;
        RECT 66.165 57.570 66.585 57.990 ;
        RECT 66.775 57.570 67.195 57.990 ;
        RECT 67.385 57.570 67.805 57.990 ;
        RECT 70.465 61.560 70.965 62.160 ;
        RECT 77.830 64.120 78.840 65.060 ;
        RECT 87.910 68.450 88.425 68.870 ;
        RECT 88.615 68.450 89.035 68.870 ;
        RECT 89.225 68.450 89.645 68.870 ;
        RECT 89.835 68.450 90.255 68.870 ;
        RECT 91.055 68.450 91.475 68.870 ;
        RECT 91.665 68.450 92.085 68.870 ;
        RECT 92.275 68.450 92.695 68.870 ;
        RECT 92.885 68.450 93.400 68.870 ;
        RECT 83.860 64.280 84.680 64.880 ;
        RECT 73.530 61.610 74.480 62.110 ;
        RECT 74.680 61.610 75.080 62.110 ;
        RECT 95.330 64.290 95.780 64.880 ;
        RECT 95.970 64.290 97.000 64.880 ;
        RECT 103.290 68.450 103.710 68.870 ;
        RECT 103.900 68.450 104.320 68.870 ;
        RECT 104.510 68.450 104.930 68.870 ;
        RECT 101.865 64.225 102.485 64.945 ;
        RECT 89.400 61.620 90.000 62.220 ;
        RECT 90.200 61.620 90.800 62.220 ;
        RECT 91.000 61.620 91.600 62.220 ;
        RECT 91.800 61.530 92.500 62.220 ;
        RECT 92.700 61.530 93.340 62.160 ;
        RECT 77.080 57.570 77.595 57.990 ;
        RECT 77.785 57.570 78.205 57.990 ;
        RECT 78.395 57.570 78.815 57.990 ;
        RECT 79.005 57.570 79.425 57.990 ;
        RECT 80.405 57.570 80.825 57.990 ;
        RECT 81.015 57.570 81.435 57.990 ;
        RECT 81.625 57.570 82.045 57.990 ;
        RECT 82.235 57.570 82.750 57.990 ;
        RECT 95.665 57.570 96.085 57.990 ;
        RECT 96.275 57.570 96.695 57.990 ;
        RECT 96.885 57.570 97.305 57.990 ;
        RECT 99.965 61.560 100.465 62.160 ;
        RECT 107.330 64.120 108.340 65.060 ;
        RECT 117.410 68.450 117.925 68.870 ;
        RECT 118.115 68.450 118.535 68.870 ;
        RECT 118.725 68.450 119.145 68.870 ;
        RECT 119.335 68.450 119.755 68.870 ;
        RECT 120.555 68.450 120.975 68.870 ;
        RECT 121.165 68.450 121.585 68.870 ;
        RECT 121.775 68.450 122.195 68.870 ;
        RECT 122.385 68.450 122.900 68.870 ;
        RECT 113.360 64.280 114.180 64.880 ;
        RECT 103.030 61.610 103.980 62.110 ;
        RECT 104.180 61.610 104.580 62.110 ;
        RECT 124.830 64.290 125.280 64.880 ;
        RECT 125.470 64.290 126.500 64.880 ;
        RECT 132.790 68.450 133.210 68.870 ;
        RECT 133.400 68.450 133.820 68.870 ;
        RECT 134.010 68.450 134.430 68.870 ;
        RECT 131.365 64.225 131.985 64.945 ;
        RECT 118.900 61.620 119.500 62.220 ;
        RECT 119.700 61.620 120.300 62.220 ;
        RECT 120.500 61.620 121.100 62.220 ;
        RECT 121.300 61.530 122.000 62.220 ;
        RECT 122.200 61.530 122.840 62.160 ;
        RECT 106.580 57.570 107.095 57.990 ;
        RECT 107.285 57.570 107.705 57.990 ;
        RECT 107.895 57.570 108.315 57.990 ;
        RECT 108.505 57.570 108.925 57.990 ;
        RECT 109.905 57.570 110.325 57.990 ;
        RECT 110.515 57.570 110.935 57.990 ;
        RECT 111.125 57.570 111.545 57.990 ;
        RECT 111.735 57.570 112.250 57.990 ;
        RECT 125.165 57.570 125.585 57.990 ;
        RECT 125.775 57.570 126.195 57.990 ;
        RECT 126.385 57.570 126.805 57.990 ;
        RECT 129.465 61.560 129.965 62.160 ;
        RECT 136.830 64.120 137.840 65.060 ;
        RECT 146.910 68.450 147.425 68.870 ;
        RECT 147.615 68.450 148.035 68.870 ;
        RECT 148.225 68.450 148.645 68.870 ;
        RECT 148.835 68.450 149.255 68.870 ;
        RECT 150.055 68.450 150.475 68.870 ;
        RECT 150.665 68.450 151.085 68.870 ;
        RECT 151.275 68.450 151.695 68.870 ;
        RECT 151.885 68.450 152.400 68.870 ;
        RECT 142.860 64.280 143.680 64.880 ;
        RECT 132.530 61.610 133.480 62.110 ;
        RECT 133.680 61.610 134.080 62.110 ;
        RECT 154.330 64.290 154.780 64.880 ;
        RECT 154.970 64.290 156.000 64.880 ;
        RECT 162.290 68.450 162.710 68.870 ;
        RECT 162.900 68.450 163.320 68.870 ;
        RECT 163.510 68.450 163.930 68.870 ;
        RECT 160.865 64.225 161.485 64.945 ;
        RECT 148.400 61.620 149.000 62.220 ;
        RECT 149.200 61.620 149.800 62.220 ;
        RECT 150.000 61.620 150.600 62.220 ;
        RECT 150.800 61.530 151.500 62.220 ;
        RECT 151.700 61.530 152.340 62.160 ;
        RECT 136.080 57.570 136.595 57.990 ;
        RECT 136.785 57.570 137.205 57.990 ;
        RECT 137.395 57.570 137.815 57.990 ;
        RECT 138.005 57.570 138.425 57.990 ;
        RECT 139.405 57.570 139.825 57.990 ;
        RECT 140.015 57.570 140.435 57.990 ;
        RECT 140.625 57.570 141.045 57.990 ;
        RECT 141.235 57.570 141.750 57.990 ;
        RECT 154.665 57.570 155.085 57.990 ;
        RECT 155.275 57.570 155.695 57.990 ;
        RECT 155.885 57.570 156.305 57.990 ;
        RECT 158.965 61.560 159.465 62.160 ;
        RECT 162.030 61.610 162.980 62.110 ;
        RECT 163.180 61.610 163.580 62.110 ;
        RECT 24.730 54.850 25.245 55.270 ;
        RECT 25.435 54.850 25.855 55.270 ;
        RECT 26.045 54.850 26.465 55.270 ;
        RECT 26.655 54.850 27.075 55.270 ;
        RECT 28.130 54.850 28.550 55.270 ;
        RECT 28.740 54.850 29.160 55.270 ;
        RECT 29.350 54.850 29.770 55.270 ;
        RECT 29.960 54.850 30.380 55.270 ;
        RECT 30.570 54.850 30.990 55.270 ;
        RECT 32.055 54.850 32.475 55.270 ;
        RECT 32.665 54.850 33.085 55.270 ;
        RECT 33.275 54.850 33.695 55.270 ;
        RECT 33.885 54.850 34.400 55.270 ;
        RECT 41.150 54.850 41.560 55.270 ;
        RECT 41.760 54.850 42.170 55.270 ;
        RECT 42.370 54.850 42.785 55.270 ;
        RECT 44.195 54.850 44.615 55.270 ;
        RECT 44.805 54.850 45.225 55.270 ;
        RECT 45.415 54.850 45.930 55.270 ;
        RECT 54.230 54.850 54.745 55.270 ;
        RECT 54.935 54.850 55.355 55.270 ;
        RECT 55.545 54.850 55.965 55.270 ;
        RECT 56.155 54.850 56.575 55.270 ;
        RECT 57.630 54.850 58.050 55.270 ;
        RECT 58.240 54.850 58.660 55.270 ;
        RECT 58.850 54.850 59.270 55.270 ;
        RECT 59.460 54.850 59.880 55.270 ;
        RECT 60.070 54.850 60.490 55.270 ;
        RECT 61.555 54.850 61.975 55.270 ;
        RECT 62.165 54.850 62.585 55.270 ;
        RECT 62.775 54.850 63.195 55.270 ;
        RECT 63.385 54.850 63.900 55.270 ;
        RECT 70.650 54.850 71.060 55.270 ;
        RECT 71.260 54.850 71.670 55.270 ;
        RECT 71.870 54.850 72.285 55.270 ;
        RECT 73.695 54.850 74.115 55.270 ;
        RECT 74.305 54.850 74.725 55.270 ;
        RECT 74.915 54.850 75.430 55.270 ;
        RECT 83.730 54.850 84.245 55.270 ;
        RECT 84.435 54.850 84.855 55.270 ;
        RECT 85.045 54.850 85.465 55.270 ;
        RECT 85.655 54.850 86.075 55.270 ;
        RECT 87.130 54.850 87.550 55.270 ;
        RECT 87.740 54.850 88.160 55.270 ;
        RECT 88.350 54.850 88.770 55.270 ;
        RECT 88.960 54.850 89.380 55.270 ;
        RECT 89.570 54.850 89.990 55.270 ;
        RECT 91.055 54.850 91.475 55.270 ;
        RECT 91.665 54.850 92.085 55.270 ;
        RECT 92.275 54.850 92.695 55.270 ;
        RECT 92.885 54.850 93.400 55.270 ;
        RECT 100.150 54.850 100.560 55.270 ;
        RECT 100.760 54.850 101.170 55.270 ;
        RECT 101.370 54.850 101.785 55.270 ;
        RECT 103.195 54.850 103.615 55.270 ;
        RECT 103.805 54.850 104.225 55.270 ;
        RECT 104.415 54.850 104.930 55.270 ;
        RECT 113.230 54.850 113.745 55.270 ;
        RECT 113.935 54.850 114.355 55.270 ;
        RECT 114.545 54.850 114.965 55.270 ;
        RECT 115.155 54.850 115.575 55.270 ;
        RECT 116.630 54.850 117.050 55.270 ;
        RECT 117.240 54.850 117.660 55.270 ;
        RECT 117.850 54.850 118.270 55.270 ;
        RECT 118.460 54.850 118.880 55.270 ;
        RECT 119.070 54.850 119.490 55.270 ;
        RECT 120.555 54.850 120.975 55.270 ;
        RECT 121.165 54.850 121.585 55.270 ;
        RECT 121.775 54.850 122.195 55.270 ;
        RECT 122.385 54.850 122.900 55.270 ;
        RECT 129.650 54.850 130.060 55.270 ;
        RECT 130.260 54.850 130.670 55.270 ;
        RECT 130.870 54.850 131.285 55.270 ;
        RECT 132.695 54.850 133.115 55.270 ;
        RECT 133.305 54.850 133.725 55.270 ;
        RECT 133.915 54.850 134.430 55.270 ;
        RECT 142.730 54.850 143.245 55.270 ;
        RECT 143.435 54.850 143.855 55.270 ;
        RECT 144.045 54.850 144.465 55.270 ;
        RECT 144.655 54.850 145.075 55.270 ;
        RECT 146.130 54.850 146.550 55.270 ;
        RECT 146.740 54.850 147.160 55.270 ;
        RECT 147.350 54.850 147.770 55.270 ;
        RECT 147.960 54.850 148.380 55.270 ;
        RECT 148.570 54.850 148.990 55.270 ;
        RECT 150.055 54.850 150.475 55.270 ;
        RECT 150.665 54.850 151.085 55.270 ;
        RECT 151.275 54.850 151.695 55.270 ;
        RECT 151.885 54.850 152.400 55.270 ;
        RECT 159.150 54.850 159.560 55.270 ;
        RECT 159.760 54.850 160.170 55.270 ;
        RECT 160.370 54.850 160.785 55.270 ;
        RECT 162.195 54.850 162.615 55.270 ;
        RECT 162.805 54.850 163.225 55.270 ;
        RECT 163.415 54.850 163.930 55.270 ;
        RECT 3.185 49.410 3.605 49.830 ;
        RECT 3.795 49.410 4.215 49.830 ;
        RECT 4.405 49.410 4.825 49.830 ;
        RECT 6.240 49.410 6.650 49.830 ;
        RECT 6.850 49.410 7.260 49.830 ;
        RECT 7.460 49.410 7.970 49.830 ;
        RECT 14.010 49.410 14.525 49.830 ;
        RECT 14.715 49.410 15.135 49.830 ;
        RECT 15.325 49.410 15.745 49.830 ;
        RECT 15.935 49.410 16.355 49.830 ;
        RECT 17.420 49.410 17.840 49.830 ;
        RECT 18.030 49.410 18.450 49.830 ;
        RECT 18.640 49.410 19.060 49.830 ;
        RECT 19.250 49.410 19.670 49.830 ;
        RECT 19.860 49.410 20.280 49.830 ;
        RECT 21.335 49.410 21.755 49.830 ;
        RECT 21.945 49.410 22.365 49.830 ;
        RECT 22.555 49.410 22.975 49.830 ;
        RECT 23.165 49.410 23.680 49.830 ;
        RECT 32.685 49.410 33.105 49.830 ;
        RECT 33.295 49.410 33.715 49.830 ;
        RECT 33.905 49.410 34.325 49.830 ;
        RECT 35.740 49.410 36.150 49.830 ;
        RECT 36.350 49.410 36.760 49.830 ;
        RECT 36.960 49.410 37.470 49.830 ;
        RECT 43.510 49.410 44.025 49.830 ;
        RECT 44.215 49.410 44.635 49.830 ;
        RECT 44.825 49.410 45.245 49.830 ;
        RECT 45.435 49.410 45.855 49.830 ;
        RECT 46.920 49.410 47.340 49.830 ;
        RECT 47.530 49.410 47.950 49.830 ;
        RECT 48.140 49.410 48.560 49.830 ;
        RECT 48.750 49.410 49.170 49.830 ;
        RECT 49.360 49.410 49.780 49.830 ;
        RECT 50.835 49.410 51.255 49.830 ;
        RECT 51.445 49.410 51.865 49.830 ;
        RECT 52.055 49.410 52.475 49.830 ;
        RECT 52.665 49.410 53.180 49.830 ;
        RECT 62.185 49.410 62.605 49.830 ;
        RECT 62.795 49.410 63.215 49.830 ;
        RECT 63.405 49.410 63.825 49.830 ;
        RECT 65.240 49.410 65.650 49.830 ;
        RECT 65.850 49.410 66.260 49.830 ;
        RECT 66.460 49.410 66.970 49.830 ;
        RECT 73.010 49.410 73.525 49.830 ;
        RECT 73.715 49.410 74.135 49.830 ;
        RECT 74.325 49.410 74.745 49.830 ;
        RECT 74.935 49.410 75.355 49.830 ;
        RECT 76.420 49.410 76.840 49.830 ;
        RECT 77.030 49.410 77.450 49.830 ;
        RECT 77.640 49.410 78.060 49.830 ;
        RECT 78.250 49.410 78.670 49.830 ;
        RECT 78.860 49.410 79.280 49.830 ;
        RECT 80.335 49.410 80.755 49.830 ;
        RECT 80.945 49.410 81.365 49.830 ;
        RECT 81.555 49.410 81.975 49.830 ;
        RECT 82.165 49.410 82.680 49.830 ;
        RECT 91.685 49.410 92.105 49.830 ;
        RECT 92.295 49.410 92.715 49.830 ;
        RECT 92.905 49.410 93.325 49.830 ;
        RECT 94.740 49.410 95.150 49.830 ;
        RECT 95.350 49.410 95.760 49.830 ;
        RECT 95.960 49.410 96.470 49.830 ;
        RECT 102.510 49.410 103.025 49.830 ;
        RECT 103.215 49.410 103.635 49.830 ;
        RECT 103.825 49.410 104.245 49.830 ;
        RECT 104.435 49.410 104.855 49.830 ;
        RECT 105.920 49.410 106.340 49.830 ;
        RECT 106.530 49.410 106.950 49.830 ;
        RECT 107.140 49.410 107.560 49.830 ;
        RECT 107.750 49.410 108.170 49.830 ;
        RECT 108.360 49.410 108.780 49.830 ;
        RECT 109.835 49.410 110.255 49.830 ;
        RECT 110.445 49.410 110.865 49.830 ;
        RECT 111.055 49.410 111.475 49.830 ;
        RECT 111.665 49.410 112.180 49.830 ;
        RECT 121.185 49.410 121.605 49.830 ;
        RECT 121.795 49.410 122.215 49.830 ;
        RECT 122.405 49.410 122.825 49.830 ;
        RECT 124.240 49.410 124.650 49.830 ;
        RECT 124.850 49.410 125.260 49.830 ;
        RECT 125.460 49.410 125.970 49.830 ;
        RECT 132.010 49.410 132.525 49.830 ;
        RECT 132.715 49.410 133.135 49.830 ;
        RECT 133.325 49.410 133.745 49.830 ;
        RECT 133.935 49.410 134.355 49.830 ;
        RECT 135.420 49.410 135.840 49.830 ;
        RECT 136.030 49.410 136.450 49.830 ;
        RECT 136.640 49.410 137.060 49.830 ;
        RECT 137.250 49.410 137.670 49.830 ;
        RECT 137.860 49.410 138.280 49.830 ;
        RECT 139.335 49.410 139.755 49.830 ;
        RECT 139.945 49.410 140.365 49.830 ;
        RECT 140.555 49.410 140.975 49.830 ;
        RECT 141.165 49.410 141.680 49.830 ;
        RECT 150.685 49.410 151.105 49.830 ;
        RECT 151.295 49.410 151.715 49.830 ;
        RECT 151.905 49.410 152.325 49.830 ;
        RECT 153.740 49.410 154.150 49.830 ;
        RECT 154.350 49.410 154.760 49.830 ;
        RECT 154.960 49.410 155.470 49.830 ;
        RECT 161.510 49.410 162.025 49.830 ;
        RECT 162.215 49.410 162.635 49.830 ;
        RECT 162.825 49.410 163.245 49.830 ;
        RECT 163.435 49.410 163.855 49.830 ;
        RECT 164.920 49.410 165.340 49.830 ;
        RECT 165.530 49.410 165.950 49.830 ;
        RECT 166.140 49.410 166.560 49.830 ;
        RECT 166.750 49.410 167.170 49.830 ;
        RECT 167.360 49.410 167.780 49.830 ;
        RECT 168.835 49.410 169.255 49.830 ;
        RECT 169.445 49.410 169.865 49.830 ;
        RECT 170.055 49.410 170.475 49.830 ;
        RECT 170.665 49.410 171.180 49.830 ;
        RECT 2.830 42.570 3.230 43.070 ;
        RECT 3.430 42.570 4.380 43.070 ;
        RECT 6.945 42.520 7.445 43.120 ;
        RECT 10.715 46.690 11.135 47.110 ;
        RECT 11.325 46.690 11.745 47.110 ;
        RECT 11.935 46.690 12.355 47.110 ;
        RECT 25.365 46.690 25.785 47.110 ;
        RECT 25.975 46.690 26.395 47.110 ;
        RECT 26.585 46.690 27.005 47.110 ;
        RECT 27.985 46.690 28.405 47.110 ;
        RECT 28.595 46.690 29.015 47.110 ;
        RECT 29.205 46.690 29.625 47.110 ;
        RECT 29.815 46.690 30.330 47.110 ;
        RECT 14.070 42.520 14.710 43.150 ;
        RECT 14.910 42.460 15.610 43.150 ;
        RECT 15.810 42.460 16.410 43.060 ;
        RECT 16.610 42.460 17.210 43.060 ;
        RECT 17.410 42.460 18.010 43.060 ;
        RECT 4.925 39.735 5.545 40.455 ;
        RECT 3.090 35.810 3.510 36.230 ;
        RECT 3.700 35.810 4.120 36.230 ;
        RECT 4.310 35.810 4.730 36.230 ;
        RECT 10.410 39.800 11.440 40.390 ;
        RECT 11.630 39.800 12.080 40.390 ;
        RECT 32.330 42.570 32.730 43.070 ;
        RECT 32.930 42.570 33.880 43.070 ;
        RECT 14.010 35.810 14.525 36.230 ;
        RECT 14.715 35.810 15.135 36.230 ;
        RECT 15.325 35.810 15.745 36.230 ;
        RECT 15.935 35.810 16.355 36.230 ;
        RECT 17.155 35.810 17.575 36.230 ;
        RECT 17.765 35.810 18.185 36.230 ;
        RECT 18.375 35.810 18.795 36.230 ;
        RECT 18.985 35.810 19.500 36.230 ;
        RECT 28.570 39.620 29.580 40.560 ;
        RECT 36.445 42.520 36.945 43.120 ;
        RECT 40.215 46.690 40.635 47.110 ;
        RECT 40.825 46.690 41.245 47.110 ;
        RECT 41.435 46.690 41.855 47.110 ;
        RECT 54.865 46.690 55.285 47.110 ;
        RECT 55.475 46.690 55.895 47.110 ;
        RECT 56.085 46.690 56.505 47.110 ;
        RECT 57.485 46.690 57.905 47.110 ;
        RECT 58.095 46.690 58.515 47.110 ;
        RECT 58.705 46.690 59.125 47.110 ;
        RECT 59.315 46.690 59.830 47.110 ;
        RECT 43.570 42.520 44.210 43.150 ;
        RECT 44.410 42.460 45.110 43.150 ;
        RECT 45.310 42.460 45.910 43.060 ;
        RECT 46.110 42.460 46.710 43.060 ;
        RECT 46.910 42.460 47.510 43.060 ;
        RECT 34.425 39.735 35.045 40.455 ;
        RECT 32.590 35.810 33.010 36.230 ;
        RECT 33.200 35.810 33.620 36.230 ;
        RECT 33.810 35.810 34.230 36.230 ;
        RECT 39.910 39.800 40.940 40.390 ;
        RECT 41.130 39.800 41.580 40.390 ;
        RECT 61.830 42.570 62.230 43.070 ;
        RECT 62.430 42.570 63.380 43.070 ;
        RECT 43.510 35.810 44.025 36.230 ;
        RECT 44.215 35.810 44.635 36.230 ;
        RECT 44.825 35.810 45.245 36.230 ;
        RECT 45.435 35.810 45.855 36.230 ;
        RECT 46.655 35.810 47.075 36.230 ;
        RECT 47.265 35.810 47.685 36.230 ;
        RECT 47.875 35.810 48.295 36.230 ;
        RECT 48.485 35.810 49.000 36.230 ;
        RECT 58.070 39.620 59.080 40.560 ;
        RECT 65.945 42.520 66.445 43.120 ;
        RECT 69.715 46.690 70.135 47.110 ;
        RECT 70.325 46.690 70.745 47.110 ;
        RECT 70.935 46.690 71.355 47.110 ;
        RECT 84.365 46.690 84.785 47.110 ;
        RECT 84.975 46.690 85.395 47.110 ;
        RECT 85.585 46.690 86.005 47.110 ;
        RECT 86.985 46.690 87.405 47.110 ;
        RECT 87.595 46.690 88.015 47.110 ;
        RECT 88.205 46.690 88.625 47.110 ;
        RECT 88.815 46.690 89.330 47.110 ;
        RECT 73.070 42.520 73.710 43.150 ;
        RECT 73.910 42.460 74.610 43.150 ;
        RECT 74.810 42.460 75.410 43.060 ;
        RECT 75.610 42.460 76.210 43.060 ;
        RECT 76.410 42.460 77.010 43.060 ;
        RECT 63.925 39.735 64.545 40.455 ;
        RECT 62.090 35.810 62.510 36.230 ;
        RECT 62.700 35.810 63.120 36.230 ;
        RECT 63.310 35.810 63.730 36.230 ;
        RECT 69.410 39.800 70.440 40.390 ;
        RECT 70.630 39.800 71.080 40.390 ;
        RECT 91.330 42.570 91.730 43.070 ;
        RECT 91.930 42.570 92.880 43.070 ;
        RECT 73.010 35.810 73.525 36.230 ;
        RECT 73.715 35.810 74.135 36.230 ;
        RECT 74.325 35.810 74.745 36.230 ;
        RECT 74.935 35.810 75.355 36.230 ;
        RECT 76.155 35.810 76.575 36.230 ;
        RECT 76.765 35.810 77.185 36.230 ;
        RECT 77.375 35.810 77.795 36.230 ;
        RECT 77.985 35.810 78.500 36.230 ;
        RECT 87.570 39.620 88.580 40.560 ;
        RECT 95.445 42.520 95.945 43.120 ;
        RECT 99.215 46.690 99.635 47.110 ;
        RECT 99.825 46.690 100.245 47.110 ;
        RECT 100.435 46.690 100.855 47.110 ;
        RECT 113.865 46.690 114.285 47.110 ;
        RECT 114.475 46.690 114.895 47.110 ;
        RECT 115.085 46.690 115.505 47.110 ;
        RECT 116.485 46.690 116.905 47.110 ;
        RECT 117.095 46.690 117.515 47.110 ;
        RECT 117.705 46.690 118.125 47.110 ;
        RECT 118.315 46.690 118.830 47.110 ;
        RECT 102.570 42.520 103.210 43.150 ;
        RECT 103.410 42.460 104.110 43.150 ;
        RECT 104.310 42.460 104.910 43.060 ;
        RECT 105.110 42.460 105.710 43.060 ;
        RECT 105.910 42.460 106.510 43.060 ;
        RECT 93.425 39.735 94.045 40.455 ;
        RECT 91.590 35.810 92.010 36.230 ;
        RECT 92.200 35.810 92.620 36.230 ;
        RECT 92.810 35.810 93.230 36.230 ;
        RECT 98.910 39.800 99.940 40.390 ;
        RECT 100.130 39.800 100.580 40.390 ;
        RECT 120.830 42.570 121.230 43.070 ;
        RECT 121.430 42.570 122.380 43.070 ;
        RECT 102.510 35.810 103.025 36.230 ;
        RECT 103.215 35.810 103.635 36.230 ;
        RECT 103.825 35.810 104.245 36.230 ;
        RECT 104.435 35.810 104.855 36.230 ;
        RECT 105.655 35.810 106.075 36.230 ;
        RECT 106.265 35.810 106.685 36.230 ;
        RECT 106.875 35.810 107.295 36.230 ;
        RECT 107.485 35.810 108.000 36.230 ;
        RECT 117.070 39.620 118.080 40.560 ;
        RECT 124.945 42.520 125.445 43.120 ;
        RECT 128.715 46.690 129.135 47.110 ;
        RECT 129.325 46.690 129.745 47.110 ;
        RECT 129.935 46.690 130.355 47.110 ;
        RECT 143.365 46.690 143.785 47.110 ;
        RECT 143.975 46.690 144.395 47.110 ;
        RECT 144.585 46.690 145.005 47.110 ;
        RECT 145.985 46.690 146.405 47.110 ;
        RECT 146.595 46.690 147.015 47.110 ;
        RECT 147.205 46.690 147.625 47.110 ;
        RECT 147.815 46.690 148.330 47.110 ;
        RECT 132.070 42.520 132.710 43.150 ;
        RECT 132.910 42.460 133.610 43.150 ;
        RECT 133.810 42.460 134.410 43.060 ;
        RECT 134.610 42.460 135.210 43.060 ;
        RECT 135.410 42.460 136.010 43.060 ;
        RECT 122.925 39.735 123.545 40.455 ;
        RECT 121.090 35.810 121.510 36.230 ;
        RECT 121.700 35.810 122.120 36.230 ;
        RECT 122.310 35.810 122.730 36.230 ;
        RECT 128.410 39.800 129.440 40.390 ;
        RECT 129.630 39.800 130.080 40.390 ;
        RECT 150.330 42.570 150.730 43.070 ;
        RECT 150.930 42.570 151.880 43.070 ;
        RECT 132.010 35.810 132.525 36.230 ;
        RECT 132.715 35.810 133.135 36.230 ;
        RECT 133.325 35.810 133.745 36.230 ;
        RECT 133.935 35.810 134.355 36.230 ;
        RECT 135.155 35.810 135.575 36.230 ;
        RECT 135.765 35.810 136.185 36.230 ;
        RECT 136.375 35.810 136.795 36.230 ;
        RECT 136.985 35.810 137.500 36.230 ;
        RECT 146.570 39.620 147.580 40.560 ;
        RECT 154.445 42.520 154.945 43.120 ;
        RECT 158.215 46.690 158.635 47.110 ;
        RECT 158.825 46.690 159.245 47.110 ;
        RECT 159.435 46.690 159.855 47.110 ;
        RECT 172.865 46.690 173.285 47.110 ;
        RECT 173.475 46.690 173.895 47.110 ;
        RECT 174.085 46.690 174.505 47.110 ;
        RECT 175.485 46.690 175.905 47.110 ;
        RECT 176.095 46.690 176.515 47.110 ;
        RECT 176.705 46.690 177.125 47.110 ;
        RECT 177.315 46.690 177.830 47.110 ;
        RECT 161.570 42.520 162.210 43.150 ;
        RECT 162.410 42.460 163.110 43.150 ;
        RECT 163.310 42.460 163.910 43.060 ;
        RECT 164.110 42.460 164.710 43.060 ;
        RECT 164.910 42.460 165.510 43.060 ;
        RECT 152.425 39.735 153.045 40.455 ;
        RECT 150.590 35.810 151.010 36.230 ;
        RECT 151.200 35.810 151.620 36.230 ;
        RECT 151.810 35.810 152.230 36.230 ;
        RECT 157.910 39.800 158.940 40.390 ;
        RECT 159.130 39.800 159.580 40.390 ;
        RECT 161.510 35.810 162.025 36.230 ;
        RECT 162.215 35.810 162.635 36.230 ;
        RECT 162.825 35.810 163.245 36.230 ;
        RECT 163.435 35.810 163.855 36.230 ;
        RECT 164.655 35.810 165.075 36.230 ;
        RECT 165.265 35.810 165.685 36.230 ;
        RECT 165.875 35.810 166.295 36.230 ;
        RECT 166.485 35.810 167.000 36.230 ;
        RECT 176.070 39.620 177.080 40.560 ;
        RECT 6.865 33.090 7.285 33.510 ;
        RECT 7.475 33.090 7.895 33.510 ;
        RECT 8.085 33.090 8.505 33.510 ;
        RECT 8.695 33.090 9.210 33.510 ;
        RECT 10.010 33.090 10.525 33.510 ;
        RECT 10.715 33.090 11.135 33.510 ;
        RECT 11.325 33.090 11.745 33.510 ;
        RECT 11.935 33.090 12.355 33.510 ;
        RECT 20.660 33.090 21.175 33.510 ;
        RECT 21.365 33.090 21.785 33.510 ;
        RECT 21.975 33.090 22.395 33.510 ;
        RECT 22.585 33.090 23.005 33.510 ;
        RECT 24.060 33.090 24.480 33.510 ;
        RECT 24.670 33.090 25.090 33.510 ;
        RECT 25.280 33.090 25.700 33.510 ;
        RECT 25.890 33.090 26.310 33.510 ;
        RECT 26.500 33.090 26.920 33.510 ;
        RECT 27.985 33.090 28.405 33.510 ;
        RECT 28.595 33.090 29.015 33.510 ;
        RECT 29.205 33.090 29.625 33.510 ;
        RECT 29.815 33.090 30.330 33.510 ;
        RECT 36.365 33.090 36.785 33.510 ;
        RECT 36.975 33.090 37.395 33.510 ;
        RECT 37.585 33.090 38.005 33.510 ;
        RECT 38.195 33.090 38.710 33.510 ;
        RECT 39.510 33.090 40.025 33.510 ;
        RECT 40.215 33.090 40.635 33.510 ;
        RECT 40.825 33.090 41.245 33.510 ;
        RECT 41.435 33.090 41.855 33.510 ;
        RECT 50.160 33.090 50.675 33.510 ;
        RECT 50.865 33.090 51.285 33.510 ;
        RECT 51.475 33.090 51.895 33.510 ;
        RECT 52.085 33.090 52.505 33.510 ;
        RECT 53.560 33.090 53.980 33.510 ;
        RECT 54.170 33.090 54.590 33.510 ;
        RECT 54.780 33.090 55.200 33.510 ;
        RECT 55.390 33.090 55.810 33.510 ;
        RECT 56.000 33.090 56.420 33.510 ;
        RECT 57.485 33.090 57.905 33.510 ;
        RECT 58.095 33.090 58.515 33.510 ;
        RECT 58.705 33.090 59.125 33.510 ;
        RECT 59.315 33.090 59.830 33.510 ;
        RECT 65.865 33.090 66.285 33.510 ;
        RECT 66.475 33.090 66.895 33.510 ;
        RECT 67.085 33.090 67.505 33.510 ;
        RECT 67.695 33.090 68.210 33.510 ;
        RECT 69.010 33.090 69.525 33.510 ;
        RECT 69.715 33.090 70.135 33.510 ;
        RECT 70.325 33.090 70.745 33.510 ;
        RECT 70.935 33.090 71.355 33.510 ;
        RECT 79.660 33.090 80.175 33.510 ;
        RECT 80.365 33.090 80.785 33.510 ;
        RECT 80.975 33.090 81.395 33.510 ;
        RECT 81.585 33.090 82.005 33.510 ;
        RECT 83.060 33.090 83.480 33.510 ;
        RECT 83.670 33.090 84.090 33.510 ;
        RECT 84.280 33.090 84.700 33.510 ;
        RECT 84.890 33.090 85.310 33.510 ;
        RECT 85.500 33.090 85.920 33.510 ;
        RECT 86.985 33.090 87.405 33.510 ;
        RECT 87.595 33.090 88.015 33.510 ;
        RECT 88.205 33.090 88.625 33.510 ;
        RECT 88.815 33.090 89.330 33.510 ;
        RECT 95.365 33.090 95.785 33.510 ;
        RECT 95.975 33.090 96.395 33.510 ;
        RECT 96.585 33.090 97.005 33.510 ;
        RECT 97.195 33.090 97.710 33.510 ;
        RECT 98.510 33.090 99.025 33.510 ;
        RECT 99.215 33.090 99.635 33.510 ;
        RECT 99.825 33.090 100.245 33.510 ;
        RECT 100.435 33.090 100.855 33.510 ;
        RECT 109.160 33.090 109.675 33.510 ;
        RECT 109.865 33.090 110.285 33.510 ;
        RECT 110.475 33.090 110.895 33.510 ;
        RECT 111.085 33.090 111.505 33.510 ;
        RECT 112.560 33.090 112.980 33.510 ;
        RECT 113.170 33.090 113.590 33.510 ;
        RECT 113.780 33.090 114.200 33.510 ;
        RECT 114.390 33.090 114.810 33.510 ;
        RECT 115.000 33.090 115.420 33.510 ;
        RECT 116.485 33.090 116.905 33.510 ;
        RECT 117.095 33.090 117.515 33.510 ;
        RECT 117.705 33.090 118.125 33.510 ;
        RECT 118.315 33.090 118.830 33.510 ;
        RECT 124.865 33.090 125.285 33.510 ;
        RECT 125.475 33.090 125.895 33.510 ;
        RECT 126.085 33.090 126.505 33.510 ;
        RECT 126.695 33.090 127.210 33.510 ;
        RECT 128.010 33.090 128.525 33.510 ;
        RECT 128.715 33.090 129.135 33.510 ;
        RECT 129.325 33.090 129.745 33.510 ;
        RECT 129.935 33.090 130.355 33.510 ;
        RECT 138.660 33.090 139.175 33.510 ;
        RECT 139.365 33.090 139.785 33.510 ;
        RECT 139.975 33.090 140.395 33.510 ;
        RECT 140.585 33.090 141.005 33.510 ;
        RECT 142.060 33.090 142.480 33.510 ;
        RECT 142.670 33.090 143.090 33.510 ;
        RECT 143.280 33.090 143.700 33.510 ;
        RECT 143.890 33.090 144.310 33.510 ;
        RECT 144.500 33.090 144.920 33.510 ;
        RECT 145.985 33.090 146.405 33.510 ;
        RECT 146.595 33.090 147.015 33.510 ;
        RECT 147.205 33.090 147.625 33.510 ;
        RECT 147.815 33.090 148.330 33.510 ;
        RECT 154.365 33.090 154.785 33.510 ;
        RECT 154.975 33.090 155.395 33.510 ;
        RECT 155.585 33.090 156.005 33.510 ;
        RECT 156.195 33.090 156.710 33.510 ;
        RECT 157.510 33.090 158.025 33.510 ;
        RECT 158.215 33.090 158.635 33.510 ;
        RECT 158.825 33.090 159.245 33.510 ;
        RECT 159.435 33.090 159.855 33.510 ;
        RECT 168.160 33.090 168.675 33.510 ;
        RECT 168.865 33.090 169.285 33.510 ;
        RECT 169.475 33.090 169.895 33.510 ;
        RECT 170.085 33.090 170.505 33.510 ;
        RECT 171.560 33.090 171.980 33.510 ;
        RECT 172.170 33.090 172.590 33.510 ;
        RECT 172.780 33.090 173.200 33.510 ;
        RECT 173.390 33.090 173.810 33.510 ;
        RECT 174.000 33.090 174.420 33.510 ;
        RECT 175.485 33.090 175.905 33.510 ;
        RECT 176.095 33.090 176.515 33.510 ;
        RECT 176.705 33.090 177.125 33.510 ;
        RECT 177.315 33.090 177.830 33.510 ;
        RECT 36.100 31.100 36.400 31.400 ;
        RECT 36.600 31.100 36.900 31.400 ;
        RECT 37.100 31.100 37.400 31.400 ;
        RECT 37.600 31.100 37.900 31.400 ;
        RECT 72.100 31.100 72.400 31.400 ;
        RECT 72.600 31.100 72.900 31.400 ;
        RECT 73.100 31.100 73.400 31.400 ;
        RECT 73.600 31.100 73.900 31.400 ;
        RECT 108.100 31.100 108.400 31.400 ;
        RECT 108.600 31.100 108.900 31.400 ;
        RECT 109.100 31.100 109.400 31.400 ;
        RECT 109.600 31.100 109.900 31.400 ;
        RECT 144.100 31.100 144.400 31.400 ;
        RECT 144.600 31.100 144.900 31.400 ;
        RECT 145.100 31.100 145.400 31.400 ;
        RECT 145.600 31.100 145.900 31.400 ;
      LAYER met1 ;
        RECT 36.000 73.000 38.000 73.500 ;
        RECT 72.000 73.000 74.000 73.500 ;
        RECT 108.000 73.000 110.000 73.500 ;
        RECT 144.000 73.000 146.000 73.500 ;
        RECT 15.790 71.140 173.000 71.620 ;
        RECT 15.510 68.420 164.900 68.900 ;
        RECT 18.800 64.915 19.930 65.140 ;
        RECT 42.805 64.915 43.545 64.975 ;
        RECT 48.300 64.915 49.430 65.140 ;
        RECT 72.305 64.915 73.045 64.975 ;
        RECT 77.800 64.915 78.930 65.140 ;
        RECT 101.805 64.915 102.545 64.975 ;
        RECT 107.300 64.915 108.430 65.140 ;
        RECT 131.305 64.915 132.045 64.975 ;
        RECT 136.800 64.915 137.930 65.140 ;
        RECT 160.805 64.915 161.545 64.975 ;
        RECT 17.350 64.255 19.930 64.915 ;
        RECT 34.570 64.910 49.430 64.915 ;
        RECT 64.070 64.910 78.930 64.915 ;
        RECT 93.570 64.910 108.430 64.915 ;
        RECT 123.070 64.910 137.930 64.915 ;
        RECT 152.570 64.910 164.950 64.915 ;
        RECT 18.800 64.040 19.930 64.255 ;
        RECT 24.800 64.255 49.430 64.910 ;
        RECT 24.800 64.250 38.060 64.255 ;
        RECT 42.805 64.195 43.545 64.255 ;
        RECT 48.300 64.040 49.430 64.255 ;
        RECT 54.300 64.255 78.930 64.910 ;
        RECT 54.300 64.250 67.560 64.255 ;
        RECT 72.305 64.195 73.045 64.255 ;
        RECT 77.800 64.040 78.930 64.255 ;
        RECT 83.800 64.255 108.430 64.910 ;
        RECT 83.800 64.250 97.060 64.255 ;
        RECT 101.805 64.195 102.545 64.255 ;
        RECT 107.300 64.040 108.430 64.255 ;
        RECT 113.300 64.255 137.930 64.910 ;
        RECT 113.300 64.250 126.560 64.255 ;
        RECT 131.305 64.195 132.045 64.255 ;
        RECT 136.800 64.040 137.930 64.255 ;
        RECT 142.800 64.255 164.950 64.910 ;
        RECT 142.800 64.250 156.060 64.255 ;
        RECT 160.805 64.195 161.545 64.255 ;
        RECT 3.330 62.980 20.000 63.460 ;
        RECT 30.300 62.220 33.600 62.250 ;
        RECT 59.800 62.220 63.100 62.250 ;
        RECT 89.300 62.220 92.600 62.250 ;
        RECT 118.800 62.220 122.100 62.250 ;
        RECT 148.300 62.220 151.600 62.250 ;
        RECT 30.300 62.160 34.400 62.220 ;
        RECT 2.390 61.790 2.710 62.110 ;
        RECT 6.310 62.010 6.730 62.040 ;
        RECT 16.510 62.010 34.400 62.160 ;
        RECT 6.310 61.710 34.400 62.010 ;
        RECT 6.310 61.680 6.730 61.710 ;
        RECT 16.510 61.560 34.400 61.710 ;
        RECT 30.300 61.500 34.400 61.560 ;
        RECT 40.935 62.160 41.495 62.220 ;
        RECT 59.800 62.160 63.900 62.220 ;
        RECT 40.935 61.560 63.900 62.160 ;
        RECT 40.935 61.500 41.495 61.560 ;
        RECT 59.800 61.500 63.900 61.560 ;
        RECT 70.435 62.160 70.995 62.220 ;
        RECT 89.300 62.160 93.400 62.220 ;
        RECT 70.435 61.560 93.400 62.160 ;
        RECT 70.435 61.500 70.995 61.560 ;
        RECT 89.300 61.500 93.400 61.560 ;
        RECT 99.935 62.160 100.495 62.220 ;
        RECT 118.800 62.160 122.900 62.220 ;
        RECT 99.935 61.560 122.900 62.160 ;
        RECT 99.935 61.500 100.495 61.560 ;
        RECT 118.800 61.500 122.900 61.560 ;
        RECT 129.435 62.160 129.995 62.220 ;
        RECT 148.300 62.160 152.400 62.220 ;
        RECT 129.435 61.560 152.400 62.160 ;
        RECT 129.435 61.500 129.995 61.560 ;
        RECT 148.300 61.500 152.400 61.560 ;
        RECT 158.935 62.160 159.495 62.220 ;
        RECT 158.935 61.560 164.950 62.160 ;
        RECT 158.935 61.500 159.495 61.560 ;
        RECT 0.000 60.260 9.475 60.740 ;
        RECT 14.515 57.540 171.950 58.020 ;
        RECT 162.000 57.535 164.000 57.540 ;
        RECT 17.400 55.290 164.900 55.300 ;
        RECT 16.510 54.810 177.040 55.290 ;
        RECT 1.510 49.380 179.950 49.860 ;
        RECT 0.000 46.660 178.955 47.140 ;
        RECT 6.915 43.120 7.475 43.180 ;
        RECT 1.510 42.520 7.475 43.120 ;
        RECT 6.915 42.460 7.475 42.520 ;
        RECT 14.010 43.120 18.110 43.180 ;
        RECT 36.415 43.120 36.975 43.180 ;
        RECT 14.010 42.520 36.975 43.120 ;
        RECT 14.010 42.460 18.110 42.520 ;
        RECT 36.415 42.460 36.975 42.520 ;
        RECT 43.510 43.120 47.610 43.180 ;
        RECT 65.915 43.120 66.475 43.180 ;
        RECT 43.510 42.520 66.475 43.120 ;
        RECT 43.510 42.460 47.610 42.520 ;
        RECT 65.915 42.460 66.475 42.520 ;
        RECT 73.010 43.120 77.110 43.180 ;
        RECT 95.415 43.120 95.975 43.180 ;
        RECT 73.010 42.520 95.975 43.120 ;
        RECT 73.010 42.460 77.110 42.520 ;
        RECT 95.415 42.460 95.975 42.520 ;
        RECT 102.510 43.120 106.610 43.180 ;
        RECT 124.915 43.120 125.475 43.180 ;
        RECT 102.510 42.520 125.475 43.120 ;
        RECT 102.510 42.460 106.610 42.520 ;
        RECT 124.915 42.460 125.475 42.520 ;
        RECT 132.010 43.120 136.110 43.180 ;
        RECT 154.415 43.120 154.975 43.180 ;
        RECT 132.010 42.520 154.975 43.120 ;
        RECT 132.010 42.460 136.110 42.520 ;
        RECT 154.415 42.460 154.975 42.520 ;
        RECT 161.510 43.120 165.610 43.180 ;
        RECT 161.510 42.520 178.510 43.120 ;
        RECT 161.510 42.460 165.610 42.520 ;
        RECT 14.810 42.430 18.110 42.460 ;
        RECT 44.310 42.430 47.610 42.460 ;
        RECT 73.810 42.430 77.110 42.460 ;
        RECT 103.310 42.430 106.610 42.460 ;
        RECT 132.810 42.430 136.110 42.460 ;
        RECT 162.310 42.430 165.610 42.460 ;
        RECT 4.865 40.425 5.605 40.485 ;
        RECT 10.350 40.425 23.610 40.430 ;
        RECT 1.510 39.770 23.610 40.425 ;
        RECT 28.480 40.425 29.610 40.640 ;
        RECT 34.365 40.425 35.105 40.485 ;
        RECT 39.850 40.425 53.110 40.430 ;
        RECT 28.480 39.770 53.110 40.425 ;
        RECT 57.980 40.425 59.110 40.640 ;
        RECT 63.865 40.425 64.605 40.485 ;
        RECT 69.350 40.425 82.610 40.430 ;
        RECT 57.980 39.770 82.610 40.425 ;
        RECT 87.480 40.425 88.610 40.640 ;
        RECT 93.365 40.425 94.105 40.485 ;
        RECT 98.850 40.425 112.110 40.430 ;
        RECT 87.480 39.770 112.110 40.425 ;
        RECT 116.980 40.425 118.110 40.640 ;
        RECT 122.865 40.425 123.605 40.485 ;
        RECT 128.350 40.425 141.610 40.430 ;
        RECT 116.980 39.770 141.610 40.425 ;
        RECT 146.480 40.425 147.610 40.640 ;
        RECT 152.365 40.425 153.105 40.485 ;
        RECT 157.850 40.425 171.110 40.430 ;
        RECT 146.480 39.770 171.110 40.425 ;
        RECT 175.980 40.425 177.110 40.640 ;
        RECT 175.980 40.395 178.510 40.425 ;
        RECT 172.150 39.795 178.510 40.395 ;
        RECT 1.510 39.765 13.840 39.770 ;
        RECT 28.480 39.765 43.340 39.770 ;
        RECT 57.980 39.765 72.840 39.770 ;
        RECT 87.480 39.765 102.340 39.770 ;
        RECT 116.980 39.765 131.840 39.770 ;
        RECT 146.480 39.765 161.340 39.770 ;
        RECT 175.980 39.765 178.510 39.795 ;
        RECT 4.865 39.705 5.605 39.765 ;
        RECT 28.480 39.540 29.610 39.765 ;
        RECT 34.365 39.705 35.105 39.765 ;
        RECT 57.980 39.540 59.110 39.765 ;
        RECT 63.865 39.705 64.605 39.765 ;
        RECT 87.480 39.540 88.610 39.765 ;
        RECT 93.365 39.705 94.105 39.765 ;
        RECT 116.980 39.540 118.110 39.765 ;
        RECT 122.865 39.705 123.605 39.765 ;
        RECT 146.480 39.540 147.610 39.765 ;
        RECT 152.365 39.705 153.105 39.765 ;
        RECT 175.980 39.540 177.110 39.765 ;
        RECT 0.000 35.780 178.950 36.260 ;
        RECT 1.510 33.060 179.950 33.540 ;
        RECT 36.000 31.000 38.000 31.500 ;
        RECT 72.000 31.000 74.000 31.500 ;
        RECT 108.000 31.000 110.000 31.500 ;
        RECT 144.000 31.000 146.000 31.500 ;
      LAYER via ;
        RECT 36.130 73.100 36.430 73.400 ;
        RECT 36.490 73.100 36.790 73.400 ;
        RECT 36.850 73.100 37.150 73.400 ;
        RECT 37.210 73.100 37.510 73.400 ;
        RECT 37.570 73.100 37.870 73.400 ;
        RECT 72.130 73.100 72.430 73.400 ;
        RECT 72.490 73.100 72.790 73.400 ;
        RECT 72.850 73.100 73.150 73.400 ;
        RECT 73.210 73.100 73.510 73.400 ;
        RECT 73.570 73.100 73.870 73.400 ;
        RECT 108.130 73.100 108.430 73.400 ;
        RECT 108.490 73.100 108.790 73.400 ;
        RECT 108.850 73.100 109.150 73.400 ;
        RECT 109.210 73.100 109.510 73.400 ;
        RECT 109.570 73.100 109.870 73.400 ;
        RECT 144.130 73.100 144.430 73.400 ;
        RECT 144.490 73.100 144.790 73.400 ;
        RECT 144.850 73.100 145.150 73.400 ;
        RECT 145.210 73.100 145.510 73.400 ;
        RECT 145.570 73.100 145.870 73.400 ;
        RECT 38.510 71.240 38.770 71.500 ;
        RECT 38.880 71.240 39.140 71.500 ;
        RECT 39.250 71.240 39.510 71.500 ;
        RECT 69.510 71.240 69.770 71.500 ;
        RECT 69.880 71.240 70.140 71.500 ;
        RECT 70.250 71.240 70.510 71.500 ;
        RECT 111.510 71.240 111.770 71.500 ;
        RECT 111.880 71.240 112.140 71.500 ;
        RECT 112.250 71.240 112.510 71.500 ;
        RECT 142.510 71.240 142.770 71.500 ;
        RECT 142.880 71.240 143.140 71.500 ;
        RECT 143.250 71.240 143.510 71.500 ;
        RECT 172.000 71.250 172.260 71.510 ;
        RECT 172.320 71.250 172.580 71.510 ;
        RECT 172.640 71.250 172.900 71.510 ;
        RECT 18.130 68.510 18.430 68.810 ;
        RECT 18.490 68.510 18.790 68.810 ;
        RECT 18.850 68.510 19.150 68.810 ;
        RECT 19.210 68.510 19.510 68.810 ;
        RECT 19.570 68.510 19.870 68.810 ;
        RECT 54.130 68.510 54.430 68.810 ;
        RECT 54.490 68.510 54.790 68.810 ;
        RECT 54.850 68.510 55.150 68.810 ;
        RECT 55.210 68.510 55.510 68.810 ;
        RECT 55.570 68.510 55.870 68.810 ;
        RECT 90.130 68.510 90.430 68.810 ;
        RECT 90.490 68.510 90.790 68.810 ;
        RECT 90.850 68.510 91.150 68.810 ;
        RECT 91.210 68.510 91.510 68.810 ;
        RECT 91.570 68.510 91.870 68.810 ;
        RECT 126.130 68.510 126.430 68.810 ;
        RECT 126.490 68.510 126.790 68.810 ;
        RECT 126.850 68.510 127.150 68.810 ;
        RECT 127.210 68.510 127.510 68.810 ;
        RECT 127.570 68.510 127.870 68.810 ;
        RECT 162.130 68.510 162.430 68.810 ;
        RECT 162.490 68.510 162.790 68.810 ;
        RECT 162.850 68.510 163.150 68.810 ;
        RECT 163.210 68.510 163.510 68.810 ;
        RECT 163.570 68.510 163.870 68.810 ;
        RECT 17.555 64.295 18.135 64.875 ;
        RECT 163.990 64.295 164.890 64.875 ;
        RECT 18.130 63.070 18.430 63.370 ;
        RECT 18.490 63.070 18.790 63.370 ;
        RECT 18.850 63.070 19.150 63.370 ;
        RECT 19.210 63.070 19.510 63.370 ;
        RECT 19.570 63.070 19.870 63.370 ;
        RECT 2.420 61.820 2.680 62.080 ;
        RECT 17.435 61.570 18.335 62.150 ;
        RECT 46.750 61.710 47.070 62.030 ;
        RECT 47.230 61.710 47.550 62.030 ;
        RECT 75.730 61.690 76.050 62.010 ;
        RECT 76.210 61.690 76.530 62.010 ;
        RECT 105.170 61.700 105.490 62.020 ;
        RECT 105.650 61.700 105.970 62.020 ;
        RECT 135.070 61.690 135.390 62.010 ;
        RECT 135.550 61.690 135.870 62.010 ;
        RECT 163.980 61.570 164.880 62.150 ;
        RECT 0.130 60.350 0.430 60.650 ;
        RECT 0.490 60.350 0.790 60.650 ;
        RECT 0.850 60.350 1.150 60.650 ;
        RECT 1.210 60.350 1.510 60.650 ;
        RECT 1.570 60.350 1.870 60.650 ;
        RECT 18.130 57.630 18.430 57.930 ;
        RECT 18.490 57.630 18.790 57.930 ;
        RECT 18.850 57.630 19.150 57.930 ;
        RECT 19.210 57.630 19.510 57.930 ;
        RECT 19.570 57.630 19.870 57.930 ;
        RECT 54.130 57.630 54.430 57.930 ;
        RECT 54.490 57.630 54.790 57.930 ;
        RECT 54.850 57.630 55.150 57.930 ;
        RECT 55.210 57.630 55.510 57.930 ;
        RECT 55.570 57.630 55.870 57.930 ;
        RECT 90.130 57.630 90.430 57.930 ;
        RECT 90.490 57.630 90.790 57.930 ;
        RECT 90.850 57.630 91.150 57.930 ;
        RECT 91.210 57.630 91.510 57.930 ;
        RECT 91.570 57.630 91.870 57.930 ;
        RECT 126.130 57.630 126.430 57.930 ;
        RECT 126.490 57.630 126.790 57.930 ;
        RECT 126.850 57.630 127.150 57.930 ;
        RECT 127.210 57.630 127.510 57.930 ;
        RECT 127.570 57.630 127.870 57.930 ;
        RECT 162.130 57.625 162.430 57.925 ;
        RECT 162.490 57.625 162.790 57.925 ;
        RECT 162.850 57.625 163.150 57.925 ;
        RECT 163.210 57.625 163.510 57.925 ;
        RECT 163.570 57.625 163.870 57.925 ;
        RECT 38.510 54.920 38.770 55.180 ;
        RECT 38.880 54.920 39.140 55.180 ;
        RECT 39.250 54.920 39.510 55.180 ;
        RECT 69.510 54.920 69.770 55.180 ;
        RECT 69.880 54.920 70.140 55.180 ;
        RECT 70.250 54.920 70.510 55.180 ;
        RECT 111.510 54.920 111.770 55.180 ;
        RECT 111.880 54.920 112.140 55.180 ;
        RECT 112.250 54.920 112.510 55.180 ;
        RECT 142.510 54.920 142.770 55.180 ;
        RECT 142.880 54.920 143.140 55.180 ;
        RECT 143.250 54.920 143.510 55.180 ;
        RECT 172.665 54.950 172.925 55.210 ;
        RECT 173.040 54.950 173.300 55.210 ;
        RECT 173.420 54.950 173.680 55.210 ;
        RECT 173.795 54.950 174.055 55.210 ;
        RECT 174.170 54.950 174.430 55.210 ;
        RECT 174.545 54.950 174.805 55.210 ;
        RECT 174.925 54.950 175.185 55.210 ;
        RECT 175.300 54.950 175.560 55.210 ;
        RECT 175.675 54.950 175.935 55.210 ;
        RECT 176.045 54.950 176.305 55.210 ;
        RECT 176.425 54.950 176.685 55.210 ;
        RECT 38.510 49.480 38.770 49.740 ;
        RECT 38.880 49.480 39.140 49.740 ;
        RECT 39.250 49.480 39.510 49.740 ;
        RECT 69.510 49.480 69.770 49.740 ;
        RECT 69.880 49.480 70.140 49.740 ;
        RECT 70.250 49.480 70.510 49.740 ;
        RECT 111.510 49.480 111.770 49.740 ;
        RECT 111.880 49.480 112.140 49.740 ;
        RECT 112.250 49.480 112.510 49.740 ;
        RECT 142.510 49.480 142.770 49.740 ;
        RECT 142.880 49.480 143.140 49.740 ;
        RECT 143.250 49.480 143.510 49.740 ;
        RECT 178.975 49.490 179.235 49.750 ;
        RECT 179.295 49.490 179.555 49.750 ;
        RECT 179.615 49.490 179.875 49.750 ;
        RECT 18.130 46.750 18.430 47.050 ;
        RECT 18.490 46.750 18.790 47.050 ;
        RECT 18.850 46.750 19.150 47.050 ;
        RECT 19.210 46.750 19.510 47.050 ;
        RECT 19.570 46.750 19.870 47.050 ;
        RECT 54.130 46.750 54.430 47.050 ;
        RECT 54.490 46.750 54.790 47.050 ;
        RECT 54.850 46.750 55.150 47.050 ;
        RECT 55.210 46.750 55.510 47.050 ;
        RECT 55.570 46.750 55.870 47.050 ;
        RECT 90.130 46.750 90.430 47.050 ;
        RECT 90.490 46.750 90.790 47.050 ;
        RECT 90.850 46.750 91.150 47.050 ;
        RECT 91.210 46.750 91.510 47.050 ;
        RECT 91.570 46.750 91.870 47.050 ;
        RECT 126.130 46.750 126.430 47.050 ;
        RECT 126.490 46.750 126.790 47.050 ;
        RECT 126.850 46.750 127.150 47.050 ;
        RECT 127.210 46.750 127.510 47.050 ;
        RECT 127.570 46.750 127.870 47.050 ;
        RECT 162.130 46.750 162.430 47.050 ;
        RECT 162.490 46.750 162.790 47.050 ;
        RECT 162.850 46.750 163.150 47.050 ;
        RECT 163.210 46.750 163.510 47.050 ;
        RECT 163.570 46.750 163.870 47.050 ;
        RECT 6.275 42.530 6.855 43.110 ;
        RECT 31.110 42.620 31.430 42.940 ;
        RECT 31.590 42.620 31.910 42.940 ;
        RECT 60.550 42.620 60.870 42.940 ;
        RECT 61.030 42.620 61.350 42.940 ;
        RECT 89.990 42.620 90.310 42.940 ;
        RECT 90.470 42.620 90.790 42.940 ;
        RECT 119.890 42.620 120.210 42.940 ;
        RECT 120.370 42.620 120.690 42.940 ;
        RECT 149.330 42.620 149.650 42.940 ;
        RECT 149.810 42.620 150.130 42.940 ;
        RECT 165.660 42.530 166.240 43.110 ;
        RECT 166.380 42.530 166.960 43.110 ;
        RECT 3.565 39.805 4.145 40.385 ;
        RECT 172.270 39.805 172.850 40.385 ;
        RECT 18.130 35.870 18.430 36.170 ;
        RECT 18.490 35.870 18.790 36.170 ;
        RECT 18.850 35.870 19.150 36.170 ;
        RECT 19.210 35.870 19.510 36.170 ;
        RECT 19.570 35.870 19.870 36.170 ;
        RECT 54.130 35.870 54.430 36.170 ;
        RECT 54.490 35.870 54.790 36.170 ;
        RECT 54.850 35.870 55.150 36.170 ;
        RECT 55.210 35.870 55.510 36.170 ;
        RECT 55.570 35.870 55.870 36.170 ;
        RECT 126.130 35.870 126.430 36.170 ;
        RECT 126.490 35.870 126.790 36.170 ;
        RECT 126.850 35.870 127.150 36.170 ;
        RECT 127.210 35.870 127.510 36.170 ;
        RECT 127.570 35.870 127.870 36.170 ;
        RECT 162.130 35.870 162.430 36.170 ;
        RECT 162.490 35.870 162.790 36.170 ;
        RECT 162.850 35.870 163.150 36.170 ;
        RECT 163.210 35.870 163.510 36.170 ;
        RECT 163.570 35.870 163.870 36.170 ;
        RECT 38.510 33.160 38.770 33.420 ;
        RECT 38.880 33.160 39.140 33.420 ;
        RECT 39.250 33.160 39.510 33.420 ;
        RECT 69.510 33.160 69.770 33.420 ;
        RECT 69.880 33.160 70.140 33.420 ;
        RECT 70.250 33.160 70.510 33.420 ;
        RECT 111.510 33.160 111.770 33.420 ;
        RECT 111.880 33.160 112.140 33.420 ;
        RECT 112.250 33.160 112.510 33.420 ;
        RECT 142.510 33.160 142.770 33.420 ;
        RECT 142.880 33.160 143.140 33.420 ;
        RECT 143.250 33.160 143.510 33.420 ;
        RECT 178.985 33.170 179.245 33.430 ;
        RECT 179.305 33.170 179.565 33.430 ;
        RECT 179.625 33.170 179.885 33.430 ;
        RECT 36.130 31.100 36.430 31.400 ;
        RECT 36.490 31.100 36.790 31.400 ;
        RECT 36.850 31.100 37.150 31.400 ;
        RECT 37.210 31.100 37.510 31.400 ;
        RECT 37.570 31.100 37.870 31.400 ;
        RECT 72.130 31.100 72.430 31.400 ;
        RECT 72.490 31.100 72.790 31.400 ;
        RECT 72.850 31.100 73.150 31.400 ;
        RECT 73.210 31.100 73.510 31.400 ;
        RECT 73.570 31.100 73.870 31.400 ;
        RECT 108.130 31.100 108.430 31.400 ;
        RECT 108.490 31.100 108.790 31.400 ;
        RECT 108.850 31.100 109.150 31.400 ;
        RECT 109.210 31.100 109.510 31.400 ;
        RECT 109.570 31.100 109.870 31.400 ;
        RECT 144.130 31.100 144.430 31.400 ;
        RECT 144.490 31.100 144.790 31.400 ;
        RECT 144.850 31.100 145.150 31.400 ;
        RECT 145.210 31.100 145.510 31.400 ;
        RECT 145.570 31.100 145.870 31.400 ;
      LAYER met2 ;
        RECT 36.000 73.000 38.000 73.500 ;
        RECT 72.000 73.000 74.000 73.500 ;
        RECT 108.000 73.000 110.000 73.500 ;
        RECT 144.000 73.000 146.000 73.500 ;
        RECT 38.510 71.170 39.510 71.570 ;
        RECT 69.510 71.170 70.510 71.570 ;
        RECT 111.510 71.170 112.510 71.570 ;
        RECT 142.510 71.170 143.510 71.570 ;
        RECT 18.000 68.420 20.000 68.900 ;
        RECT 54.000 68.420 56.000 68.900 ;
        RECT 90.000 68.420 92.000 68.900 ;
        RECT 126.000 68.420 128.000 68.900 ;
        RECT 162.000 68.420 164.000 68.900 ;
        RECT 17.400 64.935 18.295 64.965 ;
        RECT 13.930 64.235 18.295 64.935 ;
        RECT 2.370 61.760 2.730 62.140 ;
        RECT 0.000 60.260 2.000 60.740 ;
        RECT 13.930 53.350 14.630 64.235 ;
        RECT 17.400 64.205 18.295 64.235 ;
        RECT 163.980 64.935 164.900 64.965 ;
        RECT 163.980 64.235 169.000 64.935 ;
        RECT 163.980 64.205 164.900 64.235 ;
        RECT 18.000 62.980 20.000 63.460 ;
        RECT 18.000 57.540 20.000 58.020 ;
        RECT 54.000 57.540 56.000 58.020 ;
        RECT 90.000 57.540 92.000 58.020 ;
        RECT 126.000 57.540 128.000 58.020 ;
        RECT 162.000 57.535 164.000 58.020 ;
        RECT 38.510 54.850 39.510 55.250 ;
        RECT 69.510 54.850 70.510 55.250 ;
        RECT 111.510 54.850 112.510 55.250 ;
        RECT 142.510 54.850 143.510 55.250 ;
        RECT 3.510 52.650 14.630 53.350 ;
        RECT 3.510 51.835 4.210 52.650 ;
        RECT 3.505 46.265 4.210 51.835 ;
        RECT 168.300 50.935 169.000 64.235 ;
        RECT 171.950 55.540 172.950 71.670 ;
        RECT 171.950 54.740 183.010 55.540 ;
        RECT 171.950 54.540 179.950 54.740 ;
        RECT 178.950 54.000 179.945 54.540 ;
        RECT 168.300 50.235 172.910 50.935 ;
        RECT 38.510 49.410 39.510 49.810 ;
        RECT 69.510 49.410 70.510 49.810 ;
        RECT 111.510 49.410 112.510 49.810 ;
        RECT 142.510 49.410 143.510 49.810 ;
        RECT 18.000 46.660 20.000 47.140 ;
        RECT 54.000 46.660 56.000 47.140 ;
        RECT 90.000 46.660 92.000 47.140 ;
        RECT 126.000 46.660 128.000 47.140 ;
        RECT 162.000 46.660 164.000 47.140 ;
        RECT 3.505 39.715 4.205 46.265 ;
        RECT 172.210 39.745 172.910 50.235 ;
        RECT 18.000 35.780 20.000 36.260 ;
        RECT 54.000 35.780 56.000 36.260 ;
        RECT 126.000 35.780 128.000 36.260 ;
        RECT 162.000 35.780 164.000 36.260 ;
        RECT 38.510 33.090 39.510 33.490 ;
        RECT 69.510 33.090 70.510 33.490 ;
        RECT 111.510 33.090 112.510 33.490 ;
        RECT 142.510 33.090 143.510 33.490 ;
        RECT 178.950 33.010 179.950 54.000 ;
        RECT 36.000 31.000 38.000 31.500 ;
        RECT 72.000 31.000 74.000 31.500 ;
        RECT 108.000 31.000 110.000 31.500 ;
        RECT 144.000 31.000 146.000 31.500 ;
      LAYER via2 ;
        RECT 36.180 73.090 36.500 73.410 ;
        RECT 36.620 73.090 36.940 73.410 ;
        RECT 37.060 73.090 37.380 73.410 ;
        RECT 37.500 73.090 37.820 73.410 ;
        RECT 72.180 73.090 72.500 73.410 ;
        RECT 72.620 73.090 72.940 73.410 ;
        RECT 73.060 73.090 73.380 73.410 ;
        RECT 73.500 73.090 73.820 73.410 ;
        RECT 108.180 73.090 108.500 73.410 ;
        RECT 108.620 73.090 108.940 73.410 ;
        RECT 109.060 73.090 109.380 73.410 ;
        RECT 109.500 73.090 109.820 73.410 ;
        RECT 144.180 73.090 144.500 73.410 ;
        RECT 144.620 73.090 144.940 73.410 ;
        RECT 145.060 73.090 145.380 73.410 ;
        RECT 145.500 73.090 145.820 73.410 ;
        RECT 38.610 71.220 38.910 71.520 ;
        RECT 39.110 71.220 39.410 71.520 ;
        RECT 69.610 71.220 69.910 71.520 ;
        RECT 70.110 71.220 70.410 71.520 ;
        RECT 111.610 71.220 111.910 71.520 ;
        RECT 112.110 71.220 112.410 71.520 ;
        RECT 142.610 71.220 142.910 71.520 ;
        RECT 143.110 71.220 143.410 71.520 ;
        RECT 18.180 68.500 18.500 68.820 ;
        RECT 18.620 68.500 18.940 68.820 ;
        RECT 19.060 68.500 19.380 68.820 ;
        RECT 19.500 68.500 19.820 68.820 ;
        RECT 54.180 68.500 54.500 68.820 ;
        RECT 54.620 68.500 54.940 68.820 ;
        RECT 55.060 68.500 55.380 68.820 ;
        RECT 55.500 68.500 55.820 68.820 ;
        RECT 90.180 68.500 90.500 68.820 ;
        RECT 90.620 68.500 90.940 68.820 ;
        RECT 91.060 68.500 91.380 68.820 ;
        RECT 91.500 68.500 91.820 68.820 ;
        RECT 126.180 68.500 126.500 68.820 ;
        RECT 126.620 68.500 126.940 68.820 ;
        RECT 127.060 68.500 127.380 68.820 ;
        RECT 127.500 68.500 127.820 68.820 ;
        RECT 162.180 68.500 162.500 68.820 ;
        RECT 162.620 68.500 162.940 68.820 ;
        RECT 163.060 68.500 163.380 68.820 ;
        RECT 163.500 68.500 163.820 68.820 ;
        RECT 2.410 61.810 2.690 62.090 ;
        RECT 0.180 60.340 0.500 60.660 ;
        RECT 0.620 60.340 0.940 60.660 ;
        RECT 1.060 60.340 1.380 60.660 ;
        RECT 1.500 60.340 1.820 60.660 ;
        RECT 18.180 63.060 18.500 63.380 ;
        RECT 18.620 63.060 18.940 63.380 ;
        RECT 19.060 63.060 19.380 63.380 ;
        RECT 19.500 63.060 19.820 63.380 ;
        RECT 18.180 57.620 18.500 57.940 ;
        RECT 18.620 57.620 18.940 57.940 ;
        RECT 19.060 57.620 19.380 57.940 ;
        RECT 19.500 57.620 19.820 57.940 ;
        RECT 54.180 57.620 54.500 57.940 ;
        RECT 54.620 57.620 54.940 57.940 ;
        RECT 55.060 57.620 55.380 57.940 ;
        RECT 55.500 57.620 55.820 57.940 ;
        RECT 90.180 57.620 90.500 57.940 ;
        RECT 90.620 57.620 90.940 57.940 ;
        RECT 91.060 57.620 91.380 57.940 ;
        RECT 91.500 57.620 91.820 57.940 ;
        RECT 126.180 57.620 126.500 57.940 ;
        RECT 126.620 57.620 126.940 57.940 ;
        RECT 127.060 57.620 127.380 57.940 ;
        RECT 127.500 57.620 127.820 57.940 ;
        RECT 162.180 57.615 162.500 57.935 ;
        RECT 162.620 57.615 162.940 57.935 ;
        RECT 163.060 57.615 163.380 57.935 ;
        RECT 163.500 57.615 163.820 57.935 ;
        RECT 38.610 54.900 38.910 55.200 ;
        RECT 39.110 54.900 39.410 55.200 ;
        RECT 69.610 54.900 69.910 55.200 ;
        RECT 70.110 54.900 70.410 55.200 ;
        RECT 111.610 54.900 111.910 55.200 ;
        RECT 112.110 54.900 112.410 55.200 ;
        RECT 142.610 54.900 142.910 55.200 ;
        RECT 143.110 54.900 143.410 55.200 ;
        RECT 182.010 54.940 182.410 55.340 ;
        RECT 182.540 54.940 182.940 55.340 ;
        RECT 179.260 52.400 179.660 52.800 ;
        RECT 179.260 51.870 179.660 52.270 ;
        RECT 38.610 49.460 38.910 49.760 ;
        RECT 39.110 49.460 39.410 49.760 ;
        RECT 69.610 49.460 69.910 49.760 ;
        RECT 70.110 49.460 70.410 49.760 ;
        RECT 111.610 49.460 111.910 49.760 ;
        RECT 112.110 49.460 112.410 49.760 ;
        RECT 142.610 49.460 142.910 49.760 ;
        RECT 143.110 49.460 143.410 49.760 ;
        RECT 18.180 46.740 18.500 47.060 ;
        RECT 18.620 46.740 18.940 47.060 ;
        RECT 19.060 46.740 19.380 47.060 ;
        RECT 19.500 46.740 19.820 47.060 ;
        RECT 54.180 46.740 54.500 47.060 ;
        RECT 54.620 46.740 54.940 47.060 ;
        RECT 55.060 46.740 55.380 47.060 ;
        RECT 55.500 46.740 55.820 47.060 ;
        RECT 90.180 46.740 90.500 47.060 ;
        RECT 90.620 46.740 90.940 47.060 ;
        RECT 91.060 46.740 91.380 47.060 ;
        RECT 91.500 46.740 91.820 47.060 ;
        RECT 126.180 46.740 126.500 47.060 ;
        RECT 126.620 46.740 126.940 47.060 ;
        RECT 127.060 46.740 127.380 47.060 ;
        RECT 127.500 46.740 127.820 47.060 ;
        RECT 162.180 46.740 162.500 47.060 ;
        RECT 162.620 46.740 162.940 47.060 ;
        RECT 163.060 46.740 163.380 47.060 ;
        RECT 163.500 46.740 163.820 47.060 ;
        RECT 18.180 35.860 18.500 36.180 ;
        RECT 18.620 35.860 18.940 36.180 ;
        RECT 19.060 35.860 19.380 36.180 ;
        RECT 19.500 35.860 19.820 36.180 ;
        RECT 54.180 35.860 54.500 36.180 ;
        RECT 54.620 35.860 54.940 36.180 ;
        RECT 55.060 35.860 55.380 36.180 ;
        RECT 55.500 35.860 55.820 36.180 ;
        RECT 126.180 35.860 126.500 36.180 ;
        RECT 126.620 35.860 126.940 36.180 ;
        RECT 127.060 35.860 127.380 36.180 ;
        RECT 127.500 35.860 127.820 36.180 ;
        RECT 162.180 35.860 162.500 36.180 ;
        RECT 162.620 35.860 162.940 36.180 ;
        RECT 163.060 35.860 163.380 36.180 ;
        RECT 163.500 35.860 163.820 36.180 ;
        RECT 38.610 33.140 38.910 33.440 ;
        RECT 39.110 33.140 39.410 33.440 ;
        RECT 69.610 33.140 69.910 33.440 ;
        RECT 70.110 33.140 70.410 33.440 ;
        RECT 111.610 33.140 111.910 33.440 ;
        RECT 112.110 33.140 112.410 33.440 ;
        RECT 142.610 33.140 142.910 33.440 ;
        RECT 143.110 33.140 143.410 33.440 ;
        RECT 36.180 31.090 36.500 31.410 ;
        RECT 36.620 31.090 36.940 31.410 ;
        RECT 37.060 31.090 37.380 31.410 ;
        RECT 37.500 31.090 37.820 31.410 ;
        RECT 72.180 31.090 72.500 31.410 ;
        RECT 72.620 31.090 72.940 31.410 ;
        RECT 73.060 31.090 73.380 31.410 ;
        RECT 73.500 31.090 73.820 31.410 ;
        RECT 108.180 31.090 108.500 31.410 ;
        RECT 108.620 31.090 108.940 31.410 ;
        RECT 109.060 31.090 109.380 31.410 ;
        RECT 109.500 31.090 109.820 31.410 ;
        RECT 144.180 31.090 144.500 31.410 ;
        RECT 144.620 31.090 144.940 31.410 ;
        RECT 145.060 31.090 145.380 31.410 ;
        RECT 145.500 31.090 145.820 31.410 ;
      LAYER met3 ;
        RECT 5.000 103.000 177.000 105.000 ;
        RECT 0.000 99.000 182.000 101.000 ;
        RECT 36.000 73.000 38.000 73.500 ;
        RECT 72.000 73.000 74.000 73.500 ;
        RECT 108.000 73.000 110.000 73.500 ;
        RECT 144.000 73.000 146.000 73.500 ;
        RECT 18.000 68.420 20.000 68.900 ;
        RECT 54.000 68.420 56.000 68.900 ;
        RECT 90.000 68.420 92.000 68.900 ;
        RECT 126.000 68.420 128.000 68.900 ;
        RECT 162.000 68.420 164.000 68.900 ;
        RECT 18.000 62.980 20.000 63.460 ;
        RECT 0.000 60.260 2.000 60.740 ;
        RECT 18.000 57.540 20.000 58.020 ;
        RECT 54.000 57.540 56.000 58.020 ;
        RECT 90.000 57.540 92.000 58.020 ;
        RECT 126.000 57.540 128.000 58.020 ;
        RECT 162.000 57.535 164.000 58.020 ;
        RECT 18.000 46.660 20.000 47.140 ;
        RECT 54.000 46.660 56.000 47.140 ;
        RECT 90.000 46.660 92.000 47.140 ;
        RECT 126.000 46.660 128.000 47.140 ;
        RECT 162.000 46.660 164.000 47.140 ;
        RECT 18.000 35.780 20.000 36.260 ;
        RECT 54.000 35.780 56.000 36.260 ;
        RECT 126.000 35.780 128.000 36.260 ;
        RECT 162.000 35.780 164.000 36.260 ;
        RECT 36.000 31.000 38.000 31.500 ;
        RECT 72.000 31.000 74.000 31.500 ;
        RECT 108.000 31.000 110.000 31.500 ;
        RECT 144.000 31.000 146.000 31.500 ;
        RECT 0.000 4.000 182.000 6.000 ;
        RECT 5.000 0.000 177.000 2.000 ;
      LAYER via3 ;
        RECT 5.200 104.400 5.600 104.800 ;
        RECT 5.800 104.400 6.200 104.800 ;
        RECT 6.400 104.400 6.800 104.800 ;
        RECT 18.200 104.400 18.600 104.800 ;
        RECT 18.800 104.400 19.200 104.800 ;
        RECT 19.400 104.400 19.800 104.800 ;
        RECT 54.200 104.400 54.600 104.800 ;
        RECT 54.800 104.400 55.200 104.800 ;
        RECT 55.400 104.400 55.800 104.800 ;
        RECT 90.200 104.400 90.600 104.800 ;
        RECT 90.800 104.400 91.200 104.800 ;
        RECT 91.400 104.400 91.800 104.800 ;
        RECT 126.200 104.400 126.600 104.800 ;
        RECT 126.800 104.400 127.200 104.800 ;
        RECT 127.400 104.400 127.800 104.800 ;
        RECT 162.200 104.400 162.600 104.800 ;
        RECT 162.800 104.400 163.200 104.800 ;
        RECT 163.400 104.400 163.800 104.800 ;
        RECT 175.200 104.400 175.600 104.800 ;
        RECT 175.800 104.400 176.200 104.800 ;
        RECT 176.400 104.400 176.800 104.800 ;
        RECT 5.200 103.800 5.600 104.200 ;
        RECT 5.800 103.800 6.200 104.200 ;
        RECT 6.400 103.800 6.800 104.200 ;
        RECT 18.200 103.800 18.600 104.200 ;
        RECT 18.800 103.800 19.200 104.200 ;
        RECT 19.400 103.800 19.800 104.200 ;
        RECT 54.200 103.800 54.600 104.200 ;
        RECT 54.800 103.800 55.200 104.200 ;
        RECT 55.400 103.800 55.800 104.200 ;
        RECT 90.200 103.800 90.600 104.200 ;
        RECT 90.800 103.800 91.200 104.200 ;
        RECT 91.400 103.800 91.800 104.200 ;
        RECT 126.200 103.800 126.600 104.200 ;
        RECT 126.800 103.800 127.200 104.200 ;
        RECT 127.400 103.800 127.800 104.200 ;
        RECT 162.200 103.800 162.600 104.200 ;
        RECT 162.800 103.800 163.200 104.200 ;
        RECT 163.400 103.800 163.800 104.200 ;
        RECT 175.200 103.800 175.600 104.200 ;
        RECT 175.800 103.800 176.200 104.200 ;
        RECT 176.400 103.800 176.800 104.200 ;
        RECT 5.200 103.200 5.600 103.600 ;
        RECT 5.800 103.200 6.200 103.600 ;
        RECT 6.400 103.200 6.800 103.600 ;
        RECT 18.200 103.200 18.600 103.600 ;
        RECT 18.800 103.200 19.200 103.600 ;
        RECT 19.400 103.200 19.800 103.600 ;
        RECT 54.200 103.200 54.600 103.600 ;
        RECT 54.800 103.200 55.200 103.600 ;
        RECT 55.400 103.200 55.800 103.600 ;
        RECT 90.200 103.200 90.600 103.600 ;
        RECT 90.800 103.200 91.200 103.600 ;
        RECT 91.400 103.200 91.800 103.600 ;
        RECT 126.200 103.200 126.600 103.600 ;
        RECT 126.800 103.200 127.200 103.600 ;
        RECT 127.400 103.200 127.800 103.600 ;
        RECT 162.200 103.200 162.600 103.600 ;
        RECT 162.800 103.200 163.200 103.600 ;
        RECT 163.400 103.200 163.800 103.600 ;
        RECT 175.200 103.200 175.600 103.600 ;
        RECT 175.800 103.200 176.200 103.600 ;
        RECT 176.400 103.200 176.800 103.600 ;
        RECT 0.200 100.400 0.600 100.800 ;
        RECT 0.800 100.400 1.200 100.800 ;
        RECT 1.400 100.400 1.800 100.800 ;
        RECT 36.200 100.400 36.600 100.800 ;
        RECT 36.800 100.400 37.200 100.800 ;
        RECT 37.400 100.400 37.800 100.800 ;
        RECT 72.200 100.400 72.600 100.800 ;
        RECT 72.800 100.400 73.200 100.800 ;
        RECT 73.400 100.400 73.800 100.800 ;
        RECT 108.200 100.400 108.600 100.800 ;
        RECT 108.800 100.400 109.200 100.800 ;
        RECT 109.400 100.400 109.800 100.800 ;
        RECT 144.200 100.400 144.600 100.800 ;
        RECT 144.800 100.400 145.200 100.800 ;
        RECT 145.400 100.400 145.800 100.800 ;
        RECT 180.200 100.400 180.600 100.800 ;
        RECT 180.800 100.400 181.200 100.800 ;
        RECT 181.400 100.400 181.800 100.800 ;
        RECT 0.200 99.800 0.600 100.200 ;
        RECT 0.800 99.800 1.200 100.200 ;
        RECT 1.400 99.800 1.800 100.200 ;
        RECT 36.200 99.800 36.600 100.200 ;
        RECT 36.800 99.800 37.200 100.200 ;
        RECT 37.400 99.800 37.800 100.200 ;
        RECT 72.200 99.800 72.600 100.200 ;
        RECT 72.800 99.800 73.200 100.200 ;
        RECT 73.400 99.800 73.800 100.200 ;
        RECT 108.200 99.800 108.600 100.200 ;
        RECT 108.800 99.800 109.200 100.200 ;
        RECT 109.400 99.800 109.800 100.200 ;
        RECT 144.200 99.800 144.600 100.200 ;
        RECT 144.800 99.800 145.200 100.200 ;
        RECT 145.400 99.800 145.800 100.200 ;
        RECT 180.200 99.800 180.600 100.200 ;
        RECT 180.800 99.800 181.200 100.200 ;
        RECT 181.400 99.800 181.800 100.200 ;
        RECT 0.200 99.200 0.600 99.600 ;
        RECT 0.800 99.200 1.200 99.600 ;
        RECT 1.400 99.200 1.800 99.600 ;
        RECT 36.200 99.200 36.600 99.600 ;
        RECT 36.800 99.200 37.200 99.600 ;
        RECT 37.400 99.200 37.800 99.600 ;
        RECT 72.200 99.200 72.600 99.600 ;
        RECT 72.800 99.200 73.200 99.600 ;
        RECT 73.400 99.200 73.800 99.600 ;
        RECT 108.200 99.200 108.600 99.600 ;
        RECT 108.800 99.200 109.200 99.600 ;
        RECT 109.400 99.200 109.800 99.600 ;
        RECT 144.200 99.200 144.600 99.600 ;
        RECT 144.800 99.200 145.200 99.600 ;
        RECT 145.400 99.200 145.800 99.600 ;
        RECT 180.200 99.200 180.600 99.600 ;
        RECT 180.800 99.200 181.200 99.600 ;
        RECT 181.400 99.200 181.800 99.600 ;
        RECT 36.160 73.070 36.520 73.435 ;
        RECT 36.600 73.070 36.960 73.435 ;
        RECT 37.040 73.070 37.400 73.435 ;
        RECT 37.480 73.070 37.840 73.435 ;
        RECT 72.160 73.070 72.520 73.435 ;
        RECT 72.600 73.070 72.960 73.435 ;
        RECT 73.040 73.070 73.400 73.435 ;
        RECT 73.480 73.070 73.840 73.435 ;
        RECT 108.160 73.070 108.520 73.435 ;
        RECT 108.600 73.070 108.960 73.435 ;
        RECT 109.040 73.070 109.400 73.435 ;
        RECT 109.480 73.070 109.840 73.435 ;
        RECT 144.160 73.070 144.520 73.435 ;
        RECT 144.600 73.070 144.960 73.435 ;
        RECT 145.040 73.070 145.400 73.435 ;
        RECT 145.480 73.070 145.840 73.435 ;
        RECT 18.160 68.480 18.520 68.840 ;
        RECT 18.600 68.480 18.960 68.840 ;
        RECT 19.040 68.480 19.400 68.840 ;
        RECT 19.480 68.480 19.840 68.840 ;
        RECT 54.160 68.480 54.520 68.840 ;
        RECT 54.600 68.480 54.960 68.840 ;
        RECT 55.040 68.480 55.400 68.840 ;
        RECT 55.480 68.480 55.840 68.840 ;
        RECT 90.160 68.480 90.520 68.840 ;
        RECT 90.600 68.480 90.960 68.840 ;
        RECT 91.040 68.480 91.400 68.840 ;
        RECT 91.480 68.480 91.840 68.840 ;
        RECT 126.160 68.480 126.520 68.840 ;
        RECT 126.600 68.480 126.960 68.840 ;
        RECT 127.040 68.480 127.400 68.840 ;
        RECT 127.480 68.480 127.840 68.840 ;
        RECT 162.160 68.480 162.520 68.840 ;
        RECT 162.600 68.480 162.960 68.840 ;
        RECT 163.040 68.480 163.400 68.840 ;
        RECT 163.480 68.480 163.840 68.840 ;
        RECT 18.160 63.040 18.520 63.400 ;
        RECT 18.600 63.040 18.960 63.400 ;
        RECT 19.040 63.040 19.400 63.400 ;
        RECT 19.480 63.040 19.840 63.400 ;
        RECT 0.160 60.320 0.520 60.685 ;
        RECT 0.600 60.320 0.960 60.685 ;
        RECT 1.040 60.320 1.400 60.685 ;
        RECT 1.480 60.320 1.840 60.685 ;
        RECT 18.160 57.600 18.520 57.960 ;
        RECT 18.600 57.600 18.960 57.960 ;
        RECT 19.040 57.600 19.400 57.960 ;
        RECT 19.480 57.600 19.840 57.960 ;
        RECT 54.160 57.600 54.520 57.960 ;
        RECT 54.600 57.600 54.960 57.960 ;
        RECT 55.040 57.600 55.400 57.960 ;
        RECT 55.480 57.600 55.840 57.960 ;
        RECT 90.160 57.600 90.520 57.960 ;
        RECT 90.600 57.600 90.960 57.960 ;
        RECT 91.040 57.600 91.400 57.960 ;
        RECT 91.480 57.600 91.840 57.960 ;
        RECT 126.160 57.600 126.520 57.960 ;
        RECT 126.600 57.600 126.960 57.960 ;
        RECT 127.040 57.600 127.400 57.960 ;
        RECT 127.480 57.600 127.840 57.960 ;
        RECT 162.160 57.595 162.520 57.960 ;
        RECT 162.600 57.595 162.960 57.960 ;
        RECT 163.040 57.595 163.400 57.960 ;
        RECT 163.480 57.595 163.840 57.960 ;
        RECT 18.160 46.720 18.520 47.085 ;
        RECT 18.600 46.720 18.960 47.085 ;
        RECT 19.040 46.720 19.400 47.085 ;
        RECT 19.480 46.720 19.840 47.085 ;
        RECT 54.160 46.720 54.520 47.085 ;
        RECT 54.600 46.720 54.960 47.085 ;
        RECT 55.040 46.720 55.400 47.085 ;
        RECT 55.480 46.720 55.840 47.085 ;
        RECT 90.160 46.720 90.520 47.085 ;
        RECT 90.600 46.720 90.960 47.085 ;
        RECT 91.040 46.720 91.400 47.085 ;
        RECT 91.480 46.720 91.840 47.085 ;
        RECT 126.160 46.720 126.520 47.085 ;
        RECT 126.600 46.720 126.960 47.085 ;
        RECT 127.040 46.720 127.400 47.085 ;
        RECT 127.480 46.720 127.840 47.085 ;
        RECT 162.160 46.720 162.520 47.085 ;
        RECT 162.600 46.720 162.960 47.085 ;
        RECT 163.040 46.720 163.400 47.085 ;
        RECT 163.480 46.720 163.840 47.085 ;
        RECT 18.160 35.840 18.520 36.205 ;
        RECT 18.600 35.840 18.960 36.205 ;
        RECT 19.040 35.840 19.400 36.205 ;
        RECT 19.480 35.840 19.840 36.205 ;
        RECT 54.160 35.840 54.520 36.205 ;
        RECT 54.600 35.840 54.960 36.205 ;
        RECT 55.040 35.840 55.400 36.205 ;
        RECT 55.480 35.840 55.840 36.205 ;
        RECT 126.160 35.840 126.520 36.205 ;
        RECT 126.600 35.840 126.960 36.205 ;
        RECT 127.040 35.840 127.400 36.205 ;
        RECT 127.480 35.840 127.840 36.205 ;
        RECT 162.160 35.840 162.520 36.205 ;
        RECT 162.600 35.840 162.960 36.205 ;
        RECT 163.040 35.840 163.400 36.205 ;
        RECT 163.480 35.840 163.840 36.205 ;
        RECT 36.160 31.070 36.520 31.435 ;
        RECT 36.600 31.070 36.960 31.435 ;
        RECT 37.040 31.070 37.400 31.435 ;
        RECT 37.480 31.070 37.840 31.435 ;
        RECT 72.160 31.070 72.520 31.435 ;
        RECT 72.600 31.070 72.960 31.435 ;
        RECT 73.040 31.070 73.400 31.435 ;
        RECT 73.480 31.070 73.840 31.435 ;
        RECT 108.160 31.070 108.520 31.435 ;
        RECT 108.600 31.070 108.960 31.435 ;
        RECT 109.040 31.070 109.400 31.435 ;
        RECT 109.480 31.070 109.840 31.435 ;
        RECT 144.160 31.070 144.520 31.435 ;
        RECT 144.600 31.070 144.960 31.435 ;
        RECT 145.040 31.070 145.400 31.435 ;
        RECT 145.480 31.070 145.840 31.435 ;
        RECT 0.200 5.400 0.600 5.800 ;
        RECT 0.800 5.400 1.200 5.800 ;
        RECT 1.400 5.400 1.800 5.800 ;
        RECT 36.200 5.400 36.600 5.800 ;
        RECT 36.800 5.400 37.200 5.800 ;
        RECT 37.400 5.400 37.800 5.800 ;
        RECT 72.200 5.400 72.600 5.800 ;
        RECT 72.800 5.400 73.200 5.800 ;
        RECT 73.400 5.400 73.800 5.800 ;
        RECT 108.200 5.400 108.600 5.800 ;
        RECT 108.800 5.400 109.200 5.800 ;
        RECT 109.400 5.400 109.800 5.800 ;
        RECT 144.200 5.400 144.600 5.800 ;
        RECT 144.800 5.400 145.200 5.800 ;
        RECT 145.400 5.400 145.800 5.800 ;
        RECT 180.200 5.400 180.600 5.800 ;
        RECT 180.800 5.400 181.200 5.800 ;
        RECT 181.400 5.400 181.800 5.800 ;
        RECT 0.200 4.800 0.600 5.200 ;
        RECT 0.800 4.800 1.200 5.200 ;
        RECT 1.400 4.800 1.800 5.200 ;
        RECT 36.200 4.800 36.600 5.200 ;
        RECT 36.800 4.800 37.200 5.200 ;
        RECT 37.400 4.800 37.800 5.200 ;
        RECT 72.200 4.800 72.600 5.200 ;
        RECT 72.800 4.800 73.200 5.200 ;
        RECT 73.400 4.800 73.800 5.200 ;
        RECT 108.200 4.800 108.600 5.200 ;
        RECT 108.800 4.800 109.200 5.200 ;
        RECT 109.400 4.800 109.800 5.200 ;
        RECT 144.200 4.800 144.600 5.200 ;
        RECT 144.800 4.800 145.200 5.200 ;
        RECT 145.400 4.800 145.800 5.200 ;
        RECT 180.200 4.800 180.600 5.200 ;
        RECT 180.800 4.800 181.200 5.200 ;
        RECT 181.400 4.800 181.800 5.200 ;
        RECT 0.200 4.200 0.600 4.600 ;
        RECT 0.800 4.200 1.200 4.600 ;
        RECT 1.400 4.200 1.800 4.600 ;
        RECT 36.200 4.200 36.600 4.600 ;
        RECT 36.800 4.200 37.200 4.600 ;
        RECT 37.400 4.200 37.800 4.600 ;
        RECT 72.200 4.200 72.600 4.600 ;
        RECT 72.800 4.200 73.200 4.600 ;
        RECT 73.400 4.200 73.800 4.600 ;
        RECT 108.200 4.200 108.600 4.600 ;
        RECT 108.800 4.200 109.200 4.600 ;
        RECT 109.400 4.200 109.800 4.600 ;
        RECT 144.200 4.200 144.600 4.600 ;
        RECT 144.800 4.200 145.200 4.600 ;
        RECT 145.400 4.200 145.800 4.600 ;
        RECT 180.200 4.200 180.600 4.600 ;
        RECT 180.800 4.200 181.200 4.600 ;
        RECT 181.400 4.200 181.800 4.600 ;
        RECT 5.200 1.400 5.600 1.800 ;
        RECT 5.800 1.400 6.200 1.800 ;
        RECT 6.400 1.400 6.800 1.800 ;
        RECT 18.200 1.400 18.600 1.800 ;
        RECT 18.800 1.400 19.200 1.800 ;
        RECT 19.400 1.400 19.800 1.800 ;
        RECT 54.200 1.400 54.600 1.800 ;
        RECT 54.800 1.400 55.200 1.800 ;
        RECT 55.400 1.400 55.800 1.800 ;
        RECT 90.200 1.400 90.600 1.800 ;
        RECT 90.800 1.400 91.200 1.800 ;
        RECT 91.400 1.400 91.800 1.800 ;
        RECT 126.200 1.400 126.600 1.800 ;
        RECT 126.800 1.400 127.200 1.800 ;
        RECT 127.400 1.400 127.800 1.800 ;
        RECT 162.200 1.400 162.600 1.800 ;
        RECT 162.800 1.400 163.200 1.800 ;
        RECT 163.400 1.400 163.800 1.800 ;
        RECT 175.200 1.400 175.600 1.800 ;
        RECT 175.800 1.400 176.200 1.800 ;
        RECT 176.400 1.400 176.800 1.800 ;
        RECT 5.200 0.800 5.600 1.200 ;
        RECT 5.800 0.800 6.200 1.200 ;
        RECT 6.400 0.800 6.800 1.200 ;
        RECT 18.200 0.800 18.600 1.200 ;
        RECT 18.800 0.800 19.200 1.200 ;
        RECT 19.400 0.800 19.800 1.200 ;
        RECT 54.200 0.800 54.600 1.200 ;
        RECT 54.800 0.800 55.200 1.200 ;
        RECT 55.400 0.800 55.800 1.200 ;
        RECT 90.200 0.800 90.600 1.200 ;
        RECT 90.800 0.800 91.200 1.200 ;
        RECT 91.400 0.800 91.800 1.200 ;
        RECT 126.200 0.800 126.600 1.200 ;
        RECT 126.800 0.800 127.200 1.200 ;
        RECT 127.400 0.800 127.800 1.200 ;
        RECT 162.200 0.800 162.600 1.200 ;
        RECT 162.800 0.800 163.200 1.200 ;
        RECT 163.400 0.800 163.800 1.200 ;
        RECT 175.200 0.800 175.600 1.200 ;
        RECT 175.800 0.800 176.200 1.200 ;
        RECT 176.400 0.800 176.800 1.200 ;
        RECT 5.200 0.200 5.600 0.600 ;
        RECT 5.800 0.200 6.200 0.600 ;
        RECT 6.400 0.200 6.800 0.600 ;
        RECT 18.200 0.200 18.600 0.600 ;
        RECT 18.800 0.200 19.200 0.600 ;
        RECT 19.400 0.200 19.800 0.600 ;
        RECT 54.200 0.200 54.600 0.600 ;
        RECT 54.800 0.200 55.200 0.600 ;
        RECT 55.400 0.200 55.800 0.600 ;
        RECT 90.200 0.200 90.600 0.600 ;
        RECT 90.800 0.200 91.200 0.600 ;
        RECT 91.400 0.200 91.800 0.600 ;
        RECT 126.200 0.200 126.600 0.600 ;
        RECT 126.800 0.200 127.200 0.600 ;
        RECT 127.400 0.200 127.800 0.600 ;
        RECT 162.200 0.200 162.600 0.600 ;
        RECT 162.800 0.200 163.200 0.600 ;
        RECT 163.400 0.200 163.800 0.600 ;
        RECT 175.200 0.200 175.600 0.600 ;
        RECT 175.800 0.200 176.200 0.600 ;
        RECT 176.400 0.200 176.800 0.600 ;
  END
END vco
END LIBRARY

