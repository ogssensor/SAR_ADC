magic
tech sky130A
magscale 1 2
timestamp 1625495064
<< obsli1 >>
rect 1104 1785 179003 137649
<< obsm1 >>
rect 842 1572 179202 137680
<< metal2 >>
rect 1030 139200 1086 140000
rect 3146 139200 3202 140000
rect 5354 139200 5410 140000
rect 7562 139200 7618 140000
rect 9770 139200 9826 140000
rect 11978 139200 12034 140000
rect 14186 139200 14242 140000
rect 16394 139200 16450 140000
rect 18510 139200 18566 140000
rect 20718 139200 20774 140000
rect 22926 139200 22982 140000
rect 25134 139200 25190 140000
rect 27342 139200 27398 140000
rect 29550 139200 29606 140000
rect 31758 139200 31814 140000
rect 33874 139200 33930 140000
rect 36082 139200 36138 140000
rect 38290 139200 38346 140000
rect 40498 139200 40554 140000
rect 42706 139200 42762 140000
rect 44914 139200 44970 140000
rect 47122 139200 47178 140000
rect 49330 139200 49386 140000
rect 51446 139200 51502 140000
rect 53654 139200 53710 140000
rect 55862 139200 55918 140000
rect 58070 139200 58126 140000
rect 60278 139200 60334 140000
rect 62486 139200 62542 140000
rect 64694 139200 64750 140000
rect 66810 139200 66866 140000
rect 69018 139200 69074 140000
rect 71226 139200 71282 140000
rect 73434 139200 73490 140000
rect 75642 139200 75698 140000
rect 77850 139200 77906 140000
rect 80058 139200 80114 140000
rect 82266 139200 82322 140000
rect 84382 139200 84438 140000
rect 86590 139200 86646 140000
rect 88798 139200 88854 140000
rect 91006 139200 91062 140000
rect 93214 139200 93270 140000
rect 95422 139200 95478 140000
rect 97630 139200 97686 140000
rect 99746 139200 99802 140000
rect 101954 139200 102010 140000
rect 104162 139200 104218 140000
rect 106370 139200 106426 140000
rect 108578 139200 108634 140000
rect 110786 139200 110842 140000
rect 112994 139200 113050 140000
rect 115202 139200 115258 140000
rect 117318 139200 117374 140000
rect 119526 139200 119582 140000
rect 121734 139200 121790 140000
rect 123942 139200 123998 140000
rect 126150 139200 126206 140000
rect 128358 139200 128414 140000
rect 130566 139200 130622 140000
rect 132682 139200 132738 140000
rect 134890 139200 134946 140000
rect 137098 139200 137154 140000
rect 139306 139200 139362 140000
rect 141514 139200 141570 140000
rect 143722 139200 143778 140000
rect 145930 139200 145986 140000
rect 148138 139200 148194 140000
rect 150254 139200 150310 140000
rect 152462 139200 152518 140000
rect 154670 139200 154726 140000
rect 156878 139200 156934 140000
rect 159086 139200 159142 140000
rect 161294 139200 161350 140000
rect 163502 139200 163558 140000
rect 165618 139200 165674 140000
rect 167826 139200 167882 140000
rect 170034 139200 170090 140000
rect 172242 139200 172298 140000
rect 174450 139200 174506 140000
rect 176658 139200 176714 140000
rect 178866 139200 178922 140000
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5906 0 5962 800
rect 7562 0 7618 800
rect 9310 0 9366 800
rect 10966 0 11022 800
rect 12714 0 12770 800
rect 14370 0 14426 800
rect 16118 0 16174 800
rect 17774 0 17830 800
rect 19522 0 19578 800
rect 21178 0 21234 800
rect 22926 0 22982 800
rect 24582 0 24638 800
rect 26238 0 26294 800
rect 27986 0 28042 800
rect 29642 0 29698 800
rect 31390 0 31446 800
rect 33046 0 33102 800
rect 34794 0 34850 800
rect 36450 0 36506 800
rect 38198 0 38254 800
rect 39854 0 39910 800
rect 41602 0 41658 800
rect 43258 0 43314 800
rect 45006 0 45062 800
rect 46662 0 46718 800
rect 48318 0 48374 800
rect 50066 0 50122 800
rect 51722 0 51778 800
rect 53470 0 53526 800
rect 55126 0 55182 800
rect 56874 0 56930 800
rect 58530 0 58586 800
rect 60278 0 60334 800
rect 61934 0 61990 800
rect 63682 0 63738 800
rect 65338 0 65394 800
rect 67086 0 67142 800
rect 68742 0 68798 800
rect 70398 0 70454 800
rect 72146 0 72202 800
rect 73802 0 73858 800
rect 75550 0 75606 800
rect 77206 0 77262 800
rect 78954 0 79010 800
rect 80610 0 80666 800
rect 82358 0 82414 800
rect 84014 0 84070 800
rect 85762 0 85818 800
rect 87418 0 87474 800
rect 89166 0 89222 800
rect 90822 0 90878 800
rect 92478 0 92534 800
rect 94226 0 94282 800
rect 95882 0 95938 800
rect 97630 0 97686 800
rect 99286 0 99342 800
rect 101034 0 101090 800
rect 102690 0 102746 800
rect 104438 0 104494 800
rect 106094 0 106150 800
rect 107842 0 107898 800
rect 109498 0 109554 800
rect 111246 0 111302 800
rect 112902 0 112958 800
rect 114558 0 114614 800
rect 116306 0 116362 800
rect 117962 0 118018 800
rect 119710 0 119766 800
rect 121366 0 121422 800
rect 123114 0 123170 800
rect 124770 0 124826 800
rect 126518 0 126574 800
rect 128174 0 128230 800
rect 129922 0 129978 800
rect 131578 0 131634 800
rect 133326 0 133382 800
rect 134982 0 135038 800
rect 136638 0 136694 800
rect 138386 0 138442 800
rect 140042 0 140098 800
rect 141790 0 141846 800
rect 143446 0 143502 800
rect 145194 0 145250 800
rect 146850 0 146906 800
rect 148598 0 148654 800
rect 150254 0 150310 800
rect 152002 0 152058 800
rect 153658 0 153714 800
rect 155406 0 155462 800
rect 157062 0 157118 800
rect 158718 0 158774 800
rect 160466 0 160522 800
rect 162122 0 162178 800
rect 163870 0 163926 800
rect 165526 0 165582 800
rect 167274 0 167330 800
rect 168930 0 168986 800
rect 170678 0 170734 800
rect 172334 0 172390 800
rect 174082 0 174138 800
rect 175738 0 175794 800
rect 177486 0 177542 800
rect 179142 0 179198 800
<< obsm2 >>
rect 848 139144 974 139369
rect 1142 139144 3090 139369
rect 3258 139144 5298 139369
rect 5466 139144 7506 139369
rect 7674 139144 9714 139369
rect 9882 139144 11922 139369
rect 12090 139144 14130 139369
rect 14298 139144 16338 139369
rect 16506 139144 18454 139369
rect 18622 139144 20662 139369
rect 20830 139144 22870 139369
rect 23038 139144 25078 139369
rect 25246 139144 27286 139369
rect 27454 139144 29494 139369
rect 29662 139144 31702 139369
rect 31870 139144 33818 139369
rect 33986 139144 36026 139369
rect 36194 139144 38234 139369
rect 38402 139144 40442 139369
rect 40610 139144 42650 139369
rect 42818 139144 44858 139369
rect 45026 139144 47066 139369
rect 47234 139144 49274 139369
rect 49442 139144 51390 139369
rect 51558 139144 53598 139369
rect 53766 139144 55806 139369
rect 55974 139144 58014 139369
rect 58182 139144 60222 139369
rect 60390 139144 62430 139369
rect 62598 139144 64638 139369
rect 64806 139144 66754 139369
rect 66922 139144 68962 139369
rect 69130 139144 71170 139369
rect 71338 139144 73378 139369
rect 73546 139144 75586 139369
rect 75754 139144 77794 139369
rect 77962 139144 80002 139369
rect 80170 139144 82210 139369
rect 82378 139144 84326 139369
rect 84494 139144 86534 139369
rect 86702 139144 88742 139369
rect 88910 139144 90950 139369
rect 91118 139144 93158 139369
rect 93326 139144 95366 139369
rect 95534 139144 97574 139369
rect 97742 139144 99690 139369
rect 99858 139144 101898 139369
rect 102066 139144 104106 139369
rect 104274 139144 106314 139369
rect 106482 139144 108522 139369
rect 108690 139144 110730 139369
rect 110898 139144 112938 139369
rect 113106 139144 115146 139369
rect 115314 139144 117262 139369
rect 117430 139144 119470 139369
rect 119638 139144 121678 139369
rect 121846 139144 123886 139369
rect 124054 139144 126094 139369
rect 126262 139144 128302 139369
rect 128470 139144 130510 139369
rect 130678 139144 132626 139369
rect 132794 139144 134834 139369
rect 135002 139144 137042 139369
rect 137210 139144 139250 139369
rect 139418 139144 141458 139369
rect 141626 139144 143666 139369
rect 143834 139144 145874 139369
rect 146042 139144 148082 139369
rect 148250 139144 150198 139369
rect 150366 139144 152406 139369
rect 152574 139144 154614 139369
rect 154782 139144 156822 139369
rect 156990 139144 159030 139369
rect 159198 139144 161238 139369
rect 161406 139144 163446 139369
rect 163614 139144 165562 139369
rect 165730 139144 167770 139369
rect 167938 139144 169978 139369
rect 170146 139144 172186 139369
rect 172354 139144 174394 139369
rect 174562 139144 176602 139369
rect 176770 139144 178810 139369
rect 178978 139144 179196 139369
rect 848 856 179196 139144
rect 958 575 2446 856
rect 2614 575 4102 856
rect 4270 575 5850 856
rect 6018 575 7506 856
rect 7674 575 9254 856
rect 9422 575 10910 856
rect 11078 575 12658 856
rect 12826 575 14314 856
rect 14482 575 16062 856
rect 16230 575 17718 856
rect 17886 575 19466 856
rect 19634 575 21122 856
rect 21290 575 22870 856
rect 23038 575 24526 856
rect 24694 575 26182 856
rect 26350 575 27930 856
rect 28098 575 29586 856
rect 29754 575 31334 856
rect 31502 575 32990 856
rect 33158 575 34738 856
rect 34906 575 36394 856
rect 36562 575 38142 856
rect 38310 575 39798 856
rect 39966 575 41546 856
rect 41714 575 43202 856
rect 43370 575 44950 856
rect 45118 575 46606 856
rect 46774 575 48262 856
rect 48430 575 50010 856
rect 50178 575 51666 856
rect 51834 575 53414 856
rect 53582 575 55070 856
rect 55238 575 56818 856
rect 56986 575 58474 856
rect 58642 575 60222 856
rect 60390 575 61878 856
rect 62046 575 63626 856
rect 63794 575 65282 856
rect 65450 575 67030 856
rect 67198 575 68686 856
rect 68854 575 70342 856
rect 70510 575 72090 856
rect 72258 575 73746 856
rect 73914 575 75494 856
rect 75662 575 77150 856
rect 77318 575 78898 856
rect 79066 575 80554 856
rect 80722 575 82302 856
rect 82470 575 83958 856
rect 84126 575 85706 856
rect 85874 575 87362 856
rect 87530 575 89110 856
rect 89278 575 90766 856
rect 90934 575 92422 856
rect 92590 575 94170 856
rect 94338 575 95826 856
rect 95994 575 97574 856
rect 97742 575 99230 856
rect 99398 575 100978 856
rect 101146 575 102634 856
rect 102802 575 104382 856
rect 104550 575 106038 856
rect 106206 575 107786 856
rect 107954 575 109442 856
rect 109610 575 111190 856
rect 111358 575 112846 856
rect 113014 575 114502 856
rect 114670 575 116250 856
rect 116418 575 117906 856
rect 118074 575 119654 856
rect 119822 575 121310 856
rect 121478 575 123058 856
rect 123226 575 124714 856
rect 124882 575 126462 856
rect 126630 575 128118 856
rect 128286 575 129866 856
rect 130034 575 131522 856
rect 131690 575 133270 856
rect 133438 575 134926 856
rect 135094 575 136582 856
rect 136750 575 138330 856
rect 138498 575 139986 856
rect 140154 575 141734 856
rect 141902 575 143390 856
rect 143558 575 145138 856
rect 145306 575 146794 856
rect 146962 575 148542 856
rect 148710 575 150198 856
rect 150366 575 151946 856
rect 152114 575 153602 856
rect 153770 575 155350 856
rect 155518 575 157006 856
rect 157174 575 158662 856
rect 158830 575 160410 856
rect 160578 575 162066 856
rect 162234 575 163814 856
rect 163982 575 165470 856
rect 165638 575 167218 856
rect 167386 575 168874 856
rect 169042 575 170622 856
rect 170790 575 172278 856
rect 172446 575 174026 856
rect 174194 575 175682 856
rect 175850 575 177430 856
rect 177598 575 179086 856
<< metal3 >>
rect 0 139272 800 139392
rect 179200 139136 180000 139256
rect 0 138184 800 138304
rect 179200 137912 180000 138032
rect 0 136960 800 137080
rect 179200 136552 180000 136672
rect 0 135872 800 135992
rect 179200 135328 180000 135448
rect 0 134648 800 134768
rect 179200 133968 180000 134088
rect 0 133560 800 133680
rect 179200 132744 180000 132864
rect 0 132336 800 132456
rect 0 131248 800 131368
rect 179200 131384 180000 131504
rect 0 130160 800 130280
rect 179200 130160 180000 130280
rect 0 128936 800 129056
rect 179200 128936 180000 129056
rect 0 127848 800 127968
rect 179200 127576 180000 127696
rect 0 126624 800 126744
rect 179200 126352 180000 126472
rect 0 125536 800 125656
rect 179200 124992 180000 125112
rect 0 124312 800 124432
rect 179200 123768 180000 123888
rect 0 123224 800 123344
rect 179200 122408 180000 122528
rect 0 122136 800 122256
rect 179200 121184 180000 121304
rect 0 120912 800 121032
rect 0 119824 800 119944
rect 179200 119824 180000 119944
rect 0 118600 800 118720
rect 179200 118600 180000 118720
rect 0 117512 800 117632
rect 179200 117376 180000 117496
rect 0 116288 800 116408
rect 179200 116016 180000 116136
rect 0 115200 800 115320
rect 179200 114792 180000 114912
rect 0 114112 800 114232
rect 179200 113432 180000 113552
rect 0 112888 800 113008
rect 179200 112208 180000 112328
rect 0 111800 800 111920
rect 179200 110848 180000 110968
rect 0 110576 800 110696
rect 0 109488 800 109608
rect 179200 109624 180000 109744
rect 0 108264 800 108384
rect 179200 108264 180000 108384
rect 0 107176 800 107296
rect 179200 107040 180000 107160
rect 0 105952 800 106072
rect 179200 105816 180000 105936
rect 0 104864 800 104984
rect 179200 104456 180000 104576
rect 0 103776 800 103896
rect 179200 103232 180000 103352
rect 0 102552 800 102672
rect 179200 101872 180000 101992
rect 0 101464 800 101584
rect 179200 100648 180000 100768
rect 0 100240 800 100360
rect 0 99152 800 99272
rect 179200 99288 180000 99408
rect 0 97928 800 98048
rect 179200 98064 180000 98184
rect 0 96840 800 96960
rect 179200 96840 180000 96960
rect 0 95752 800 95872
rect 179200 95480 180000 95600
rect 0 94528 800 94648
rect 179200 94256 180000 94376
rect 0 93440 800 93560
rect 179200 92896 180000 93016
rect 0 92216 800 92336
rect 179200 91672 180000 91792
rect 0 91128 800 91248
rect 179200 90312 180000 90432
rect 0 89904 800 90024
rect 179200 89088 180000 89208
rect 0 88816 800 88936
rect 0 87728 800 87848
rect 179200 87728 180000 87848
rect 0 86504 800 86624
rect 179200 86504 180000 86624
rect 0 85416 800 85536
rect 179200 85280 180000 85400
rect 0 84192 800 84312
rect 179200 83920 180000 84040
rect 0 83104 800 83224
rect 179200 82696 180000 82816
rect 0 81880 800 82000
rect 179200 81336 180000 81456
rect 0 80792 800 80912
rect 179200 80112 180000 80232
rect 0 79568 800 79688
rect 179200 78752 180000 78872
rect 0 78480 800 78600
rect 0 77392 800 77512
rect 179200 77528 180000 77648
rect 0 76168 800 76288
rect 179200 76168 180000 76288
rect 0 75080 800 75200
rect 179200 74944 180000 75064
rect 0 73856 800 73976
rect 179200 73720 180000 73840
rect 0 72768 800 72888
rect 179200 72360 180000 72480
rect 0 71544 800 71664
rect 179200 71136 180000 71256
rect 0 70456 800 70576
rect 179200 69776 180000 69896
rect 0 69368 800 69488
rect 179200 68552 180000 68672
rect 0 68144 800 68264
rect 0 67056 800 67176
rect 179200 67192 180000 67312
rect 0 65832 800 65952
rect 179200 65968 180000 66088
rect 0 64744 800 64864
rect 179200 64744 180000 64864
rect 0 63520 800 63640
rect 179200 63384 180000 63504
rect 0 62432 800 62552
rect 179200 62160 180000 62280
rect 0 61344 800 61464
rect 179200 60800 180000 60920
rect 0 60120 800 60240
rect 179200 59576 180000 59696
rect 0 59032 800 59152
rect 179200 58216 180000 58336
rect 0 57808 800 57928
rect 179200 56992 180000 57112
rect 0 56720 800 56840
rect 0 55496 800 55616
rect 179200 55632 180000 55752
rect 0 54408 800 54528
rect 179200 54408 180000 54528
rect 0 53184 800 53304
rect 179200 53184 180000 53304
rect 0 52096 800 52216
rect 179200 51824 180000 51944
rect 0 51008 800 51128
rect 179200 50600 180000 50720
rect 0 49784 800 49904
rect 179200 49240 180000 49360
rect 0 48696 800 48816
rect 179200 48016 180000 48136
rect 0 47472 800 47592
rect 179200 46656 180000 46776
rect 0 46384 800 46504
rect 179200 45432 180000 45552
rect 0 45160 800 45280
rect 0 44072 800 44192
rect 179200 44072 180000 44192
rect 0 42984 800 43104
rect 179200 42848 180000 42968
rect 0 41760 800 41880
rect 179200 41624 180000 41744
rect 0 40672 800 40792
rect 179200 40264 180000 40384
rect 0 39448 800 39568
rect 179200 39040 180000 39160
rect 0 38360 800 38480
rect 179200 37680 180000 37800
rect 0 37136 800 37256
rect 179200 36456 180000 36576
rect 0 36048 800 36168
rect 0 34960 800 35080
rect 179200 35096 180000 35216
rect 0 33736 800 33856
rect 179200 33872 180000 33992
rect 0 32648 800 32768
rect 179200 32648 180000 32768
rect 0 31424 800 31544
rect 179200 31288 180000 31408
rect 0 30336 800 30456
rect 179200 30064 180000 30184
rect 0 29112 800 29232
rect 179200 28704 180000 28824
rect 0 28024 800 28144
rect 179200 27480 180000 27600
rect 0 26800 800 26920
rect 179200 26120 180000 26240
rect 0 25712 800 25832
rect 179200 24896 180000 25016
rect 0 24624 800 24744
rect 0 23400 800 23520
rect 179200 23536 180000 23656
rect 0 22312 800 22432
rect 179200 22312 180000 22432
rect 0 21088 800 21208
rect 179200 21088 180000 21208
rect 0 20000 800 20120
rect 179200 19728 180000 19848
rect 0 18776 800 18896
rect 179200 18504 180000 18624
rect 0 17688 800 17808
rect 179200 17144 180000 17264
rect 0 16600 800 16720
rect 179200 15920 180000 16040
rect 0 15376 800 15496
rect 179200 14560 180000 14680
rect 0 14288 800 14408
rect 179200 13336 180000 13456
rect 0 13064 800 13184
rect 0 11976 800 12096
rect 179200 11976 180000 12096
rect 0 10752 800 10872
rect 179200 10752 180000 10872
rect 0 9664 800 9784
rect 179200 9528 180000 9648
rect 0 8576 800 8696
rect 179200 8168 180000 8288
rect 0 7352 800 7472
rect 179200 6944 180000 7064
rect 0 6264 800 6384
rect 179200 5584 180000 5704
rect 0 5040 800 5160
rect 179200 4360 180000 4480
rect 0 3952 800 4072
rect 179200 3000 180000 3120
rect 0 2728 800 2848
rect 0 1640 800 1760
rect 179200 1776 180000 1896
rect 0 552 800 672
rect 179200 552 180000 672
<< obsm3 >>
rect 880 139336 179200 139365
rect 880 139192 179120 139336
rect 800 139056 179120 139192
rect 800 138384 179200 139056
rect 880 138112 179200 138384
rect 880 138104 179120 138112
rect 800 137832 179120 138104
rect 800 137160 179200 137832
rect 880 136880 179200 137160
rect 800 136752 179200 136880
rect 800 136472 179120 136752
rect 800 136072 179200 136472
rect 880 135792 179200 136072
rect 800 135528 179200 135792
rect 800 135248 179120 135528
rect 800 134848 179200 135248
rect 880 134568 179200 134848
rect 800 134168 179200 134568
rect 800 133888 179120 134168
rect 800 133760 179200 133888
rect 880 133480 179200 133760
rect 800 132944 179200 133480
rect 800 132664 179120 132944
rect 800 132536 179200 132664
rect 880 132256 179200 132536
rect 800 131584 179200 132256
rect 800 131448 179120 131584
rect 880 131304 179120 131448
rect 880 131168 179200 131304
rect 800 130360 179200 131168
rect 880 130080 179120 130360
rect 800 129136 179200 130080
rect 880 128856 179120 129136
rect 800 128048 179200 128856
rect 880 127776 179200 128048
rect 880 127768 179120 127776
rect 800 127496 179120 127768
rect 800 126824 179200 127496
rect 880 126552 179200 126824
rect 880 126544 179120 126552
rect 800 126272 179120 126544
rect 800 125736 179200 126272
rect 880 125456 179200 125736
rect 800 125192 179200 125456
rect 800 124912 179120 125192
rect 800 124512 179200 124912
rect 880 124232 179200 124512
rect 800 123968 179200 124232
rect 800 123688 179120 123968
rect 800 123424 179200 123688
rect 880 123144 179200 123424
rect 800 122608 179200 123144
rect 800 122336 179120 122608
rect 880 122328 179120 122336
rect 880 122056 179200 122328
rect 800 121384 179200 122056
rect 800 121112 179120 121384
rect 880 121104 179120 121112
rect 880 120832 179200 121104
rect 800 120024 179200 120832
rect 880 119744 179120 120024
rect 800 118800 179200 119744
rect 880 118520 179120 118800
rect 800 117712 179200 118520
rect 880 117576 179200 117712
rect 880 117432 179120 117576
rect 800 117296 179120 117432
rect 800 116488 179200 117296
rect 880 116216 179200 116488
rect 880 116208 179120 116216
rect 800 115936 179120 116208
rect 800 115400 179200 115936
rect 880 115120 179200 115400
rect 800 114992 179200 115120
rect 800 114712 179120 114992
rect 800 114312 179200 114712
rect 880 114032 179200 114312
rect 800 113632 179200 114032
rect 800 113352 179120 113632
rect 800 113088 179200 113352
rect 880 112808 179200 113088
rect 800 112408 179200 112808
rect 800 112128 179120 112408
rect 800 112000 179200 112128
rect 880 111720 179200 112000
rect 800 111048 179200 111720
rect 800 110776 179120 111048
rect 880 110768 179120 110776
rect 880 110496 179200 110768
rect 800 109824 179200 110496
rect 800 109688 179120 109824
rect 880 109544 179120 109688
rect 880 109408 179200 109544
rect 800 108464 179200 109408
rect 880 108184 179120 108464
rect 800 107376 179200 108184
rect 880 107240 179200 107376
rect 880 107096 179120 107240
rect 800 106960 179120 107096
rect 800 106152 179200 106960
rect 880 106016 179200 106152
rect 880 105872 179120 106016
rect 800 105736 179120 105872
rect 800 105064 179200 105736
rect 880 104784 179200 105064
rect 800 104656 179200 104784
rect 800 104376 179120 104656
rect 800 103976 179200 104376
rect 880 103696 179200 103976
rect 800 103432 179200 103696
rect 800 103152 179120 103432
rect 800 102752 179200 103152
rect 880 102472 179200 102752
rect 800 102072 179200 102472
rect 800 101792 179120 102072
rect 800 101664 179200 101792
rect 880 101384 179200 101664
rect 800 100848 179200 101384
rect 800 100568 179120 100848
rect 800 100440 179200 100568
rect 880 100160 179200 100440
rect 800 99488 179200 100160
rect 800 99352 179120 99488
rect 880 99208 179120 99352
rect 880 99072 179200 99208
rect 800 98264 179200 99072
rect 800 98128 179120 98264
rect 880 97984 179120 98128
rect 880 97848 179200 97984
rect 800 97040 179200 97848
rect 880 96760 179120 97040
rect 800 95952 179200 96760
rect 880 95680 179200 95952
rect 880 95672 179120 95680
rect 800 95400 179120 95672
rect 800 94728 179200 95400
rect 880 94456 179200 94728
rect 880 94448 179120 94456
rect 800 94176 179120 94448
rect 800 93640 179200 94176
rect 880 93360 179200 93640
rect 800 93096 179200 93360
rect 800 92816 179120 93096
rect 800 92416 179200 92816
rect 880 92136 179200 92416
rect 800 91872 179200 92136
rect 800 91592 179120 91872
rect 800 91328 179200 91592
rect 880 91048 179200 91328
rect 800 90512 179200 91048
rect 800 90232 179120 90512
rect 800 90104 179200 90232
rect 880 89824 179200 90104
rect 800 89288 179200 89824
rect 800 89016 179120 89288
rect 880 89008 179120 89016
rect 880 88736 179200 89008
rect 800 87928 179200 88736
rect 880 87648 179120 87928
rect 800 86704 179200 87648
rect 880 86424 179120 86704
rect 800 85616 179200 86424
rect 880 85480 179200 85616
rect 880 85336 179120 85480
rect 800 85200 179120 85336
rect 800 84392 179200 85200
rect 880 84120 179200 84392
rect 880 84112 179120 84120
rect 800 83840 179120 84112
rect 800 83304 179200 83840
rect 880 83024 179200 83304
rect 800 82896 179200 83024
rect 800 82616 179120 82896
rect 800 82080 179200 82616
rect 880 81800 179200 82080
rect 800 81536 179200 81800
rect 800 81256 179120 81536
rect 800 80992 179200 81256
rect 880 80712 179200 80992
rect 800 80312 179200 80712
rect 800 80032 179120 80312
rect 800 79768 179200 80032
rect 880 79488 179200 79768
rect 800 78952 179200 79488
rect 800 78680 179120 78952
rect 880 78672 179120 78680
rect 880 78400 179200 78672
rect 800 77728 179200 78400
rect 800 77592 179120 77728
rect 880 77448 179120 77592
rect 880 77312 179200 77448
rect 800 76368 179200 77312
rect 880 76088 179120 76368
rect 800 75280 179200 76088
rect 880 75144 179200 75280
rect 880 75000 179120 75144
rect 800 74864 179120 75000
rect 800 74056 179200 74864
rect 880 73920 179200 74056
rect 880 73776 179120 73920
rect 800 73640 179120 73776
rect 800 72968 179200 73640
rect 880 72688 179200 72968
rect 800 72560 179200 72688
rect 800 72280 179120 72560
rect 800 71744 179200 72280
rect 880 71464 179200 71744
rect 800 71336 179200 71464
rect 800 71056 179120 71336
rect 800 70656 179200 71056
rect 880 70376 179200 70656
rect 800 69976 179200 70376
rect 800 69696 179120 69976
rect 800 69568 179200 69696
rect 880 69288 179200 69568
rect 800 68752 179200 69288
rect 800 68472 179120 68752
rect 800 68344 179200 68472
rect 880 68064 179200 68344
rect 800 67392 179200 68064
rect 800 67256 179120 67392
rect 880 67112 179120 67256
rect 880 66976 179200 67112
rect 800 66168 179200 66976
rect 800 66032 179120 66168
rect 880 65888 179120 66032
rect 880 65752 179200 65888
rect 800 64944 179200 65752
rect 880 64664 179120 64944
rect 800 63720 179200 64664
rect 880 63584 179200 63720
rect 880 63440 179120 63584
rect 800 63304 179120 63440
rect 800 62632 179200 63304
rect 880 62360 179200 62632
rect 880 62352 179120 62360
rect 800 62080 179120 62352
rect 800 61544 179200 62080
rect 880 61264 179200 61544
rect 800 61000 179200 61264
rect 800 60720 179120 61000
rect 800 60320 179200 60720
rect 880 60040 179200 60320
rect 800 59776 179200 60040
rect 800 59496 179120 59776
rect 800 59232 179200 59496
rect 880 58952 179200 59232
rect 800 58416 179200 58952
rect 800 58136 179120 58416
rect 800 58008 179200 58136
rect 880 57728 179200 58008
rect 800 57192 179200 57728
rect 800 56920 179120 57192
rect 880 56912 179120 56920
rect 880 56640 179200 56912
rect 800 55832 179200 56640
rect 800 55696 179120 55832
rect 880 55552 179120 55696
rect 880 55416 179200 55552
rect 800 54608 179200 55416
rect 880 54328 179120 54608
rect 800 53384 179200 54328
rect 880 53104 179120 53384
rect 800 52296 179200 53104
rect 880 52024 179200 52296
rect 880 52016 179120 52024
rect 800 51744 179120 52016
rect 800 51208 179200 51744
rect 880 50928 179200 51208
rect 800 50800 179200 50928
rect 800 50520 179120 50800
rect 800 49984 179200 50520
rect 880 49704 179200 49984
rect 800 49440 179200 49704
rect 800 49160 179120 49440
rect 800 48896 179200 49160
rect 880 48616 179200 48896
rect 800 48216 179200 48616
rect 800 47936 179120 48216
rect 800 47672 179200 47936
rect 880 47392 179200 47672
rect 800 46856 179200 47392
rect 800 46584 179120 46856
rect 880 46576 179120 46584
rect 880 46304 179200 46576
rect 800 45632 179200 46304
rect 800 45360 179120 45632
rect 880 45352 179120 45360
rect 880 45080 179200 45352
rect 800 44272 179200 45080
rect 880 43992 179120 44272
rect 800 43184 179200 43992
rect 880 43048 179200 43184
rect 880 42904 179120 43048
rect 800 42768 179120 42904
rect 800 41960 179200 42768
rect 880 41824 179200 41960
rect 880 41680 179120 41824
rect 800 41544 179120 41680
rect 800 40872 179200 41544
rect 880 40592 179200 40872
rect 800 40464 179200 40592
rect 800 40184 179120 40464
rect 800 39648 179200 40184
rect 880 39368 179200 39648
rect 800 39240 179200 39368
rect 800 38960 179120 39240
rect 800 38560 179200 38960
rect 880 38280 179200 38560
rect 800 37880 179200 38280
rect 800 37600 179120 37880
rect 800 37336 179200 37600
rect 880 37056 179200 37336
rect 800 36656 179200 37056
rect 800 36376 179120 36656
rect 800 36248 179200 36376
rect 880 35968 179200 36248
rect 800 35296 179200 35968
rect 800 35160 179120 35296
rect 880 35016 179120 35160
rect 880 34880 179200 35016
rect 800 34072 179200 34880
rect 800 33936 179120 34072
rect 880 33792 179120 33936
rect 880 33656 179200 33792
rect 800 32848 179200 33656
rect 880 32568 179120 32848
rect 800 31624 179200 32568
rect 880 31488 179200 31624
rect 880 31344 179120 31488
rect 800 31208 179120 31344
rect 800 30536 179200 31208
rect 880 30264 179200 30536
rect 880 30256 179120 30264
rect 800 29984 179120 30256
rect 800 29312 179200 29984
rect 880 29032 179200 29312
rect 800 28904 179200 29032
rect 800 28624 179120 28904
rect 800 28224 179200 28624
rect 880 27944 179200 28224
rect 800 27680 179200 27944
rect 800 27400 179120 27680
rect 800 27000 179200 27400
rect 880 26720 179200 27000
rect 800 26320 179200 26720
rect 800 26040 179120 26320
rect 800 25912 179200 26040
rect 880 25632 179200 25912
rect 800 25096 179200 25632
rect 800 24824 179120 25096
rect 880 24816 179120 24824
rect 880 24544 179200 24816
rect 800 23736 179200 24544
rect 800 23600 179120 23736
rect 880 23456 179120 23600
rect 880 23320 179200 23456
rect 800 22512 179200 23320
rect 880 22232 179120 22512
rect 800 21288 179200 22232
rect 880 21008 179120 21288
rect 800 20200 179200 21008
rect 880 19928 179200 20200
rect 880 19920 179120 19928
rect 800 19648 179120 19920
rect 800 18976 179200 19648
rect 880 18704 179200 18976
rect 880 18696 179120 18704
rect 800 18424 179120 18696
rect 800 17888 179200 18424
rect 880 17608 179200 17888
rect 800 17344 179200 17608
rect 800 17064 179120 17344
rect 800 16800 179200 17064
rect 880 16520 179200 16800
rect 800 16120 179200 16520
rect 800 15840 179120 16120
rect 800 15576 179200 15840
rect 880 15296 179200 15576
rect 800 14760 179200 15296
rect 800 14488 179120 14760
rect 880 14480 179120 14488
rect 880 14208 179200 14480
rect 800 13536 179200 14208
rect 800 13264 179120 13536
rect 880 13256 179120 13264
rect 880 12984 179200 13256
rect 800 12176 179200 12984
rect 880 11896 179120 12176
rect 800 10952 179200 11896
rect 880 10672 179120 10952
rect 800 9864 179200 10672
rect 880 9728 179200 9864
rect 880 9584 179120 9728
rect 800 9448 179120 9584
rect 800 8776 179200 9448
rect 880 8496 179200 8776
rect 800 8368 179200 8496
rect 800 8088 179120 8368
rect 800 7552 179200 8088
rect 880 7272 179200 7552
rect 800 7144 179200 7272
rect 800 6864 179120 7144
rect 800 6464 179200 6864
rect 880 6184 179200 6464
rect 800 5784 179200 6184
rect 800 5504 179120 5784
rect 800 5240 179200 5504
rect 880 4960 179200 5240
rect 800 4560 179200 4960
rect 800 4280 179120 4560
rect 800 4152 179200 4280
rect 880 3872 179200 4152
rect 800 3200 179200 3872
rect 800 2928 179120 3200
rect 880 2920 179120 2928
rect 880 2648 179200 2920
rect 800 1976 179200 2648
rect 800 1840 179120 1976
rect 880 1696 179120 1840
rect 880 1560 179200 1696
rect 800 752 179200 1560
rect 880 579 179120 752
<< metal4 >>
rect 4208 2128 4528 137680
rect 4868 2176 5188 137632
rect 5528 2176 5848 137632
rect 6188 2176 6508 137632
rect 19568 2128 19888 137680
rect 20228 2176 20548 137632
rect 20888 2176 21208 137632
rect 21548 2176 21868 137632
rect 34928 2128 35248 137680
rect 35588 2176 35908 137632
rect 36248 2176 36568 137632
rect 36908 2176 37228 137632
rect 50288 2128 50608 137680
rect 50948 2176 51268 137632
rect 51608 2176 51928 137632
rect 52268 2176 52588 137632
rect 65648 2128 65968 137680
rect 66308 2176 66628 137632
rect 66968 2176 67288 137632
rect 67628 2176 67948 137632
rect 81008 2128 81328 137680
rect 81668 2176 81988 137632
rect 82328 2176 82648 137632
rect 82988 2176 83308 137632
rect 96368 2128 96688 137680
rect 97028 2176 97348 137632
rect 97688 2176 98008 137632
rect 98348 2176 98668 137632
rect 111728 2128 112048 137680
rect 112388 2176 112708 137632
rect 113048 2176 113368 137632
rect 113708 2176 114028 137632
rect 127088 2128 127408 137680
rect 127748 2176 128068 137632
rect 128408 2176 128728 137632
rect 129068 2176 129388 137632
rect 142448 2128 142768 137680
rect 143108 2176 143428 137632
rect 143768 2176 144088 137632
rect 144428 2176 144748 137632
rect 157808 2128 158128 137680
rect 158468 2176 158788 137632
rect 159128 2176 159448 137632
rect 159788 2176 160108 137632
rect 173168 2128 173488 137680
rect 173828 2176 174148 137632
rect 174488 2176 174808 137632
rect 175148 2176 175468 137632
<< obsm4 >>
rect 80007 2891 80928 137189
rect 81408 2891 81588 137189
rect 82068 2891 82248 137189
rect 82728 2891 82908 137189
rect 83388 2891 96288 137189
rect 96768 2891 96948 137189
rect 97428 2891 97608 137189
rect 98088 2891 98268 137189
rect 98748 2891 111648 137189
rect 112128 2891 112308 137189
rect 112788 2891 112968 137189
rect 113448 2891 113628 137189
rect 114108 2891 127008 137189
rect 127488 2891 127668 137189
rect 128148 2891 128328 137189
rect 128808 2891 128988 137189
rect 129468 2891 142368 137189
rect 142848 2891 143028 137189
rect 143508 2891 143688 137189
rect 144168 2891 144348 137189
rect 144828 2891 157728 137189
rect 158208 2891 158388 137189
rect 158868 2891 159048 137189
rect 159528 2891 159708 137189
rect 160188 2891 173088 137189
rect 173568 2891 173748 137189
rect 174228 2891 174408 137189
rect 174888 2891 175068 137189
rect 175548 2891 177869 137189
<< labels >>
rlabel metal3 s 179200 552 180000 672 6 adc0_dat_i[0]
port 1 nsew signal input
rlabel metal3 s 179200 42848 180000 42968 6 adc0_dat_i[10]
port 2 nsew signal input
rlabel metal3 s 179200 46656 180000 46776 6 adc0_dat_i[11]
port 3 nsew signal input
rlabel metal3 s 179200 50600 180000 50720 6 adc0_dat_i[12]
port 4 nsew signal input
rlabel metal3 s 179200 54408 180000 54528 6 adc0_dat_i[13]
port 5 nsew signal input
rlabel metal3 s 179200 58216 180000 58336 6 adc0_dat_i[14]
port 6 nsew signal input
rlabel metal3 s 179200 62160 180000 62280 6 adc0_dat_i[15]
port 7 nsew signal input
rlabel metal3 s 179200 65968 180000 66088 6 adc0_dat_i[16]
port 8 nsew signal input
rlabel metal3 s 179200 69776 180000 69896 6 adc0_dat_i[17]
port 9 nsew signal input
rlabel metal3 s 179200 73720 180000 73840 6 adc0_dat_i[18]
port 10 nsew signal input
rlabel metal3 s 179200 77528 180000 77648 6 adc0_dat_i[19]
port 11 nsew signal input
rlabel metal3 s 179200 5584 180000 5704 6 adc0_dat_i[1]
port 12 nsew signal input
rlabel metal3 s 179200 81336 180000 81456 6 adc0_dat_i[20]
port 13 nsew signal input
rlabel metal3 s 179200 85280 180000 85400 6 adc0_dat_i[21]
port 14 nsew signal input
rlabel metal3 s 179200 89088 180000 89208 6 adc0_dat_i[22]
port 15 nsew signal input
rlabel metal3 s 179200 92896 180000 93016 6 adc0_dat_i[23]
port 16 nsew signal input
rlabel metal3 s 179200 96840 180000 96960 6 adc0_dat_i[24]
port 17 nsew signal input
rlabel metal3 s 179200 100648 180000 100768 6 adc0_dat_i[25]
port 18 nsew signal input
rlabel metal3 s 179200 104456 180000 104576 6 adc0_dat_i[26]
port 19 nsew signal input
rlabel metal3 s 179200 108264 180000 108384 6 adc0_dat_i[27]
port 20 nsew signal input
rlabel metal3 s 179200 112208 180000 112328 6 adc0_dat_i[28]
port 21 nsew signal input
rlabel metal3 s 179200 116016 180000 116136 6 adc0_dat_i[29]
port 22 nsew signal input
rlabel metal3 s 179200 10752 180000 10872 6 adc0_dat_i[2]
port 23 nsew signal input
rlabel metal3 s 179200 119824 180000 119944 6 adc0_dat_i[30]
port 24 nsew signal input
rlabel metal3 s 179200 123768 180000 123888 6 adc0_dat_i[31]
port 25 nsew signal input
rlabel metal3 s 179200 15920 180000 16040 6 adc0_dat_i[3]
port 26 nsew signal input
rlabel metal3 s 179200 19728 180000 19848 6 adc0_dat_i[4]
port 27 nsew signal input
rlabel metal3 s 179200 23536 180000 23656 6 adc0_dat_i[5]
port 28 nsew signal input
rlabel metal3 s 179200 27480 180000 27600 6 adc0_dat_i[6]
port 29 nsew signal input
rlabel metal3 s 179200 31288 180000 31408 6 adc0_dat_i[7]
port 30 nsew signal input
rlabel metal3 s 179200 35096 180000 35216 6 adc0_dat_i[8]
port 31 nsew signal input
rlabel metal3 s 179200 39040 180000 39160 6 adc0_dat_i[9]
port 32 nsew signal input
rlabel metal3 s 179200 1776 180000 1896 6 adc1_dat_i[0]
port 33 nsew signal input
rlabel metal3 s 179200 44072 180000 44192 6 adc1_dat_i[10]
port 34 nsew signal input
rlabel metal3 s 179200 48016 180000 48136 6 adc1_dat_i[11]
port 35 nsew signal input
rlabel metal3 s 179200 51824 180000 51944 6 adc1_dat_i[12]
port 36 nsew signal input
rlabel metal3 s 179200 55632 180000 55752 6 adc1_dat_i[13]
port 37 nsew signal input
rlabel metal3 s 179200 59576 180000 59696 6 adc1_dat_i[14]
port 38 nsew signal input
rlabel metal3 s 179200 63384 180000 63504 6 adc1_dat_i[15]
port 39 nsew signal input
rlabel metal3 s 179200 67192 180000 67312 6 adc1_dat_i[16]
port 40 nsew signal input
rlabel metal3 s 179200 71136 180000 71256 6 adc1_dat_i[17]
port 41 nsew signal input
rlabel metal3 s 179200 74944 180000 75064 6 adc1_dat_i[18]
port 42 nsew signal input
rlabel metal3 s 179200 78752 180000 78872 6 adc1_dat_i[19]
port 43 nsew signal input
rlabel metal3 s 179200 6944 180000 7064 6 adc1_dat_i[1]
port 44 nsew signal input
rlabel metal3 s 179200 82696 180000 82816 6 adc1_dat_i[20]
port 45 nsew signal input
rlabel metal3 s 179200 86504 180000 86624 6 adc1_dat_i[21]
port 46 nsew signal input
rlabel metal3 s 179200 90312 180000 90432 6 adc1_dat_i[22]
port 47 nsew signal input
rlabel metal3 s 179200 94256 180000 94376 6 adc1_dat_i[23]
port 48 nsew signal input
rlabel metal3 s 179200 98064 180000 98184 6 adc1_dat_i[24]
port 49 nsew signal input
rlabel metal3 s 179200 101872 180000 101992 6 adc1_dat_i[25]
port 50 nsew signal input
rlabel metal3 s 179200 105816 180000 105936 6 adc1_dat_i[26]
port 51 nsew signal input
rlabel metal3 s 179200 109624 180000 109744 6 adc1_dat_i[27]
port 52 nsew signal input
rlabel metal3 s 179200 113432 180000 113552 6 adc1_dat_i[28]
port 53 nsew signal input
rlabel metal3 s 179200 117376 180000 117496 6 adc1_dat_i[29]
port 54 nsew signal input
rlabel metal3 s 179200 11976 180000 12096 6 adc1_dat_i[2]
port 55 nsew signal input
rlabel metal3 s 179200 121184 180000 121304 6 adc1_dat_i[30]
port 56 nsew signal input
rlabel metal3 s 179200 124992 180000 125112 6 adc1_dat_i[31]
port 57 nsew signal input
rlabel metal3 s 179200 17144 180000 17264 6 adc1_dat_i[3]
port 58 nsew signal input
rlabel metal3 s 179200 21088 180000 21208 6 adc1_dat_i[4]
port 59 nsew signal input
rlabel metal3 s 179200 24896 180000 25016 6 adc1_dat_i[5]
port 60 nsew signal input
rlabel metal3 s 179200 28704 180000 28824 6 adc1_dat_i[6]
port 61 nsew signal input
rlabel metal3 s 179200 32648 180000 32768 6 adc1_dat_i[7]
port 62 nsew signal input
rlabel metal3 s 179200 36456 180000 36576 6 adc1_dat_i[8]
port 63 nsew signal input
rlabel metal3 s 179200 40264 180000 40384 6 adc1_dat_i[9]
port 64 nsew signal input
rlabel metal3 s 179200 3000 180000 3120 6 adc2_dat_i[0]
port 65 nsew signal input
rlabel metal3 s 179200 45432 180000 45552 6 adc2_dat_i[10]
port 66 nsew signal input
rlabel metal3 s 179200 49240 180000 49360 6 adc2_dat_i[11]
port 67 nsew signal input
rlabel metal3 s 179200 53184 180000 53304 6 adc2_dat_i[12]
port 68 nsew signal input
rlabel metal3 s 179200 56992 180000 57112 6 adc2_dat_i[13]
port 69 nsew signal input
rlabel metal3 s 179200 60800 180000 60920 6 adc2_dat_i[14]
port 70 nsew signal input
rlabel metal3 s 179200 64744 180000 64864 6 adc2_dat_i[15]
port 71 nsew signal input
rlabel metal3 s 179200 68552 180000 68672 6 adc2_dat_i[16]
port 72 nsew signal input
rlabel metal3 s 179200 72360 180000 72480 6 adc2_dat_i[17]
port 73 nsew signal input
rlabel metal3 s 179200 76168 180000 76288 6 adc2_dat_i[18]
port 74 nsew signal input
rlabel metal3 s 179200 80112 180000 80232 6 adc2_dat_i[19]
port 75 nsew signal input
rlabel metal3 s 179200 8168 180000 8288 6 adc2_dat_i[1]
port 76 nsew signal input
rlabel metal3 s 179200 83920 180000 84040 6 adc2_dat_i[20]
port 77 nsew signal input
rlabel metal3 s 179200 87728 180000 87848 6 adc2_dat_i[21]
port 78 nsew signal input
rlabel metal3 s 179200 91672 180000 91792 6 adc2_dat_i[22]
port 79 nsew signal input
rlabel metal3 s 179200 95480 180000 95600 6 adc2_dat_i[23]
port 80 nsew signal input
rlabel metal3 s 179200 99288 180000 99408 6 adc2_dat_i[24]
port 81 nsew signal input
rlabel metal3 s 179200 103232 180000 103352 6 adc2_dat_i[25]
port 82 nsew signal input
rlabel metal3 s 179200 107040 180000 107160 6 adc2_dat_i[26]
port 83 nsew signal input
rlabel metal3 s 179200 110848 180000 110968 6 adc2_dat_i[27]
port 84 nsew signal input
rlabel metal3 s 179200 114792 180000 114912 6 adc2_dat_i[28]
port 85 nsew signal input
rlabel metal3 s 179200 118600 180000 118720 6 adc2_dat_i[29]
port 86 nsew signal input
rlabel metal3 s 179200 13336 180000 13456 6 adc2_dat_i[2]
port 87 nsew signal input
rlabel metal3 s 179200 122408 180000 122528 6 adc2_dat_i[30]
port 88 nsew signal input
rlabel metal3 s 179200 126352 180000 126472 6 adc2_dat_i[31]
port 89 nsew signal input
rlabel metal3 s 179200 18504 180000 18624 6 adc2_dat_i[3]
port 90 nsew signal input
rlabel metal3 s 179200 22312 180000 22432 6 adc2_dat_i[4]
port 91 nsew signal input
rlabel metal3 s 179200 26120 180000 26240 6 adc2_dat_i[5]
port 92 nsew signal input
rlabel metal3 s 179200 30064 180000 30184 6 adc2_dat_i[6]
port 93 nsew signal input
rlabel metal3 s 179200 33872 180000 33992 6 adc2_dat_i[7]
port 94 nsew signal input
rlabel metal3 s 179200 37680 180000 37800 6 adc2_dat_i[8]
port 95 nsew signal input
rlabel metal3 s 179200 41624 180000 41744 6 adc2_dat_i[9]
port 96 nsew signal input
rlabel metal3 s 179200 4360 180000 4480 6 adc_dvalid_i[0]
port 97 nsew signal input
rlabel metal3 s 179200 9528 180000 9648 6 adc_dvalid_i[1]
port 98 nsew signal input
rlabel metal3 s 179200 14560 180000 14680 6 adc_dvalid_i[2]
port 99 nsew signal input
rlabel metal2 s 1030 139200 1086 140000 6 io_oeb[0]
port 100 nsew signal output
rlabel metal2 s 44914 139200 44970 140000 6 io_oeb[10]
port 101 nsew signal output
rlabel metal2 s 49330 139200 49386 140000 6 io_oeb[11]
port 102 nsew signal output
rlabel metal2 s 53654 139200 53710 140000 6 io_oeb[12]
port 103 nsew signal output
rlabel metal2 s 58070 139200 58126 140000 6 io_oeb[13]
port 104 nsew signal output
rlabel metal2 s 62486 139200 62542 140000 6 io_oeb[14]
port 105 nsew signal output
rlabel metal2 s 66810 139200 66866 140000 6 io_oeb[15]
port 106 nsew signal output
rlabel metal2 s 71226 139200 71282 140000 6 io_oeb[16]
port 107 nsew signal output
rlabel metal2 s 75642 139200 75698 140000 6 io_oeb[17]
port 108 nsew signal output
rlabel metal2 s 80058 139200 80114 140000 6 io_oeb[18]
port 109 nsew signal output
rlabel metal2 s 84382 139200 84438 140000 6 io_oeb[19]
port 110 nsew signal output
rlabel metal2 s 5354 139200 5410 140000 6 io_oeb[1]
port 111 nsew signal output
rlabel metal2 s 88798 139200 88854 140000 6 io_oeb[20]
port 112 nsew signal output
rlabel metal2 s 93214 139200 93270 140000 6 io_oeb[21]
port 113 nsew signal output
rlabel metal2 s 97630 139200 97686 140000 6 io_oeb[22]
port 114 nsew signal output
rlabel metal2 s 101954 139200 102010 140000 6 io_oeb[23]
port 115 nsew signal output
rlabel metal2 s 106370 139200 106426 140000 6 io_oeb[24]
port 116 nsew signal output
rlabel metal2 s 110786 139200 110842 140000 6 io_oeb[25]
port 117 nsew signal output
rlabel metal2 s 115202 139200 115258 140000 6 io_oeb[26]
port 118 nsew signal output
rlabel metal2 s 119526 139200 119582 140000 6 io_oeb[27]
port 119 nsew signal output
rlabel metal2 s 123942 139200 123998 140000 6 io_oeb[28]
port 120 nsew signal output
rlabel metal2 s 128358 139200 128414 140000 6 io_oeb[29]
port 121 nsew signal output
rlabel metal2 s 9770 139200 9826 140000 6 io_oeb[2]
port 122 nsew signal output
rlabel metal2 s 132682 139200 132738 140000 6 io_oeb[30]
port 123 nsew signal output
rlabel metal2 s 137098 139200 137154 140000 6 io_oeb[31]
port 124 nsew signal output
rlabel metal2 s 141514 139200 141570 140000 6 io_oeb[32]
port 125 nsew signal output
rlabel metal2 s 145930 139200 145986 140000 6 io_oeb[33]
port 126 nsew signal output
rlabel metal2 s 150254 139200 150310 140000 6 io_oeb[34]
port 127 nsew signal output
rlabel metal2 s 154670 139200 154726 140000 6 io_oeb[35]
port 128 nsew signal output
rlabel metal2 s 159086 139200 159142 140000 6 io_oeb[36]
port 129 nsew signal output
rlabel metal2 s 163502 139200 163558 140000 6 io_oeb[37]
port 130 nsew signal output
rlabel metal2 s 14186 139200 14242 140000 6 io_oeb[3]
port 131 nsew signal output
rlabel metal2 s 18510 139200 18566 140000 6 io_oeb[4]
port 132 nsew signal output
rlabel metal2 s 22926 139200 22982 140000 6 io_oeb[5]
port 133 nsew signal output
rlabel metal2 s 27342 139200 27398 140000 6 io_oeb[6]
port 134 nsew signal output
rlabel metal2 s 31758 139200 31814 140000 6 io_oeb[7]
port 135 nsew signal output
rlabel metal2 s 36082 139200 36138 140000 6 io_oeb[8]
port 136 nsew signal output
rlabel metal2 s 40498 139200 40554 140000 6 io_oeb[9]
port 137 nsew signal output
rlabel metal2 s 3146 139200 3202 140000 6 io_out[0]
port 138 nsew signal output
rlabel metal2 s 47122 139200 47178 140000 6 io_out[10]
port 139 nsew signal output
rlabel metal2 s 51446 139200 51502 140000 6 io_out[11]
port 140 nsew signal output
rlabel metal2 s 55862 139200 55918 140000 6 io_out[12]
port 141 nsew signal output
rlabel metal2 s 60278 139200 60334 140000 6 io_out[13]
port 142 nsew signal output
rlabel metal2 s 64694 139200 64750 140000 6 io_out[14]
port 143 nsew signal output
rlabel metal2 s 69018 139200 69074 140000 6 io_out[15]
port 144 nsew signal output
rlabel metal2 s 73434 139200 73490 140000 6 io_out[16]
port 145 nsew signal output
rlabel metal2 s 77850 139200 77906 140000 6 io_out[17]
port 146 nsew signal output
rlabel metal2 s 82266 139200 82322 140000 6 io_out[18]
port 147 nsew signal output
rlabel metal2 s 86590 139200 86646 140000 6 io_out[19]
port 148 nsew signal output
rlabel metal2 s 7562 139200 7618 140000 6 io_out[1]
port 149 nsew signal output
rlabel metal2 s 91006 139200 91062 140000 6 io_out[20]
port 150 nsew signal output
rlabel metal2 s 95422 139200 95478 140000 6 io_out[21]
port 151 nsew signal output
rlabel metal2 s 99746 139200 99802 140000 6 io_out[22]
port 152 nsew signal output
rlabel metal2 s 104162 139200 104218 140000 6 io_out[23]
port 153 nsew signal output
rlabel metal2 s 108578 139200 108634 140000 6 io_out[24]
port 154 nsew signal output
rlabel metal2 s 112994 139200 113050 140000 6 io_out[25]
port 155 nsew signal output
rlabel metal2 s 117318 139200 117374 140000 6 io_out[26]
port 156 nsew signal output
rlabel metal2 s 121734 139200 121790 140000 6 io_out[27]
port 157 nsew signal output
rlabel metal2 s 126150 139200 126206 140000 6 io_out[28]
port 158 nsew signal output
rlabel metal2 s 130566 139200 130622 140000 6 io_out[29]
port 159 nsew signal output
rlabel metal2 s 11978 139200 12034 140000 6 io_out[2]
port 160 nsew signal output
rlabel metal2 s 134890 139200 134946 140000 6 io_out[30]
port 161 nsew signal output
rlabel metal2 s 139306 139200 139362 140000 6 io_out[31]
port 162 nsew signal output
rlabel metal2 s 143722 139200 143778 140000 6 io_out[32]
port 163 nsew signal output
rlabel metal2 s 148138 139200 148194 140000 6 io_out[33]
port 164 nsew signal output
rlabel metal2 s 152462 139200 152518 140000 6 io_out[34]
port 165 nsew signal output
rlabel metal2 s 156878 139200 156934 140000 6 io_out[35]
port 166 nsew signal output
rlabel metal2 s 161294 139200 161350 140000 6 io_out[36]
port 167 nsew signal output
rlabel metal2 s 165618 139200 165674 140000 6 io_out[37]
port 168 nsew signal output
rlabel metal2 s 16394 139200 16450 140000 6 io_out[3]
port 169 nsew signal output
rlabel metal2 s 20718 139200 20774 140000 6 io_out[4]
port 170 nsew signal output
rlabel metal2 s 25134 139200 25190 140000 6 io_out[5]
port 171 nsew signal output
rlabel metal2 s 29550 139200 29606 140000 6 io_out[6]
port 172 nsew signal output
rlabel metal2 s 33874 139200 33930 140000 6 io_out[7]
port 173 nsew signal output
rlabel metal2 s 38290 139200 38346 140000 6 io_out[8]
port 174 nsew signal output
rlabel metal2 s 42706 139200 42762 140000 6 io_out[9]
port 175 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 mem1_data_i[0]
port 176 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 mem1_data_i[10]
port 177 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 mem1_data_i[11]
port 178 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 mem1_data_i[12]
port 179 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 mem1_data_i[13]
port 180 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 mem1_data_i[14]
port 181 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 mem1_data_i[15]
port 182 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 mem1_data_i[16]
port 183 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 mem1_data_i[17]
port 184 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 mem1_data_i[18]
port 185 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 mem1_data_i[19]
port 186 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 mem1_data_i[1]
port 187 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 mem1_data_i[20]
port 188 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 mem1_data_i[21]
port 189 nsew signal input
rlabel metal3 s 0 105952 800 106072 6 mem1_data_i[22]
port 190 nsew signal input
rlabel metal3 s 0 109488 800 109608 6 mem1_data_i[23]
port 191 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 mem1_data_i[24]
port 192 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 mem1_data_i[25]
port 193 nsew signal input
rlabel metal3 s 0 119824 800 119944 6 mem1_data_i[26]
port 194 nsew signal input
rlabel metal3 s 0 123224 800 123344 6 mem1_data_i[27]
port 195 nsew signal input
rlabel metal3 s 0 126624 800 126744 6 mem1_data_i[28]
port 196 nsew signal input
rlabel metal3 s 0 130160 800 130280 6 mem1_data_i[29]
port 197 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 mem1_data_i[2]
port 198 nsew signal input
rlabel metal3 s 0 133560 800 133680 6 mem1_data_i[30]
port 199 nsew signal input
rlabel metal3 s 0 136960 800 137080 6 mem1_data_i[31]
port 200 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 mem1_data_i[3]
port 201 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 mem1_data_i[4]
port 202 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 mem1_data_i[5]
port 203 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 mem1_data_i[6]
port 204 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 mem1_data_i[7]
port 205 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 mem1_data_i[8]
port 206 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 mem1_data_i[9]
port 207 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 mem_data_i[0]
port 208 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 mem_data_i[10]
port 209 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 mem_data_i[11]
port 210 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 mem_data_i[12]
port 211 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 mem_data_i[13]
port 212 nsew signal input
rlabel metal3 s 0 79568 800 79688 6 mem_data_i[14]
port 213 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 mem_data_i[15]
port 214 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 mem_data_i[16]
port 215 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 mem_data_i[17]
port 216 nsew signal input
rlabel metal3 s 0 93440 800 93560 6 mem_data_i[18]
port 217 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 mem_data_i[19]
port 218 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 mem_data_i[1]
port 219 nsew signal input
rlabel metal3 s 0 100240 800 100360 6 mem_data_i[20]
port 220 nsew signal input
rlabel metal3 s 0 103776 800 103896 6 mem_data_i[21]
port 221 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 mem_data_i[22]
port 222 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 mem_data_i[23]
port 223 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 mem_data_i[24]
port 224 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 mem_data_i[25]
port 225 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 mem_data_i[26]
port 226 nsew signal input
rlabel metal3 s 0 124312 800 124432 6 mem_data_i[27]
port 227 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 mem_data_i[28]
port 228 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 mem_data_i[29]
port 229 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 mem_data_i[2]
port 230 nsew signal input
rlabel metal3 s 0 134648 800 134768 6 mem_data_i[30]
port 231 nsew signal input
rlabel metal3 s 0 138184 800 138304 6 mem_data_i[31]
port 232 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 mem_data_i[3]
port 233 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 mem_data_i[4]
port 234 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 mem_data_i[5]
port 235 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 mem_data_i[6]
port 236 nsew signal input
rlabel metal3 s 0 51008 800 51128 6 mem_data_i[7]
port 237 nsew signal input
rlabel metal3 s 0 56720 800 56840 6 mem_data_i[8]
port 238 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 mem_data_i[9]
port 239 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 mem_data_o[0]
port 240 nsew signal output
rlabel metal3 s 0 67056 800 67176 6 mem_data_o[10]
port 241 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 mem_data_o[11]
port 242 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 mem_data_o[12]
port 243 nsew signal output
rlabel metal3 s 0 77392 800 77512 6 mem_data_o[13]
port 244 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 mem_data_o[14]
port 245 nsew signal output
rlabel metal3 s 0 84192 800 84312 6 mem_data_o[15]
port 246 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 mem_data_o[16]
port 247 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 mem_data_o[17]
port 248 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 mem_data_o[18]
port 249 nsew signal output
rlabel metal3 s 0 97928 800 98048 6 mem_data_o[19]
port 250 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 mem_data_o[1]
port 251 nsew signal output
rlabel metal3 s 0 101464 800 101584 6 mem_data_o[20]
port 252 nsew signal output
rlabel metal3 s 0 104864 800 104984 6 mem_data_o[21]
port 253 nsew signal output
rlabel metal3 s 0 108264 800 108384 6 mem_data_o[22]
port 254 nsew signal output
rlabel metal3 s 0 111800 800 111920 6 mem_data_o[23]
port 255 nsew signal output
rlabel metal3 s 0 115200 800 115320 6 mem_data_o[24]
port 256 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 mem_data_o[25]
port 257 nsew signal output
rlabel metal3 s 0 122136 800 122256 6 mem_data_o[26]
port 258 nsew signal output
rlabel metal3 s 0 125536 800 125656 6 mem_data_o[27]
port 259 nsew signal output
rlabel metal3 s 0 128936 800 129056 6 mem_data_o[28]
port 260 nsew signal output
rlabel metal3 s 0 132336 800 132456 6 mem_data_o[29]
port 261 nsew signal output
rlabel metal3 s 0 23400 800 23520 6 mem_data_o[2]
port 262 nsew signal output
rlabel metal3 s 0 135872 800 135992 6 mem_data_o[30]
port 263 nsew signal output
rlabel metal3 s 0 139272 800 139392 6 mem_data_o[31]
port 264 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 mem_data_o[3]
port 265 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 mem_data_o[4]
port 266 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 mem_data_o[5]
port 267 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 mem_data_o[6]
port 268 nsew signal output
rlabel metal3 s 0 52096 800 52216 6 mem_data_o[7]
port 269 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 mem_data_o[8]
port 270 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 mem_data_o[9]
port 271 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 mem_raddr_o[0]
port 272 nsew signal output
rlabel metal3 s 0 16600 800 16720 6 mem_raddr_o[1]
port 273 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 mem_raddr_o[2]
port 274 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 mem_raddr_o[3]
port 275 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 mem_raddr_o[4]
port 276 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 mem_raddr_o[5]
port 277 nsew signal output
rlabel metal3 s 0 47472 800 47592 6 mem_raddr_o[6]
port 278 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 mem_raddr_o[7]
port 279 nsew signal output
rlabel metal3 s 0 59032 800 59152 6 mem_raddr_o[8]
port 280 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 mem_renb_o[0]
port 281 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 mem_renb_o[1]
port 282 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 mem_waddr_o[0]
port 283 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 mem_waddr_o[1]
port 284 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 mem_waddr_o[2]
port 285 nsew signal output
rlabel metal3 s 0 31424 800 31544 6 mem_waddr_o[3]
port 286 nsew signal output
rlabel metal3 s 0 37136 800 37256 6 mem_waddr_o[4]
port 287 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 mem_waddr_o[5]
port 288 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 mem_waddr_o[6]
port 289 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 mem_waddr_o[7]
port 290 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 mem_waddr_o[8]
port 291 nsew signal output
rlabel metal3 s 0 11976 800 12096 6 mem_wenb_o[0]
port 292 nsew signal output
rlabel metal3 s 0 20000 800 20120 6 mem_wenb_o[1]
port 293 nsew signal output
rlabel metal3 s 179200 127576 180000 127696 6 oversample_o[0]
port 294 nsew signal output
rlabel metal3 s 179200 128936 180000 129056 6 oversample_o[1]
port 295 nsew signal output
rlabel metal3 s 179200 130160 180000 130280 6 oversample_o[2]
port 296 nsew signal output
rlabel metal3 s 179200 131384 180000 131504 6 oversample_o[3]
port 297 nsew signal output
rlabel metal3 s 179200 132744 180000 132864 6 oversample_o[4]
port 298 nsew signal output
rlabel metal3 s 179200 133968 180000 134088 6 oversample_o[5]
port 299 nsew signal output
rlabel metal3 s 179200 135328 180000 135448 6 oversample_o[6]
port 300 nsew signal output
rlabel metal3 s 179200 136552 180000 136672 6 oversample_o[7]
port 301 nsew signal output
rlabel metal3 s 179200 137912 180000 138032 6 oversample_o[8]
port 302 nsew signal output
rlabel metal3 s 179200 139136 180000 139256 6 oversample_o[9]
port 303 nsew signal output
rlabel metal2 s 174450 139200 174506 140000 6 sinc3_en_o[0]
port 304 nsew signal output
rlabel metal2 s 176658 139200 176714 140000 6 sinc3_en_o[1]
port 305 nsew signal output
rlabel metal2 s 178866 139200 178922 140000 6 sinc3_en_o[2]
port 306 nsew signal output
rlabel metal2 s 167826 139200 167882 140000 6 vco_enb_o[0]
port 307 nsew signal output
rlabel metal2 s 170034 139200 170090 140000 6 vco_enb_o[1]
port 308 nsew signal output
rlabel metal2 s 172242 139200 172298 140000 6 vco_enb_o[2]
port 309 nsew signal output
rlabel metal2 s 846 0 902 800 6 wb_clk_i
port 310 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wb_rst_i
port 311 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_ack_o
port 312 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[0]
port 313 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 wbs_adr_i[10]
port 314 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 wbs_adr_i[11]
port 315 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_adr_i[12]
port 316 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_adr_i[13]
port 317 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[14]
port 318 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 wbs_adr_i[15]
port 319 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 wbs_adr_i[16]
port 320 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_adr_i[17]
port 321 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 wbs_adr_i[18]
port 322 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 wbs_adr_i[19]
port 323 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[1]
port 324 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 wbs_adr_i[20]
port 325 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 wbs_adr_i[21]
port 326 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 wbs_adr_i[22]
port 327 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 wbs_adr_i[23]
port 328 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 wbs_adr_i[24]
port 329 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 wbs_adr_i[25]
port 330 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 wbs_adr_i[26]
port 331 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 wbs_adr_i[27]
port 332 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 wbs_adr_i[28]
port 333 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 wbs_adr_i[29]
port 334 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[2]
port 335 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 wbs_adr_i[30]
port 336 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 wbs_adr_i[31]
port 337 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[3]
port 338 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[4]
port 339 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_adr_i[5]
port 340 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[6]
port 341 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_adr_i[7]
port 342 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_adr_i[8]
port 343 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 wbs_adr_i[9]
port 344 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_cyc_i
port 345 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[0]
port 346 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wbs_dat_i[10]
port 347 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_i[11]
port 348 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_i[12]
port 349 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_i[13]
port 350 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_i[14]
port 351 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 wbs_dat_i[15]
port 352 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 wbs_dat_i[16]
port 353 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 wbs_dat_i[17]
port 354 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 wbs_dat_i[18]
port 355 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 wbs_dat_i[19]
port 356 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[1]
port 357 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 wbs_dat_i[20]
port 358 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_i[21]
port 359 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 wbs_dat_i[22]
port 360 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 wbs_dat_i[23]
port 361 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 wbs_dat_i[24]
port 362 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 wbs_dat_i[25]
port 363 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 wbs_dat_i[26]
port 364 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 wbs_dat_i[27]
port 365 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 wbs_dat_i[28]
port 366 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 wbs_dat_i[29]
port 367 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[2]
port 368 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 wbs_dat_i[30]
port 369 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 wbs_dat_i[31]
port 370 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[3]
port 371 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_i[4]
port 372 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_i[5]
port 373 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_i[6]
port 374 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[7]
port 375 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 wbs_dat_i[8]
port 376 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[9]
port 377 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[0]
port 378 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[10]
port 379 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 wbs_dat_o[11]
port 380 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_o[12]
port 381 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_o[13]
port 382 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_o[14]
port 383 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 wbs_dat_o[15]
port 384 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 wbs_dat_o[16]
port 385 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 wbs_dat_o[17]
port 386 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 wbs_dat_o[18]
port 387 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 wbs_dat_o[19]
port 388 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[1]
port 389 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 wbs_dat_o[20]
port 390 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 wbs_dat_o[21]
port 391 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 wbs_dat_o[22]
port 392 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 wbs_dat_o[23]
port 393 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 wbs_dat_o[24]
port 394 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 wbs_dat_o[25]
port 395 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 wbs_dat_o[26]
port 396 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 wbs_dat_o[27]
port 397 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 wbs_dat_o[28]
port 398 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 wbs_dat_o[29]
port 399 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[2]
port 400 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 wbs_dat_o[30]
port 401 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 wbs_dat_o[31]
port 402 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_o[3]
port 403 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[4]
port 404 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[5]
port 405 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[6]
port 406 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[7]
port 407 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_o[8]
port 408 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 wbs_dat_o[9]
port 409 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_sel_i[0]
port 410 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_sel_i[1]
port 411 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_sel_i[2]
port 412 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_sel_i[3]
port 413 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_stb_i
port 414 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_we_i
port 415 nsew signal input
rlabel metal3 s 0 552 800 672 6 wmask_o[0]
port 416 nsew signal output
rlabel metal3 s 0 1640 800 1760 6 wmask_o[1]
port 417 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 wmask_o[2]
port 418 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 wmask_o[3]
port 419 nsew signal output
rlabel metal4 s 157808 2128 158128 137680 6 vccd1
port 420 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 421 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 422 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 423 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 424 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 425 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 137680 6 vssd1
port 426 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 137680 6 vssd1
port 427 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 428 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 429 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 430 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 431 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 137632 6 vccd2
port 432 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 137632 6 vccd2
port 433 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 137632 6 vccd2
port 434 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 137632 6 vccd2
port 435 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 137632 6 vccd2
port 436 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 137632 6 vccd2
port 437 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 137632 6 vssd2
port 438 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 137632 6 vssd2
port 439 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 137632 6 vssd2
port 440 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 137632 6 vssd2
port 441 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 137632 6 vssd2
port 442 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 137632 6 vssd2
port 443 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 137632 6 vdda1
port 444 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 137632 6 vdda1
port 445 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 137632 6 vdda1
port 446 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 137632 6 vdda1
port 447 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 137632 6 vdda1
port 448 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 137632 6 vdda1
port 449 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 137632 6 vssa1
port 450 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 137632 6 vssa1
port 451 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 137632 6 vssa1
port 452 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 137632 6 vssa1
port 453 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 137632 6 vssa1
port 454 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 137632 6 vssa1
port 455 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 137632 6 vdda2
port 456 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 137632 6 vdda2
port 457 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 137632 6 vdda2
port 458 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 137632 6 vdda2
port 459 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 137632 6 vdda2
port 460 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 137632 6 vdda2
port 461 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 137632 6 vssa2
port 462 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 137632 6 vssa2
port 463 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 137632 6 vssa2
port 464 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 137632 6 vssa2
port 465 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 137632 6 vssa2
port 466 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 137632 6 vssa2
port 467 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 140000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 10066530
string GDS_START 602518
<< end >>

