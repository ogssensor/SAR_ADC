magic
tech sky130A
timestamp 1622045257
<< metal1 >>
rect 19800 8413 20000 8461
rect 9000 8141 9200 8189
rect 10800 8141 11000 8189
rect 12600 8141 12800 8189
rect 16200 8141 16400 8189
rect 23400 8141 23600 8189
rect 22996 7325 25424 7373
rect 9000 7053 9200 7101
rect 10800 7053 11000 7101
rect 12600 7053 12800 7101
rect 19800 7053 20000 7101
rect 23400 6780 23600 6828
rect 23400 6237 23600 6285
rect 9000 5965 9200 6013
rect 10800 5965 11000 6013
rect 12600 5965 12800 6013
rect 16200 5965 16400 6013
rect 19800 5965 20000 6013
rect 9000 4877 9200 4925
rect 10800 4877 11000 4925
rect 12600 4877 12800 4925
rect 19800 4877 20000 4925
rect 23400 4877 23600 4925
<< metal2 >>
rect 11833 8466 11913 8566
rect 14783 8466 14863 8566
rect 17733 8466 17813 8566
rect 20683 8466 20763 8566
rect 19800 8413 20000 8461
rect 9000 8141 9200 8189
rect 10800 8141 11000 8189
rect 12600 8141 12800 8189
rect 16200 8141 16400 8189
rect 23400 8141 23600 8189
rect 25200 7325 25400 7373
rect 25201 7168 25301 7248
rect 9000 7053 9200 7101
rect 10800 7053 11000 7101
rect 12600 7053 12800 7101
rect 19800 7053 20000 7101
rect 23400 6780 23600 6828
rect 23400 6237 23600 6285
rect 9000 5965 9200 6013
rect 10800 5965 11000 6013
rect 12600 5965 12800 6013
rect 16200 5965 16400 6013
rect 19800 5965 20000 6013
rect 9000 4877 9200 4925
rect 10800 4877 11000 4925
rect 12600 4877 12800 4925
rect 19800 4877 20000 4925
rect 23400 4877 23600 4925
rect 8478 4500 8558 4600
rect 10278 4500 10358 4600
rect 13228 4500 13308 4600
rect 16178 4500 16258 4600
rect 19128 4500 19208 4600
rect 22078 4500 22158 4600
rect 23787 4500 23867 4600
<< metal3 >>
rect 19800 8455 20000 8461
rect 19800 8419 19816 8455
rect 19852 8419 19860 8455
rect 19896 8419 19904 8455
rect 19940 8419 19948 8455
rect 19984 8419 20000 8455
rect 19800 8413 20000 8419
rect 9000 8183 9200 8189
rect 9000 8147 9016 8183
rect 9052 8147 9060 8183
rect 9096 8147 9104 8183
rect 9140 8147 9148 8183
rect 9184 8147 9200 8183
rect 9000 8141 9200 8147
rect 10800 8183 11000 8189
rect 10800 8147 10816 8183
rect 10852 8147 10860 8183
rect 10896 8147 10904 8183
rect 10940 8147 10948 8183
rect 10984 8147 11000 8183
rect 10800 8141 11000 8147
rect 12600 8183 12800 8189
rect 12600 8147 12616 8183
rect 12652 8147 12660 8183
rect 12696 8147 12704 8183
rect 12740 8147 12748 8183
rect 12784 8147 12800 8183
rect 12600 8141 12800 8147
rect 16200 8183 16400 8189
rect 16200 8147 16216 8183
rect 16252 8147 16260 8183
rect 16296 8147 16304 8183
rect 16340 8147 16348 8183
rect 16384 8147 16400 8183
rect 16200 8141 16400 8147
rect 23400 8183 23600 8189
rect 23400 8147 23416 8183
rect 23452 8147 23460 8183
rect 23496 8147 23504 8183
rect 23540 8147 23548 8183
rect 23584 8147 23600 8183
rect 23400 8141 23600 8147
rect 25200 7367 25400 7373
rect 25200 7331 25216 7367
rect 25252 7331 25260 7367
rect 25296 7331 25304 7367
rect 25340 7331 25348 7367
rect 25384 7331 25400 7367
rect 25200 7325 25400 7331
rect 9000 7095 9200 7101
rect 9000 7059 9016 7095
rect 9052 7059 9060 7095
rect 9096 7059 9104 7095
rect 9140 7059 9148 7095
rect 9184 7059 9200 7095
rect 9000 7053 9200 7059
rect 10800 7095 11000 7101
rect 10800 7059 10816 7095
rect 10852 7059 10860 7095
rect 10896 7059 10904 7095
rect 10940 7059 10948 7095
rect 10984 7059 11000 7095
rect 10800 7053 11000 7059
rect 12600 7095 12800 7101
rect 12600 7059 12616 7095
rect 12652 7059 12660 7095
rect 12696 7059 12704 7095
rect 12740 7059 12748 7095
rect 12784 7059 12800 7095
rect 12600 7053 12800 7059
rect 19800 7095 20000 7101
rect 19800 7059 19816 7095
rect 19852 7059 19860 7095
rect 19896 7059 19904 7095
rect 19940 7059 19948 7095
rect 19984 7059 20000 7095
rect 19800 7053 20000 7059
rect 23400 6822 23600 6828
rect 23400 6786 23416 6822
rect 23452 6786 23460 6822
rect 23496 6786 23504 6822
rect 23540 6786 23548 6822
rect 23584 6786 23600 6822
rect 23400 6780 23600 6786
rect 23400 6279 23600 6285
rect 23400 6243 23416 6279
rect 23452 6243 23460 6279
rect 23496 6243 23504 6279
rect 23540 6243 23548 6279
rect 23584 6243 23600 6279
rect 23400 6237 23600 6243
rect 9000 6007 9200 6013
rect 9000 5971 9016 6007
rect 9052 5971 9060 6007
rect 9096 5971 9104 6007
rect 9140 5971 9148 6007
rect 9184 5971 9200 6007
rect 9000 5965 9200 5971
rect 10800 6007 11000 6013
rect 10800 5971 10816 6007
rect 10852 5971 10860 6007
rect 10896 5971 10904 6007
rect 10940 5971 10948 6007
rect 10984 5971 11000 6007
rect 10800 5965 11000 5971
rect 12600 6007 12800 6013
rect 12600 5971 12616 6007
rect 12652 5971 12660 6007
rect 12696 5971 12704 6007
rect 12740 5971 12748 6007
rect 12784 5971 12800 6007
rect 12600 5965 12800 5971
rect 16200 6007 16400 6013
rect 16200 5971 16216 6007
rect 16252 5971 16260 6007
rect 16296 5971 16304 6007
rect 16340 5971 16348 6007
rect 16384 5971 16400 6007
rect 16200 5965 16400 5971
rect 19800 6007 20000 6013
rect 19800 5971 19816 6007
rect 19852 5971 19860 6007
rect 19896 5971 19904 6007
rect 19940 5971 19948 6007
rect 19984 5971 20000 6007
rect 19800 5965 20000 5971
rect 9000 4919 9200 4925
rect 9000 4883 9016 4919
rect 9052 4883 9060 4919
rect 9096 4883 9104 4919
rect 9140 4883 9148 4919
rect 9184 4883 9200 4919
rect 9000 4877 9200 4883
rect 10800 4919 11000 4925
rect 10800 4883 10816 4919
rect 10852 4883 10860 4919
rect 10896 4883 10904 4919
rect 10940 4883 10948 4919
rect 10984 4883 11000 4919
rect 10800 4877 11000 4883
rect 12600 4919 12800 4925
rect 12600 4883 12616 4919
rect 12652 4883 12660 4919
rect 12696 4883 12704 4919
rect 12740 4883 12748 4919
rect 12784 4883 12800 4919
rect 12600 4877 12800 4883
rect 19800 4919 20000 4925
rect 19800 4883 19816 4919
rect 19852 4883 19860 4919
rect 19896 4883 19904 4919
rect 19940 4883 19948 4919
rect 19984 4883 20000 4919
rect 19800 4877 20000 4883
rect 23400 4919 23600 4925
rect 23400 4883 23416 4919
rect 23452 4883 23460 4919
rect 23496 4883 23504 4919
rect 23540 4883 23548 4919
rect 23584 4883 23600 4919
rect 23400 4877 23600 4883
<< via3 >>
rect 19816 8419 19852 8455
rect 19860 8419 19896 8455
rect 19904 8419 19940 8455
rect 19948 8419 19984 8455
rect 9016 8147 9052 8183
rect 9060 8147 9096 8183
rect 9104 8147 9140 8183
rect 9148 8147 9184 8183
rect 10816 8147 10852 8183
rect 10860 8147 10896 8183
rect 10904 8147 10940 8183
rect 10948 8147 10984 8183
rect 12616 8147 12652 8183
rect 12660 8147 12696 8183
rect 12704 8147 12740 8183
rect 12748 8147 12784 8183
rect 16216 8147 16252 8183
rect 16260 8147 16296 8183
rect 16304 8147 16340 8183
rect 16348 8147 16384 8183
rect 23416 8147 23452 8183
rect 23460 8147 23496 8183
rect 23504 8147 23540 8183
rect 23548 8147 23584 8183
rect 25216 7331 25252 7367
rect 25260 7331 25296 7367
rect 25304 7331 25340 7367
rect 25348 7331 25384 7367
rect 9016 7059 9052 7095
rect 9060 7059 9096 7095
rect 9104 7059 9140 7095
rect 9148 7059 9184 7095
rect 10816 7059 10852 7095
rect 10860 7059 10896 7095
rect 10904 7059 10940 7095
rect 10948 7059 10984 7095
rect 12616 7059 12652 7095
rect 12660 7059 12696 7095
rect 12704 7059 12740 7095
rect 12748 7059 12784 7095
rect 19816 7059 19852 7095
rect 19860 7059 19896 7095
rect 19904 7059 19940 7095
rect 19948 7059 19984 7095
rect 23416 6786 23452 6822
rect 23460 6786 23496 6822
rect 23504 6786 23540 6822
rect 23548 6786 23584 6822
rect 23416 6243 23452 6279
rect 23460 6243 23496 6279
rect 23504 6243 23540 6279
rect 23548 6243 23584 6279
rect 9016 5971 9052 6007
rect 9060 5971 9096 6007
rect 9104 5971 9140 6007
rect 9148 5971 9184 6007
rect 10816 5971 10852 6007
rect 10860 5971 10896 6007
rect 10904 5971 10940 6007
rect 10948 5971 10984 6007
rect 12616 5971 12652 6007
rect 12660 5971 12696 6007
rect 12704 5971 12740 6007
rect 12748 5971 12784 6007
rect 16216 5971 16252 6007
rect 16260 5971 16296 6007
rect 16304 5971 16340 6007
rect 16348 5971 16384 6007
rect 19816 5971 19852 6007
rect 19860 5971 19896 6007
rect 19904 5971 19940 6007
rect 19948 5971 19984 6007
rect 9016 4883 9052 4919
rect 9060 4883 9096 4919
rect 9104 4883 9140 4919
rect 9148 4883 9184 4919
rect 10816 4883 10852 4919
rect 10860 4883 10896 4919
rect 10904 4883 10940 4919
rect 10948 4883 10984 4919
rect 12616 4883 12652 4919
rect 12660 4883 12696 4919
rect 12704 4883 12740 4919
rect 12748 4883 12784 4919
rect 19816 4883 19852 4919
rect 19860 4883 19896 4919
rect 19904 4883 19940 4919
rect 19948 4883 19984 4919
rect 23416 4883 23452 4919
rect 23460 4883 23496 4919
rect 23504 4883 23540 4919
rect 23548 4883 23584 4919
<< metal4 >>
rect 19800 8455 20000 8461
rect 19800 8419 19816 8455
rect 19852 8419 19860 8455
rect 19896 8419 19904 8455
rect 19940 8419 19948 8455
rect 19984 8419 20000 8455
rect 19800 8413 20000 8419
rect 9000 8183 9200 8189
rect 9000 8147 9016 8183
rect 9052 8147 9060 8183
rect 9096 8147 9104 8183
rect 9140 8147 9148 8183
rect 9184 8147 9200 8183
rect 9000 8141 9200 8147
rect 10800 8183 11000 8189
rect 10800 8147 10816 8183
rect 10852 8147 10860 8183
rect 10896 8147 10904 8183
rect 10940 8147 10948 8183
rect 10984 8147 11000 8183
rect 10800 8141 11000 8147
rect 12600 8183 12800 8189
rect 12600 8147 12616 8183
rect 12652 8147 12660 8183
rect 12696 8147 12704 8183
rect 12740 8147 12748 8183
rect 12784 8147 12800 8183
rect 12600 8141 12800 8147
rect 16200 8183 16400 8189
rect 16200 8147 16216 8183
rect 16252 8147 16260 8183
rect 16296 8147 16304 8183
rect 16340 8147 16348 8183
rect 16384 8147 16400 8183
rect 16200 8141 16400 8147
rect 23400 8183 23600 8189
rect 23400 8147 23416 8183
rect 23452 8147 23460 8183
rect 23496 8147 23504 8183
rect 23540 8147 23548 8183
rect 23584 8147 23600 8183
rect 23400 8141 23600 8147
rect 25200 7367 25400 7373
rect 25200 7331 25216 7367
rect 25252 7331 25260 7367
rect 25296 7331 25304 7367
rect 25340 7331 25348 7367
rect 25384 7331 25400 7367
rect 25200 7325 25400 7331
rect 9000 7095 9200 7101
rect 9000 7059 9016 7095
rect 9052 7059 9060 7095
rect 9096 7059 9104 7095
rect 9140 7059 9148 7095
rect 9184 7059 9200 7095
rect 9000 7053 9200 7059
rect 10800 7095 11000 7101
rect 10800 7059 10816 7095
rect 10852 7059 10860 7095
rect 10896 7059 10904 7095
rect 10940 7059 10948 7095
rect 10984 7059 11000 7095
rect 10800 7053 11000 7059
rect 12600 7095 12800 7101
rect 12600 7059 12616 7095
rect 12652 7059 12660 7095
rect 12696 7059 12704 7095
rect 12740 7059 12748 7095
rect 12784 7059 12800 7095
rect 12600 7053 12800 7059
rect 19800 7095 20000 7101
rect 19800 7059 19816 7095
rect 19852 7059 19860 7095
rect 19896 7059 19904 7095
rect 19940 7059 19948 7095
rect 19984 7059 20000 7095
rect 19800 7053 20000 7059
rect 23400 6822 23600 6828
rect 23400 6786 23416 6822
rect 23452 6786 23460 6822
rect 23496 6786 23504 6822
rect 23540 6786 23548 6822
rect 23584 6786 23600 6822
rect 23400 6780 23600 6786
rect 23400 6279 23600 6285
rect 23400 6243 23416 6279
rect 23452 6243 23460 6279
rect 23496 6243 23504 6279
rect 23540 6243 23548 6279
rect 23584 6243 23600 6279
rect 23400 6237 23600 6243
rect 9000 6007 9200 6013
rect 9000 5971 9016 6007
rect 9052 5971 9060 6007
rect 9096 5971 9104 6007
rect 9140 5971 9148 6007
rect 9184 5971 9200 6007
rect 9000 5965 9200 5971
rect 10800 6007 11000 6013
rect 10800 5971 10816 6007
rect 10852 5971 10860 6007
rect 10896 5971 10904 6007
rect 10940 5971 10948 6007
rect 10984 5971 11000 6007
rect 10800 5965 11000 5971
rect 12600 6007 12800 6013
rect 12600 5971 12616 6007
rect 12652 5971 12660 6007
rect 12696 5971 12704 6007
rect 12740 5971 12748 6007
rect 12784 5971 12800 6007
rect 12600 5965 12800 5971
rect 16200 6007 16400 6013
rect 16200 5971 16216 6007
rect 16252 5971 16260 6007
rect 16296 5971 16304 6007
rect 16340 5971 16348 6007
rect 16384 5971 16400 6007
rect 16200 5965 16400 5971
rect 19800 6007 20000 6013
rect 19800 5971 19816 6007
rect 19852 5971 19860 6007
rect 19896 5971 19904 6007
rect 19940 5971 19948 6007
rect 19984 5971 20000 6007
rect 19800 5965 20000 5971
rect 9000 4919 9200 4925
rect 9000 4883 9016 4919
rect 9052 4883 9060 4919
rect 9096 4883 9104 4919
rect 9140 4883 9148 4919
rect 9184 4883 9200 4919
rect 9000 4877 9200 4883
rect 10800 4919 11000 4925
rect 10800 4883 10816 4919
rect 10852 4883 10860 4919
rect 10896 4883 10904 4919
rect 10940 4883 10948 4919
rect 10984 4883 11000 4919
rect 10800 4877 11000 4883
rect 12600 4919 12800 4925
rect 12600 4883 12616 4919
rect 12652 4883 12660 4919
rect 12696 4883 12704 4919
rect 12740 4883 12748 4919
rect 12784 4883 12800 4919
rect 12600 4877 12800 4883
rect 19800 4919 20000 4925
rect 19800 4883 19816 4919
rect 19852 4883 19860 4919
rect 19896 4883 19904 4919
rect 19940 4883 19948 4919
rect 19984 4883 20000 4919
rect 19800 4877 20000 4883
rect 23400 4919 23600 4925
rect 23400 4883 23416 4919
rect 23452 4883 23460 4919
rect 23496 4883 23504 4919
rect 23540 4883 23548 4919
rect 23584 4883 23600 4919
rect 23400 4877 23600 4883
<< metal5 >>
rect 28000 13100 28500 13300
rect 27500 12600 28000 12800
use power_ring  power_ring_0
timestamp 1622042232
transform 1 0 -6300 0 1 2400
box 6300 -2400 35400 10900
use ring_osc_3-1  ring_osc_3-1_0
timestamp 1622022171
transform 1 0 7151 0 1 4629
box 0 -129 18150 3937
<< labels >>
flabel metal5 s 28000 13100 28500 13300 1 FreeSans 1200 0 0 0 vccd1
port 13 nsew power bidirectional abutment
flabel metal5 s 27500 12600 28000 12800 1 FreeSans 1200 0 0 0 vssd1
port 14 nsew ground bidirectional abutment
flabel metal2 25201 7168 25301 7248 1 FreeSans 1 0 0 0 input_analog
port 12 nsew signal input
flabel metal2 22078 4500 22158 4600 1 FreeSans 1 0 0 0 p[0]
port 1 nsew signal output
flabel metal2 19128 4500 19208 4600 1 FreeSans 1 0 0 0 p[1]
port 2 nsew signal output
flabel metal2 16178 4500 16258 4600 1 FreeSans 1 0 0 0 p[2]
port 3 nsew signal output
flabel metal2 13228 4500 13308 4600 1 FreeSans 1 0 0 0 p[3]
port 4 nsew signal output
flabel metal2 10278 4500 10358 4600 1 FreeSans 1 0 0 0 p[4]
port 5 nsew signal output
flabel metal2 8478 4500 8558 4600 1 FreeSans 1 0 0 0 p[5]
port 6 nsew signal output
flabel metal2 11833 8466 11913 8566 1 FreeSans 1 0 0 0 p[6]
port 7 nsew signal output
flabel metal2 14783 8466 14863 8566 1 FreeSans 1 0 0 0 p[7]
port 8 nsew signal output
flabel metal2 17733 8466 17813 8566 1 FreeSans 1 0 0 0 p[8]
port 9 nsew signal output
flabel metal2 20683 8466 20763 8566 1 FreeSans 1 0 0 0 p[9]
port 10 nsew signal output
flabel metal2 23787 4500 23867 4600 1 FreeSans 1 0 0 0 p[10]
port 11 nsew signal output
<< end >>
