MACRO vco_r100
  CLASS BLOCK ;
  FOREIGN vco_r100 ;
  ORIGIN 0.000 0.000 ;
  SIZE 183.510 BY 105.000 ;
  PIN p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.680500 ;
    PORT
      LAYER met2 ;
        RECT 16.630 61.510 18.375 62.210 ;
        RECT 16.630 50.650 17.330 61.510 ;
        RECT 6.215 49.950 17.330 50.650 ;
        RECT 6.215 43.010 6.915 49.950 ;
        RECT 6.140 42.550 7.060 43.010 ;
        RECT 6.215 42.470 6.915 42.550 ;
    END
  END p[0]
  PIN p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 30.590 42.550 31.510 43.010 ;
    END
  END p[1]
  PIN p[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 46.230 61.630 47.150 62.090 ;
    END
  END p[2]
  PIN p[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 60.030 42.550 60.950 43.010 ;
    END
  END p[3]
  PIN p[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 75.670 61.630 76.590 62.090 ;
    END
  END p[4]
  PIN p[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 89.470 42.550 90.390 43.010 ;
    END
  END p[5]
  PIN p[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 105.110 61.630 106.030 62.090 ;
    END
  END p[6]
  PIN p[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 119.370 42.550 120.290 43.010 ;
    END
  END p[7]
  PIN p[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 134.550 61.630 135.470 62.090 ;
    END
  END p[8]
  PIN p[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 148.810 42.550 149.730 43.010 ;
    END
  END p[9]
  PIN p[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 70.199997 ;
    ANTENNADIFFAREA 6.235000 ;
    PORT
      LAYER met2 ;
        RECT 163.960 61.510 166.300 62.210 ;
        RECT 165.600 43.170 166.300 61.510 ;
        RECT 165.600 42.440 166.970 43.170 ;
    END
  END p[10]
  PIN input_analog
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.080 58.690 183.510 59.490 ;
    END
  END input_analog
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER nwell ;
        RECT 3.140 61.805 5.820 63.640 ;
        RECT 7.310 61.805 9.070 63.640 ;
        RECT 17.900 57.545 23.750 63.420 ;
        RECT 28.730 63.080 34.580 68.935 ;
        RECT 42.350 63.610 46.110 68.885 ;
        RECT 35.875 57.550 39.635 62.860 ;
        RECT 47.400 57.545 53.250 63.420 ;
        RECT 58.230 63.080 64.080 68.935 ;
        RECT 71.850 63.610 75.610 68.885 ;
        RECT 65.375 57.550 69.135 62.860 ;
        RECT 76.900 57.545 82.750 63.420 ;
        RECT 87.730 63.080 93.580 68.935 ;
        RECT 101.350 63.610 105.110 68.885 ;
        RECT 94.875 57.550 98.635 62.860 ;
        RECT 106.400 57.545 112.250 63.420 ;
        RECT 117.230 63.080 123.080 68.935 ;
        RECT 130.850 63.610 134.610 68.885 ;
        RECT 124.375 57.550 128.135 62.860 ;
        RECT 135.900 57.545 141.750 63.420 ;
        RECT 146.730 63.080 152.580 68.935 ;
        RECT 160.350 63.610 164.110 68.885 ;
        RECT 153.875 57.550 157.635 62.860 ;
        RECT 8.775 41.820 12.535 47.130 ;
        RECT 2.300 35.795 6.060 41.070 ;
        RECT 13.830 35.745 19.680 41.600 ;
        RECT 24.660 41.260 30.510 47.135 ;
        RECT 38.275 41.820 42.035 47.130 ;
        RECT 31.800 35.795 35.560 41.070 ;
        RECT 43.330 35.745 49.180 41.600 ;
        RECT 54.160 41.260 60.010 47.135 ;
        RECT 67.775 41.820 71.535 47.130 ;
        RECT 61.300 35.795 65.060 41.070 ;
        RECT 72.830 35.745 78.680 41.600 ;
        RECT 83.660 41.260 89.510 47.135 ;
        RECT 97.275 41.820 101.035 47.130 ;
        RECT 90.800 35.795 94.560 41.070 ;
        RECT 102.330 35.745 108.180 41.600 ;
        RECT 113.160 41.260 119.010 47.135 ;
        RECT 126.775 41.820 130.535 47.130 ;
        RECT 120.300 35.795 124.060 41.070 ;
        RECT 131.830 35.745 137.680 41.600 ;
        RECT 142.660 41.260 148.510 47.135 ;
        RECT 156.275 41.820 160.035 47.130 ;
        RECT 149.800 35.795 153.560 41.070 ;
        RECT 161.330 35.745 167.180 41.600 ;
        RECT 172.160 41.260 178.010 47.135 ;
      LAYER met4 ;
        RECT 5.000 0.000 7.000 105.000 ;
        RECT 18.000 0.000 20.000 105.000 ;
        RECT 54.000 0.000 56.000 105.000 ;
        RECT 90.000 0.000 92.000 105.000 ;
        RECT 126.000 0.000 128.000 105.000 ;
        RECT 162.000 0.000 164.000 105.000 ;
        RECT 175.000 0.000 177.000 105.000 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met4 ;
        RECT 0.000 4.000 2.000 101.000 ;
        RECT 36.000 4.000 38.000 101.000 ;
        RECT 72.000 4.000 74.000 101.000 ;
        RECT 108.000 4.000 110.000 101.000 ;
        RECT 144.000 4.000 146.000 101.000 ;
        RECT 180.000 4.000 182.000 101.000 ;
    END
  END vssd2
  PIN enb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.223500 ;
    PORT
      LAYER met3 ;
        RECT 2.350 61.770 2.710 63.180 ;
    END
  END enb
  OBS
      LAYER pwell ;
        RECT 17.900 65.610 27.930 71.670 ;
        RECT 35.875 65.570 41.725 71.670 ;
        RECT 47.400 65.610 57.430 71.670 ;
        RECT 65.375 65.570 71.225 71.670 ;
        RECT 76.900 65.610 86.930 71.670 ;
        RECT 94.875 65.570 100.725 71.670 ;
        RECT 106.400 65.610 116.430 71.670 ;
        RECT 124.375 65.570 130.225 71.670 ;
        RECT 135.900 65.610 145.930 71.670 ;
        RECT 153.875 65.570 159.725 71.670 ;
        RECT 3.820 61.285 5.625 61.515 ;
        RECT 3.335 60.605 5.625 61.285 ;
        RECT 3.480 60.415 3.650 60.605 ;
        RECT 7.645 60.415 7.815 60.585 ;
        RECT 24.550 54.760 34.580 61.160 ;
        RECT 40.255 59.925 46.105 60.865 ;
        RECT 40.255 59.875 46.110 59.925 ;
        RECT 40.260 54.765 46.110 59.875 ;
        RECT 54.050 54.760 64.080 61.160 ;
        RECT 69.755 59.925 75.605 60.865 ;
        RECT 69.755 59.875 75.610 59.925 ;
        RECT 69.760 54.765 75.610 59.875 ;
        RECT 83.550 54.760 93.580 61.160 ;
        RECT 99.255 59.925 105.105 60.865 ;
        RECT 99.255 59.875 105.110 59.925 ;
        RECT 99.260 54.765 105.110 59.875 ;
        RECT 113.050 54.760 123.080 61.160 ;
        RECT 128.755 59.925 134.605 60.865 ;
        RECT 128.755 59.875 134.610 59.925 ;
        RECT 128.760 54.765 134.610 59.875 ;
        RECT 142.550 54.760 152.580 61.160 ;
        RECT 158.255 59.925 164.105 60.865 ;
        RECT 158.255 59.875 164.110 59.925 ;
        RECT 158.260 54.765 164.110 59.875 ;
        RECT 171.100 53.580 177.890 60.580 ;
        RECT 2.300 44.805 8.150 49.915 ;
        RECT 2.300 44.755 8.155 44.805 ;
        RECT 2.305 43.815 8.155 44.755 ;
        RECT 13.830 43.520 23.860 49.920 ;
        RECT 31.800 44.805 37.650 49.915 ;
        RECT 31.800 44.755 37.655 44.805 ;
        RECT 31.805 43.815 37.655 44.755 ;
        RECT 43.330 43.520 53.360 49.920 ;
        RECT 61.300 44.805 67.150 49.915 ;
        RECT 61.300 44.755 67.155 44.805 ;
        RECT 61.305 43.815 67.155 44.755 ;
        RECT 72.830 43.520 82.860 49.920 ;
        RECT 90.800 44.805 96.650 49.915 ;
        RECT 90.800 44.755 96.655 44.805 ;
        RECT 90.805 43.815 96.655 44.755 ;
        RECT 102.330 43.520 112.360 49.920 ;
        RECT 120.300 44.805 126.150 49.915 ;
        RECT 120.300 44.755 126.155 44.805 ;
        RECT 120.305 43.815 126.155 44.755 ;
        RECT 131.830 43.520 141.860 49.920 ;
        RECT 149.800 44.805 155.650 49.915 ;
        RECT 149.800 44.755 155.655 44.805 ;
        RECT 149.805 43.815 155.655 44.755 ;
        RECT 161.330 43.520 171.360 49.920 ;
        RECT 6.685 33.010 12.535 39.110 ;
        RECT 20.480 33.010 30.510 39.070 ;
        RECT 36.185 33.010 42.035 39.110 ;
        RECT 49.980 33.010 60.010 39.070 ;
        RECT 65.685 33.010 71.535 39.110 ;
        RECT 79.480 33.010 89.510 39.070 ;
        RECT 95.185 33.010 101.035 39.110 ;
        RECT 108.980 33.010 119.010 39.070 ;
        RECT 124.685 33.010 130.535 39.110 ;
        RECT 138.480 33.010 148.510 39.070 ;
        RECT 154.185 33.010 160.035 39.110 ;
        RECT 167.980 33.010 178.010 39.070 ;
      LAYER li1 ;
        RECT 15.430 73.000 166.090 73.500 ;
        RECT 3.850 63.305 4.820 63.460 ;
        RECT 7.850 63.305 8.820 63.460 ;
        RECT 3.330 63.135 5.630 63.305 ;
        RECT 7.500 63.135 8.880 63.305 ;
        RECT 3.415 62.565 3.675 62.965 ;
        RECT 3.845 62.735 4.780 63.135 ;
        RECT 4.950 62.625 5.545 62.965 ;
        RECT 3.415 62.395 4.780 62.565 ;
        RECT 3.415 62.100 3.875 62.225 ;
        RECT 2.380 61.800 3.875 62.100 ;
        RECT 3.415 61.495 3.875 61.800 ;
        RECT 4.045 61.325 4.780 62.395 ;
        RECT 3.415 61.155 4.780 61.325 ;
        RECT 4.950 61.305 5.125 62.625 ;
        RECT 5.840 62.455 7.290 62.675 ;
        RECT 5.305 62.375 7.290 62.455 ;
        RECT 7.775 62.410 8.105 63.135 ;
        RECT 5.305 62.155 6.140 62.375 ;
        RECT 6.990 62.240 7.290 62.375 ;
        RECT 5.305 61.475 5.545 62.155 ;
        RECT 4.950 61.175 5.545 61.305 ;
        RECT 6.370 61.175 6.670 62.010 ;
        RECT 6.990 61.940 8.105 62.240 ;
        RECT 3.415 60.755 3.675 61.155 ;
        RECT 3.845 60.585 4.780 60.985 ;
        RECT 4.950 60.875 6.670 61.175 ;
        RECT 4.950 60.755 5.545 60.875 ;
        RECT 7.585 60.755 8.105 61.940 ;
        RECT 8.275 61.415 8.795 62.965 ;
        RECT 8.275 60.585 8.615 61.245 ;
        RECT 3.330 60.415 5.630 60.585 ;
        RECT 7.500 60.415 8.880 60.585 ;
        RECT 15.510 53.500 16.010 73.000 ;
        RECT 18.080 71.140 20.425 71.620 ;
        RECT 21.490 71.140 24.350 71.620 ;
        RECT 25.405 71.140 27.750 71.620 ;
        RECT 36.055 71.140 38.400 71.620 ;
        RECT 39.200 71.140 41.545 71.620 ;
        RECT 47.580 71.140 49.925 71.620 ;
        RECT 50.990 71.140 53.850 71.620 ;
        RECT 54.905 71.140 57.250 71.620 ;
        RECT 65.555 71.140 67.900 71.620 ;
        RECT 68.700 71.140 71.045 71.620 ;
        RECT 77.080 71.140 79.425 71.620 ;
        RECT 80.490 71.140 83.350 71.620 ;
        RECT 84.405 71.140 86.750 71.620 ;
        RECT 95.055 71.140 97.400 71.620 ;
        RECT 98.200 71.140 100.545 71.620 ;
        RECT 106.580 71.140 108.925 71.620 ;
        RECT 109.990 71.140 112.850 71.620 ;
        RECT 113.905 71.140 116.250 71.620 ;
        RECT 124.555 71.140 126.900 71.620 ;
        RECT 127.700 71.140 130.045 71.620 ;
        RECT 136.080 71.140 138.425 71.620 ;
        RECT 139.490 71.140 142.350 71.620 ;
        RECT 143.405 71.140 145.750 71.620 ;
        RECT 154.055 71.140 156.400 71.620 ;
        RECT 157.200 71.140 159.545 71.620 ;
        RECT 18.590 66.545 18.880 71.140 ;
        RECT 18.650 66.300 18.820 66.545 ;
        RECT 18.800 64.090 19.930 65.090 ;
        RECT 20.680 64.780 20.970 70.840 ;
        RECT 22.770 66.545 23.060 71.140 ;
        RECT 22.830 66.300 23.000 66.545 ;
        RECT 24.860 64.880 25.150 70.840 ;
        RECT 26.950 66.545 27.240 71.140 ;
        RECT 28.910 68.755 31.255 68.900 ;
        RECT 32.055 68.755 34.400 68.900 ;
        RECT 28.910 68.585 34.400 68.755 ;
        RECT 28.910 68.420 31.255 68.585 ;
        RECT 32.055 68.420 34.400 68.585 ;
        RECT 27.010 66.535 27.205 66.545 ;
        RECT 27.010 66.300 27.180 66.535 ;
        RECT 24.860 64.780 25.680 64.880 ;
        RECT 20.680 64.280 25.680 64.780 ;
        RECT 18.080 58.020 18.250 62.875 ;
        RECT 18.590 58.020 18.880 62.870 ;
        RECT 20.680 58.330 20.970 64.280 ;
        RECT 28.910 63.760 29.080 68.420 ;
        RECT 29.420 63.590 29.710 68.420 ;
        RECT 31.510 63.150 31.800 68.150 ;
        RECT 33.600 63.590 33.890 68.420 ;
        RECT 34.230 63.820 34.400 68.420 ;
        RECT 36.565 66.790 36.855 71.140 ;
        RECT 36.800 64.880 38.000 65.190 ;
        RECT 36.300 64.260 38.000 64.880 ;
        RECT 36.800 64.060 38.000 64.260 ;
        RECT 38.650 63.150 38.945 70.830 ;
        RECT 40.745 66.790 41.035 71.140 ;
        RECT 43.835 68.870 45.930 68.900 ;
        RECT 43.680 68.705 45.930 68.870 ;
        RECT 42.530 68.535 45.930 68.705 ;
        RECT 42.530 65.560 42.700 68.535 ;
        RECT 43.680 68.450 45.930 68.535 ;
        RECT 43.835 68.420 45.930 68.450 ;
        RECT 43.035 64.975 43.330 68.050 ;
        RECT 42.805 64.195 43.545 64.975 ;
        RECT 22.770 58.020 23.060 62.870 ;
        RECT 23.400 58.020 23.570 62.875 ;
        RECT 28.870 62.650 41.465 63.150 ;
        RECT 28.870 61.210 29.370 62.650 ;
        RECT 30.400 61.620 34.400 62.220 ;
        RECT 32.400 61.500 34.400 61.620 ;
        RECT 27.330 60.920 31.800 61.210 ;
        RECT 32.400 60.920 33.600 61.500 ;
        RECT 25.300 59.895 25.470 60.130 ;
        RECT 25.275 59.885 25.470 59.895 ;
        RECT 18.080 57.895 20.425 58.020 ;
        RECT 21.225 57.990 23.570 58.020 ;
        RECT 21.225 57.895 23.750 57.990 ;
        RECT 18.080 57.725 23.750 57.895 ;
        RECT 18.080 57.540 20.425 57.725 ;
        RECT 21.225 57.570 23.750 57.725 ;
        RECT 21.225 57.540 23.570 57.570 ;
        RECT 25.240 55.300 25.530 59.885 ;
        RECT 27.330 55.590 27.620 60.920 ;
        RECT 29.480 59.885 29.650 60.110 ;
        RECT 29.420 55.300 29.710 59.885 ;
        RECT 31.510 55.590 31.800 60.920 ;
        RECT 33.660 59.885 33.830 60.110 ;
        RECT 33.600 55.300 33.890 59.885 ;
        RECT 36.055 58.020 36.225 61.945 ;
        RECT 36.565 58.020 36.855 62.090 ;
        RECT 38.655 58.385 38.950 62.650 ;
        RECT 36.055 57.990 38.150 58.020 ;
        RECT 36.055 57.900 38.305 57.990 ;
        RECT 39.285 57.900 39.455 61.935 ;
        RECT 40.965 61.500 41.465 62.650 ;
        RECT 36.055 57.730 39.455 57.900 ;
        RECT 36.055 57.570 38.305 57.730 ;
        RECT 36.055 57.540 38.150 57.570 ;
        RECT 40.950 55.300 41.240 59.645 ;
        RECT 43.035 55.605 43.330 64.195 ;
        RECT 45.130 64.010 45.420 68.420 ;
        RECT 45.760 64.005 45.930 68.420 ;
        RECT 48.090 66.545 48.380 71.140 ;
        RECT 48.150 66.300 48.320 66.545 ;
        RECT 48.300 64.090 49.430 65.090 ;
        RECT 50.180 64.780 50.470 70.840 ;
        RECT 52.270 66.545 52.560 71.140 ;
        RECT 52.330 66.300 52.500 66.545 ;
        RECT 54.360 64.880 54.650 70.840 ;
        RECT 56.450 66.545 56.740 71.140 ;
        RECT 58.410 68.755 60.755 68.900 ;
        RECT 61.555 68.755 63.900 68.900 ;
        RECT 58.410 68.585 63.900 68.755 ;
        RECT 58.410 68.420 60.755 68.585 ;
        RECT 61.555 68.420 63.900 68.585 ;
        RECT 56.510 66.535 56.705 66.545 ;
        RECT 56.510 66.300 56.680 66.535 ;
        RECT 54.360 64.780 55.180 64.880 ;
        RECT 50.180 64.280 55.180 64.780 ;
        RECT 43.950 62.160 45.130 62.360 ;
        RECT 43.950 61.560 45.630 62.160 ;
        RECT 43.950 61.280 45.130 61.560 ;
        RECT 45.130 55.300 45.420 59.645 ;
        RECT 47.580 58.020 47.750 62.875 ;
        RECT 48.090 58.020 48.380 62.870 ;
        RECT 50.180 58.330 50.470 64.280 ;
        RECT 58.410 63.760 58.580 68.420 ;
        RECT 58.920 63.590 59.210 68.420 ;
        RECT 61.010 63.150 61.300 68.150 ;
        RECT 63.100 63.590 63.390 68.420 ;
        RECT 63.730 63.820 63.900 68.420 ;
        RECT 66.065 66.790 66.355 71.140 ;
        RECT 66.300 64.880 67.500 65.190 ;
        RECT 65.800 64.260 67.500 64.880 ;
        RECT 66.300 64.060 67.500 64.260 ;
        RECT 68.150 63.150 68.445 70.830 ;
        RECT 70.245 66.790 70.535 71.140 ;
        RECT 73.335 68.870 75.430 68.900 ;
        RECT 73.180 68.705 75.430 68.870 ;
        RECT 72.030 68.535 75.430 68.705 ;
        RECT 72.030 65.560 72.200 68.535 ;
        RECT 73.180 68.450 75.430 68.535 ;
        RECT 73.335 68.420 75.430 68.450 ;
        RECT 72.535 64.975 72.830 68.050 ;
        RECT 72.305 64.195 73.045 64.975 ;
        RECT 52.270 58.020 52.560 62.870 ;
        RECT 52.900 58.020 53.070 62.875 ;
        RECT 58.370 62.650 70.965 63.150 ;
        RECT 58.370 61.210 58.870 62.650 ;
        RECT 59.900 61.620 63.900 62.220 ;
        RECT 61.900 61.500 63.900 61.620 ;
        RECT 56.830 60.920 61.300 61.210 ;
        RECT 61.900 60.920 63.100 61.500 ;
        RECT 54.800 59.895 54.970 60.130 ;
        RECT 54.775 59.885 54.970 59.895 ;
        RECT 47.580 57.895 49.925 58.020 ;
        RECT 50.725 57.990 53.070 58.020 ;
        RECT 50.725 57.895 53.250 57.990 ;
        RECT 47.580 57.725 53.250 57.895 ;
        RECT 47.580 57.540 49.925 57.725 ;
        RECT 50.725 57.570 53.250 57.725 ;
        RECT 50.725 57.540 53.070 57.570 ;
        RECT 54.740 55.300 55.030 59.885 ;
        RECT 56.830 55.590 57.120 60.920 ;
        RECT 58.980 59.885 59.150 60.110 ;
        RECT 58.920 55.300 59.210 59.885 ;
        RECT 61.010 55.590 61.300 60.920 ;
        RECT 63.160 59.885 63.330 60.110 ;
        RECT 63.100 55.300 63.390 59.885 ;
        RECT 65.555 58.020 65.725 61.945 ;
        RECT 66.065 58.020 66.355 62.090 ;
        RECT 68.155 58.385 68.450 62.650 ;
        RECT 65.555 57.990 67.650 58.020 ;
        RECT 65.555 57.900 67.805 57.990 ;
        RECT 68.785 57.900 68.955 61.935 ;
        RECT 70.465 61.500 70.965 62.650 ;
        RECT 65.555 57.730 68.955 57.900 ;
        RECT 65.555 57.570 67.805 57.730 ;
        RECT 65.555 57.540 67.650 57.570 ;
        RECT 70.450 55.300 70.740 59.645 ;
        RECT 72.535 55.605 72.830 64.195 ;
        RECT 74.630 64.010 74.920 68.420 ;
        RECT 75.260 64.005 75.430 68.420 ;
        RECT 77.590 66.545 77.880 71.140 ;
        RECT 77.650 66.300 77.820 66.545 ;
        RECT 77.800 64.090 78.930 65.090 ;
        RECT 79.680 64.780 79.970 70.840 ;
        RECT 81.770 66.545 82.060 71.140 ;
        RECT 81.830 66.300 82.000 66.545 ;
        RECT 83.860 64.880 84.150 70.840 ;
        RECT 85.950 66.545 86.240 71.140 ;
        RECT 87.910 68.755 90.255 68.900 ;
        RECT 91.055 68.755 93.400 68.900 ;
        RECT 87.910 68.585 93.400 68.755 ;
        RECT 87.910 68.420 90.255 68.585 ;
        RECT 91.055 68.420 93.400 68.585 ;
        RECT 86.010 66.535 86.205 66.545 ;
        RECT 86.010 66.300 86.180 66.535 ;
        RECT 83.860 64.780 84.680 64.880 ;
        RECT 79.680 64.280 84.680 64.780 ;
        RECT 73.450 62.160 74.630 62.360 ;
        RECT 73.450 61.560 75.130 62.160 ;
        RECT 73.450 61.280 74.630 61.560 ;
        RECT 74.630 55.300 74.920 59.645 ;
        RECT 77.080 58.020 77.250 62.875 ;
        RECT 77.590 58.020 77.880 62.870 ;
        RECT 79.680 58.330 79.970 64.280 ;
        RECT 87.910 63.760 88.080 68.420 ;
        RECT 88.420 63.590 88.710 68.420 ;
        RECT 90.510 63.150 90.800 68.150 ;
        RECT 92.600 63.590 92.890 68.420 ;
        RECT 93.230 63.820 93.400 68.420 ;
        RECT 95.565 66.790 95.855 71.140 ;
        RECT 95.800 64.880 97.000 65.190 ;
        RECT 95.300 64.260 97.000 64.880 ;
        RECT 95.800 64.060 97.000 64.260 ;
        RECT 97.650 63.150 97.945 70.830 ;
        RECT 99.745 66.790 100.035 71.140 ;
        RECT 102.835 68.870 104.930 68.900 ;
        RECT 102.680 68.705 104.930 68.870 ;
        RECT 101.530 68.535 104.930 68.705 ;
        RECT 101.530 65.560 101.700 68.535 ;
        RECT 102.680 68.450 104.930 68.535 ;
        RECT 102.835 68.420 104.930 68.450 ;
        RECT 102.035 64.975 102.330 68.050 ;
        RECT 101.805 64.195 102.545 64.975 ;
        RECT 81.770 58.020 82.060 62.870 ;
        RECT 82.400 58.020 82.570 62.875 ;
        RECT 87.870 62.650 100.465 63.150 ;
        RECT 87.870 61.210 88.370 62.650 ;
        RECT 89.400 61.620 93.400 62.220 ;
        RECT 91.400 61.500 93.400 61.620 ;
        RECT 86.330 60.920 90.800 61.210 ;
        RECT 91.400 60.920 92.600 61.500 ;
        RECT 84.300 59.895 84.470 60.130 ;
        RECT 84.275 59.885 84.470 59.895 ;
        RECT 77.080 57.895 79.425 58.020 ;
        RECT 80.225 57.990 82.570 58.020 ;
        RECT 80.225 57.895 82.750 57.990 ;
        RECT 77.080 57.725 82.750 57.895 ;
        RECT 77.080 57.540 79.425 57.725 ;
        RECT 80.225 57.570 82.750 57.725 ;
        RECT 80.225 57.540 82.570 57.570 ;
        RECT 84.240 55.300 84.530 59.885 ;
        RECT 86.330 55.590 86.620 60.920 ;
        RECT 88.480 59.885 88.650 60.110 ;
        RECT 88.420 55.300 88.710 59.885 ;
        RECT 90.510 55.590 90.800 60.920 ;
        RECT 92.660 59.885 92.830 60.110 ;
        RECT 92.600 55.300 92.890 59.885 ;
        RECT 95.055 58.020 95.225 61.945 ;
        RECT 95.565 58.020 95.855 62.090 ;
        RECT 97.655 58.385 97.950 62.650 ;
        RECT 95.055 57.990 97.150 58.020 ;
        RECT 95.055 57.900 97.305 57.990 ;
        RECT 98.285 57.900 98.455 61.935 ;
        RECT 99.965 61.500 100.465 62.650 ;
        RECT 95.055 57.730 98.455 57.900 ;
        RECT 95.055 57.570 97.305 57.730 ;
        RECT 95.055 57.540 97.150 57.570 ;
        RECT 99.950 55.300 100.240 59.645 ;
        RECT 102.035 55.605 102.330 64.195 ;
        RECT 104.130 64.010 104.420 68.420 ;
        RECT 104.760 64.005 104.930 68.420 ;
        RECT 107.090 66.545 107.380 71.140 ;
        RECT 107.150 66.300 107.320 66.545 ;
        RECT 107.300 64.090 108.430 65.090 ;
        RECT 109.180 64.780 109.470 70.840 ;
        RECT 111.270 66.545 111.560 71.140 ;
        RECT 111.330 66.300 111.500 66.545 ;
        RECT 113.360 64.880 113.650 70.840 ;
        RECT 115.450 66.545 115.740 71.140 ;
        RECT 117.410 68.755 119.755 68.900 ;
        RECT 120.555 68.755 122.900 68.900 ;
        RECT 117.410 68.585 122.900 68.755 ;
        RECT 117.410 68.420 119.755 68.585 ;
        RECT 120.555 68.420 122.900 68.585 ;
        RECT 115.510 66.535 115.705 66.545 ;
        RECT 115.510 66.300 115.680 66.535 ;
        RECT 113.360 64.780 114.180 64.880 ;
        RECT 109.180 64.280 114.180 64.780 ;
        RECT 102.950 62.160 104.130 62.360 ;
        RECT 102.950 61.560 104.630 62.160 ;
        RECT 102.950 61.280 104.130 61.560 ;
        RECT 104.130 55.300 104.420 59.645 ;
        RECT 106.580 58.020 106.750 62.875 ;
        RECT 107.090 58.020 107.380 62.870 ;
        RECT 109.180 58.330 109.470 64.280 ;
        RECT 117.410 63.760 117.580 68.420 ;
        RECT 117.920 63.590 118.210 68.420 ;
        RECT 120.010 63.150 120.300 68.150 ;
        RECT 122.100 63.590 122.390 68.420 ;
        RECT 122.730 63.820 122.900 68.420 ;
        RECT 125.065 66.790 125.355 71.140 ;
        RECT 125.300 64.880 126.500 65.190 ;
        RECT 124.800 64.260 126.500 64.880 ;
        RECT 125.300 64.060 126.500 64.260 ;
        RECT 127.150 63.150 127.445 70.830 ;
        RECT 129.245 66.790 129.535 71.140 ;
        RECT 132.335 68.870 134.430 68.900 ;
        RECT 132.180 68.705 134.430 68.870 ;
        RECT 131.030 68.535 134.430 68.705 ;
        RECT 131.030 65.560 131.200 68.535 ;
        RECT 132.180 68.450 134.430 68.535 ;
        RECT 132.335 68.420 134.430 68.450 ;
        RECT 131.535 64.975 131.830 68.050 ;
        RECT 131.305 64.195 132.045 64.975 ;
        RECT 111.270 58.020 111.560 62.870 ;
        RECT 111.900 58.020 112.070 62.875 ;
        RECT 117.370 62.650 129.965 63.150 ;
        RECT 117.370 61.210 117.870 62.650 ;
        RECT 118.900 61.620 122.900 62.220 ;
        RECT 120.900 61.500 122.900 61.620 ;
        RECT 115.830 60.920 120.300 61.210 ;
        RECT 120.900 60.920 122.100 61.500 ;
        RECT 113.800 59.895 113.970 60.130 ;
        RECT 113.775 59.885 113.970 59.895 ;
        RECT 106.580 57.895 108.925 58.020 ;
        RECT 109.725 57.990 112.070 58.020 ;
        RECT 109.725 57.895 112.250 57.990 ;
        RECT 106.580 57.725 112.250 57.895 ;
        RECT 106.580 57.540 108.925 57.725 ;
        RECT 109.725 57.570 112.250 57.725 ;
        RECT 109.725 57.540 112.070 57.570 ;
        RECT 113.740 55.300 114.030 59.885 ;
        RECT 115.830 55.590 116.120 60.920 ;
        RECT 117.980 59.885 118.150 60.110 ;
        RECT 117.920 55.300 118.210 59.885 ;
        RECT 120.010 55.590 120.300 60.920 ;
        RECT 122.160 59.885 122.330 60.110 ;
        RECT 122.100 55.300 122.390 59.885 ;
        RECT 124.555 58.020 124.725 61.945 ;
        RECT 125.065 58.020 125.355 62.090 ;
        RECT 127.155 58.385 127.450 62.650 ;
        RECT 124.555 57.990 126.650 58.020 ;
        RECT 124.555 57.900 126.805 57.990 ;
        RECT 127.785 57.900 127.955 61.935 ;
        RECT 129.465 61.500 129.965 62.650 ;
        RECT 124.555 57.730 127.955 57.900 ;
        RECT 124.555 57.570 126.805 57.730 ;
        RECT 124.555 57.540 126.650 57.570 ;
        RECT 129.450 55.300 129.740 59.645 ;
        RECT 131.535 55.605 131.830 64.195 ;
        RECT 133.630 64.010 133.920 68.420 ;
        RECT 134.260 64.005 134.430 68.420 ;
        RECT 136.590 66.545 136.880 71.140 ;
        RECT 136.650 66.300 136.820 66.545 ;
        RECT 136.800 64.090 137.930 65.090 ;
        RECT 138.680 64.780 138.970 70.840 ;
        RECT 140.770 66.545 141.060 71.140 ;
        RECT 140.830 66.300 141.000 66.545 ;
        RECT 142.860 64.880 143.150 70.840 ;
        RECT 144.950 66.545 145.240 71.140 ;
        RECT 146.910 68.755 149.255 68.900 ;
        RECT 150.055 68.755 152.400 68.900 ;
        RECT 146.910 68.585 152.400 68.755 ;
        RECT 146.910 68.420 149.255 68.585 ;
        RECT 150.055 68.420 152.400 68.585 ;
        RECT 145.010 66.535 145.205 66.545 ;
        RECT 145.010 66.300 145.180 66.535 ;
        RECT 142.860 64.780 143.680 64.880 ;
        RECT 138.680 64.280 143.680 64.780 ;
        RECT 132.450 62.160 133.630 62.360 ;
        RECT 132.450 61.560 134.130 62.160 ;
        RECT 132.450 61.280 133.630 61.560 ;
        RECT 133.630 55.300 133.920 59.645 ;
        RECT 136.080 58.020 136.250 62.875 ;
        RECT 136.590 58.020 136.880 62.870 ;
        RECT 138.680 58.330 138.970 64.280 ;
        RECT 146.910 63.760 147.080 68.420 ;
        RECT 147.420 63.590 147.710 68.420 ;
        RECT 149.510 63.150 149.800 68.150 ;
        RECT 151.600 63.590 151.890 68.420 ;
        RECT 152.230 63.820 152.400 68.420 ;
        RECT 154.565 66.790 154.855 71.140 ;
        RECT 154.800 64.880 156.000 65.190 ;
        RECT 154.300 64.260 156.000 64.880 ;
        RECT 154.800 64.060 156.000 64.260 ;
        RECT 156.650 63.150 156.945 70.830 ;
        RECT 158.745 66.790 159.035 71.140 ;
        RECT 161.835 68.870 163.930 68.900 ;
        RECT 161.680 68.705 163.930 68.870 ;
        RECT 160.530 68.535 163.930 68.705 ;
        RECT 160.530 65.560 160.700 68.535 ;
        RECT 161.680 68.450 163.930 68.535 ;
        RECT 161.835 68.420 163.930 68.450 ;
        RECT 161.035 64.975 161.330 68.050 ;
        RECT 160.805 64.195 161.545 64.975 ;
        RECT 140.770 58.020 141.060 62.870 ;
        RECT 141.400 58.020 141.570 62.875 ;
        RECT 146.870 62.650 159.465 63.150 ;
        RECT 146.870 61.210 147.370 62.650 ;
        RECT 148.400 61.620 152.400 62.220 ;
        RECT 150.400 61.500 152.400 61.620 ;
        RECT 145.330 60.920 149.800 61.210 ;
        RECT 150.400 60.920 151.600 61.500 ;
        RECT 143.300 59.895 143.470 60.130 ;
        RECT 143.275 59.885 143.470 59.895 ;
        RECT 136.080 57.895 138.425 58.020 ;
        RECT 139.225 57.990 141.570 58.020 ;
        RECT 139.225 57.895 141.750 57.990 ;
        RECT 136.080 57.725 141.750 57.895 ;
        RECT 136.080 57.540 138.425 57.725 ;
        RECT 139.225 57.570 141.750 57.725 ;
        RECT 139.225 57.540 141.570 57.570 ;
        RECT 143.240 55.300 143.530 59.885 ;
        RECT 145.330 55.590 145.620 60.920 ;
        RECT 147.480 59.885 147.650 60.110 ;
        RECT 147.420 55.300 147.710 59.885 ;
        RECT 149.510 55.590 149.800 60.920 ;
        RECT 151.660 59.885 151.830 60.110 ;
        RECT 151.600 55.300 151.890 59.885 ;
        RECT 154.055 58.020 154.225 61.945 ;
        RECT 154.565 58.020 154.855 62.090 ;
        RECT 156.655 58.385 156.950 62.650 ;
        RECT 154.055 57.990 156.150 58.020 ;
        RECT 154.055 57.900 156.305 57.990 ;
        RECT 157.285 57.900 157.455 61.935 ;
        RECT 158.965 61.500 159.465 62.650 ;
        RECT 154.055 57.730 157.455 57.900 ;
        RECT 154.055 57.570 156.305 57.730 ;
        RECT 154.055 57.540 156.150 57.570 ;
        RECT 158.950 55.300 159.240 59.645 ;
        RECT 161.035 55.605 161.330 64.195 ;
        RECT 163.130 64.010 163.420 68.420 ;
        RECT 163.760 64.005 163.930 68.420 ;
        RECT 161.950 62.160 163.130 62.360 ;
        RECT 161.950 61.560 163.630 62.160 ;
        RECT 161.950 61.280 163.130 61.560 ;
        RECT 163.130 55.300 163.420 59.645 ;
        RECT 24.730 54.820 27.080 55.300 ;
        RECT 28.130 54.820 30.990 55.300 ;
        RECT 32.055 54.820 34.400 55.300 ;
        RECT 40.440 55.270 42.780 55.300 ;
        RECT 43.590 55.270 45.930 55.300 ;
        RECT 40.440 54.850 42.785 55.270 ;
        RECT 43.585 54.850 45.930 55.270 ;
        RECT 40.440 54.820 42.780 54.850 ;
        RECT 43.590 54.820 45.930 54.850 ;
        RECT 54.230 54.820 56.580 55.300 ;
        RECT 57.630 54.820 60.490 55.300 ;
        RECT 61.555 54.820 63.900 55.300 ;
        RECT 69.940 55.270 72.280 55.300 ;
        RECT 73.090 55.270 75.430 55.300 ;
        RECT 69.940 54.850 72.285 55.270 ;
        RECT 73.085 54.850 75.430 55.270 ;
        RECT 69.940 54.820 72.280 54.850 ;
        RECT 73.090 54.820 75.430 54.850 ;
        RECT 83.730 54.820 86.080 55.300 ;
        RECT 87.130 54.820 89.990 55.300 ;
        RECT 91.055 54.820 93.400 55.300 ;
        RECT 99.440 55.270 101.780 55.300 ;
        RECT 102.590 55.270 104.930 55.300 ;
        RECT 99.440 54.850 101.785 55.270 ;
        RECT 102.585 54.850 104.930 55.270 ;
        RECT 99.440 54.820 101.780 54.850 ;
        RECT 102.590 54.820 104.930 54.850 ;
        RECT 113.230 54.820 115.580 55.300 ;
        RECT 116.630 54.820 119.490 55.300 ;
        RECT 120.555 54.820 122.900 55.300 ;
        RECT 128.940 55.270 131.280 55.300 ;
        RECT 132.090 55.270 134.430 55.300 ;
        RECT 128.940 54.850 131.285 55.270 ;
        RECT 132.085 54.850 134.430 55.270 ;
        RECT 128.940 54.820 131.280 54.850 ;
        RECT 132.090 54.820 134.430 54.850 ;
        RECT 142.730 54.820 145.080 55.300 ;
        RECT 146.130 54.820 148.990 55.300 ;
        RECT 150.055 54.820 152.400 55.300 ;
        RECT 158.440 55.270 160.780 55.300 ;
        RECT 161.590 55.270 163.930 55.300 ;
        RECT 158.440 54.850 160.785 55.270 ;
        RECT 161.585 54.850 163.930 55.270 ;
        RECT 158.440 54.820 160.780 54.850 ;
        RECT 161.590 54.820 163.930 54.850 ;
        RECT 165.510 53.500 166.010 73.000 ;
        RECT 171.930 59.500 173.930 59.670 ;
        RECT 172.010 59.470 173.850 59.500 ;
        RECT 175.060 59.040 177.060 59.210 ;
        RECT 175.140 59.010 176.980 59.040 ;
        RECT 172.010 55.120 173.850 55.150 ;
        RECT 171.930 54.950 173.930 55.120 ;
        RECT 175.140 54.660 176.980 54.690 ;
        RECT 175.060 54.490 177.060 54.660 ;
        RECT 15.430 53.000 166.090 53.500 ;
        RECT 0.430 51.000 180.090 51.500 ;
        RECT 0.510 31.500 1.010 51.000 ;
        RECT 2.480 49.830 4.820 49.860 ;
        RECT 5.630 49.830 7.970 49.860 ;
        RECT 2.480 49.410 4.825 49.830 ;
        RECT 5.625 49.410 7.970 49.830 ;
        RECT 2.480 49.380 4.820 49.410 ;
        RECT 5.630 49.380 7.970 49.410 ;
        RECT 14.010 49.380 16.355 49.860 ;
        RECT 17.420 49.380 20.280 49.860 ;
        RECT 21.330 49.380 23.680 49.860 ;
        RECT 31.980 49.830 34.320 49.860 ;
        RECT 35.130 49.830 37.470 49.860 ;
        RECT 31.980 49.410 34.325 49.830 ;
        RECT 35.125 49.410 37.470 49.830 ;
        RECT 31.980 49.380 34.320 49.410 ;
        RECT 35.130 49.380 37.470 49.410 ;
        RECT 43.510 49.380 45.855 49.860 ;
        RECT 46.920 49.380 49.780 49.860 ;
        RECT 50.830 49.380 53.180 49.860 ;
        RECT 61.480 49.830 63.820 49.860 ;
        RECT 64.630 49.830 66.970 49.860 ;
        RECT 61.480 49.410 63.825 49.830 ;
        RECT 64.625 49.410 66.970 49.830 ;
        RECT 61.480 49.380 63.820 49.410 ;
        RECT 64.630 49.380 66.970 49.410 ;
        RECT 73.010 49.380 75.355 49.860 ;
        RECT 76.420 49.380 79.280 49.860 ;
        RECT 80.330 49.380 82.680 49.860 ;
        RECT 90.980 49.830 93.320 49.860 ;
        RECT 94.130 49.830 96.470 49.860 ;
        RECT 90.980 49.410 93.325 49.830 ;
        RECT 94.125 49.410 96.470 49.830 ;
        RECT 90.980 49.380 93.320 49.410 ;
        RECT 94.130 49.380 96.470 49.410 ;
        RECT 102.510 49.380 104.855 49.860 ;
        RECT 105.920 49.380 108.780 49.860 ;
        RECT 109.830 49.380 112.180 49.860 ;
        RECT 120.480 49.830 122.820 49.860 ;
        RECT 123.630 49.830 125.970 49.860 ;
        RECT 120.480 49.410 122.825 49.830 ;
        RECT 123.625 49.410 125.970 49.830 ;
        RECT 120.480 49.380 122.820 49.410 ;
        RECT 123.630 49.380 125.970 49.410 ;
        RECT 132.010 49.380 134.355 49.860 ;
        RECT 135.420 49.380 138.280 49.860 ;
        RECT 139.330 49.380 141.680 49.860 ;
        RECT 149.980 49.830 152.320 49.860 ;
        RECT 153.130 49.830 155.470 49.860 ;
        RECT 149.980 49.410 152.325 49.830 ;
        RECT 153.125 49.410 155.470 49.830 ;
        RECT 149.980 49.380 152.320 49.410 ;
        RECT 153.130 49.380 155.470 49.410 ;
        RECT 161.510 49.380 163.855 49.860 ;
        RECT 164.920 49.380 167.780 49.860 ;
        RECT 168.830 49.380 171.180 49.860 ;
        RECT 2.990 45.035 3.280 49.380 ;
        RECT 3.280 43.120 4.460 43.400 ;
        RECT 2.780 42.520 4.460 43.120 ;
        RECT 3.280 42.320 4.460 42.520 ;
        RECT 2.480 36.260 2.650 40.675 ;
        RECT 2.990 36.260 3.280 40.670 ;
        RECT 5.080 40.485 5.375 49.075 ;
        RECT 7.170 45.035 7.460 49.380 ;
        RECT 10.260 47.110 12.355 47.140 ;
        RECT 10.105 46.950 12.355 47.110 ;
        RECT 8.955 46.780 12.355 46.950 ;
        RECT 6.945 42.030 7.445 43.180 ;
        RECT 8.955 42.745 9.125 46.780 ;
        RECT 10.105 46.690 12.355 46.780 ;
        RECT 10.260 46.660 12.355 46.690 ;
        RECT 9.460 42.030 9.755 46.295 ;
        RECT 11.555 42.590 11.845 46.660 ;
        RECT 12.185 42.735 12.355 46.660 ;
        RECT 14.520 44.795 14.810 49.380 ;
        RECT 14.580 44.570 14.750 44.795 ;
        RECT 16.610 43.760 16.900 49.090 ;
        RECT 18.700 44.795 18.990 49.380 ;
        RECT 18.760 44.570 18.930 44.795 ;
        RECT 20.790 43.760 21.080 49.090 ;
        RECT 22.880 44.795 23.170 49.380 ;
        RECT 24.840 47.110 27.185 47.140 ;
        RECT 24.660 46.955 27.185 47.110 ;
        RECT 27.985 46.955 30.330 47.140 ;
        RECT 24.660 46.785 30.330 46.955 ;
        RECT 24.660 46.690 27.185 46.785 ;
        RECT 24.840 46.660 27.185 46.690 ;
        RECT 27.985 46.660 30.330 46.785 ;
        RECT 22.940 44.785 23.135 44.795 ;
        RECT 22.940 44.550 23.110 44.785 ;
        RECT 14.810 43.180 16.010 43.760 ;
        RECT 16.610 43.470 21.080 43.760 ;
        RECT 14.010 43.060 16.010 43.180 ;
        RECT 14.010 42.460 18.010 43.060 ;
        RECT 19.040 42.030 19.540 43.470 ;
        RECT 6.945 41.530 19.540 42.030 ;
        RECT 24.840 41.805 25.010 46.660 ;
        RECT 25.350 41.810 25.640 46.660 ;
        RECT 4.865 39.705 5.605 40.485 ;
        RECT 5.080 36.630 5.375 39.705 ;
        RECT 2.480 36.230 4.575 36.260 ;
        RECT 2.480 36.145 4.730 36.230 ;
        RECT 5.710 36.145 5.880 39.120 ;
        RECT 2.480 35.975 5.880 36.145 ;
        RECT 2.480 35.810 4.730 35.975 ;
        RECT 2.480 35.780 4.575 35.810 ;
        RECT 7.375 33.540 7.665 37.890 ;
        RECT 9.465 33.850 9.760 41.530 ;
        RECT 10.410 40.420 11.610 40.620 ;
        RECT 10.410 39.800 12.110 40.420 ;
        RECT 10.410 39.490 11.610 39.800 ;
        RECT 11.555 33.540 11.845 37.890 ;
        RECT 14.010 36.260 14.180 40.860 ;
        RECT 14.520 36.260 14.810 41.090 ;
        RECT 16.610 36.530 16.900 41.530 ;
        RECT 18.700 36.260 18.990 41.090 ;
        RECT 19.330 36.260 19.500 40.920 ;
        RECT 27.440 40.400 27.730 46.350 ;
        RECT 29.530 41.810 29.820 46.660 ;
        RECT 30.160 41.805 30.330 46.660 ;
        RECT 32.490 45.035 32.780 49.380 ;
        RECT 32.780 43.120 33.960 43.400 ;
        RECT 32.280 42.520 33.960 43.120 ;
        RECT 32.780 42.320 33.960 42.520 ;
        RECT 22.730 39.900 27.730 40.400 ;
        RECT 22.730 39.800 23.550 39.900 ;
        RECT 21.230 38.145 21.400 38.380 ;
        RECT 21.205 38.135 21.400 38.145 ;
        RECT 14.010 36.095 16.355 36.260 ;
        RECT 17.155 36.095 19.500 36.260 ;
        RECT 14.010 35.925 19.500 36.095 ;
        RECT 14.010 35.780 16.355 35.925 ;
        RECT 17.155 35.780 19.500 35.925 ;
        RECT 21.170 33.540 21.460 38.135 ;
        RECT 23.260 33.840 23.550 39.800 ;
        RECT 25.410 38.135 25.580 38.380 ;
        RECT 25.350 33.540 25.640 38.135 ;
        RECT 27.440 33.840 27.730 39.900 ;
        RECT 28.480 39.590 29.610 40.590 ;
        RECT 29.590 38.135 29.760 38.380 ;
        RECT 29.530 33.540 29.820 38.135 ;
        RECT 31.980 36.260 32.150 40.675 ;
        RECT 32.490 36.260 32.780 40.670 ;
        RECT 34.580 40.485 34.875 49.075 ;
        RECT 36.670 45.035 36.960 49.380 ;
        RECT 39.760 47.110 41.855 47.140 ;
        RECT 39.605 46.950 41.855 47.110 ;
        RECT 38.455 46.780 41.855 46.950 ;
        RECT 36.445 42.030 36.945 43.180 ;
        RECT 38.455 42.745 38.625 46.780 ;
        RECT 39.605 46.690 41.855 46.780 ;
        RECT 39.760 46.660 41.855 46.690 ;
        RECT 38.960 42.030 39.255 46.295 ;
        RECT 41.055 42.590 41.345 46.660 ;
        RECT 41.685 42.735 41.855 46.660 ;
        RECT 44.020 44.795 44.310 49.380 ;
        RECT 44.080 44.570 44.250 44.795 ;
        RECT 46.110 43.760 46.400 49.090 ;
        RECT 48.200 44.795 48.490 49.380 ;
        RECT 48.260 44.570 48.430 44.795 ;
        RECT 50.290 43.760 50.580 49.090 ;
        RECT 52.380 44.795 52.670 49.380 ;
        RECT 54.340 47.110 56.685 47.140 ;
        RECT 54.160 46.955 56.685 47.110 ;
        RECT 57.485 46.955 59.830 47.140 ;
        RECT 54.160 46.785 59.830 46.955 ;
        RECT 54.160 46.690 56.685 46.785 ;
        RECT 54.340 46.660 56.685 46.690 ;
        RECT 57.485 46.660 59.830 46.785 ;
        RECT 52.440 44.785 52.635 44.795 ;
        RECT 52.440 44.550 52.610 44.785 ;
        RECT 44.310 43.180 45.510 43.760 ;
        RECT 46.110 43.470 50.580 43.760 ;
        RECT 43.510 43.060 45.510 43.180 ;
        RECT 43.510 42.460 47.510 43.060 ;
        RECT 48.540 42.030 49.040 43.470 ;
        RECT 36.445 41.530 49.040 42.030 ;
        RECT 54.340 41.805 54.510 46.660 ;
        RECT 54.850 41.810 55.140 46.660 ;
        RECT 34.365 39.705 35.105 40.485 ;
        RECT 34.580 36.630 34.875 39.705 ;
        RECT 31.980 36.230 34.075 36.260 ;
        RECT 31.980 36.145 34.230 36.230 ;
        RECT 35.210 36.145 35.380 39.120 ;
        RECT 31.980 35.975 35.380 36.145 ;
        RECT 31.980 35.810 34.230 35.975 ;
        RECT 31.980 35.780 34.075 35.810 ;
        RECT 36.875 33.540 37.165 37.890 ;
        RECT 38.965 33.850 39.260 41.530 ;
        RECT 39.910 40.420 41.110 40.620 ;
        RECT 39.910 39.800 41.610 40.420 ;
        RECT 39.910 39.490 41.110 39.800 ;
        RECT 41.055 33.540 41.345 37.890 ;
        RECT 43.510 36.260 43.680 40.860 ;
        RECT 44.020 36.260 44.310 41.090 ;
        RECT 46.110 36.530 46.400 41.530 ;
        RECT 48.200 36.260 48.490 41.090 ;
        RECT 48.830 36.260 49.000 40.920 ;
        RECT 56.940 40.400 57.230 46.350 ;
        RECT 59.030 41.810 59.320 46.660 ;
        RECT 59.660 41.805 59.830 46.660 ;
        RECT 61.990 45.035 62.280 49.380 ;
        RECT 62.280 43.120 63.460 43.400 ;
        RECT 61.780 42.520 63.460 43.120 ;
        RECT 62.280 42.320 63.460 42.520 ;
        RECT 52.230 39.900 57.230 40.400 ;
        RECT 52.230 39.800 53.050 39.900 ;
        RECT 50.730 38.145 50.900 38.380 ;
        RECT 50.705 38.135 50.900 38.145 ;
        RECT 43.510 36.095 45.855 36.260 ;
        RECT 46.655 36.095 49.000 36.260 ;
        RECT 43.510 35.925 49.000 36.095 ;
        RECT 43.510 35.780 45.855 35.925 ;
        RECT 46.655 35.780 49.000 35.925 ;
        RECT 50.670 33.540 50.960 38.135 ;
        RECT 52.760 33.840 53.050 39.800 ;
        RECT 54.910 38.135 55.080 38.380 ;
        RECT 54.850 33.540 55.140 38.135 ;
        RECT 56.940 33.840 57.230 39.900 ;
        RECT 57.980 39.590 59.110 40.590 ;
        RECT 59.090 38.135 59.260 38.380 ;
        RECT 59.030 33.540 59.320 38.135 ;
        RECT 61.480 36.260 61.650 40.675 ;
        RECT 61.990 36.260 62.280 40.670 ;
        RECT 64.080 40.485 64.375 49.075 ;
        RECT 66.170 45.035 66.460 49.380 ;
        RECT 69.260 47.110 71.355 47.140 ;
        RECT 69.105 46.950 71.355 47.110 ;
        RECT 67.955 46.780 71.355 46.950 ;
        RECT 65.945 42.030 66.445 43.180 ;
        RECT 67.955 42.745 68.125 46.780 ;
        RECT 69.105 46.690 71.355 46.780 ;
        RECT 69.260 46.660 71.355 46.690 ;
        RECT 68.460 42.030 68.755 46.295 ;
        RECT 70.555 42.590 70.845 46.660 ;
        RECT 71.185 42.735 71.355 46.660 ;
        RECT 73.520 44.795 73.810 49.380 ;
        RECT 73.580 44.570 73.750 44.795 ;
        RECT 75.610 43.760 75.900 49.090 ;
        RECT 77.700 44.795 77.990 49.380 ;
        RECT 77.760 44.570 77.930 44.795 ;
        RECT 79.790 43.760 80.080 49.090 ;
        RECT 81.880 44.795 82.170 49.380 ;
        RECT 83.840 47.110 86.185 47.140 ;
        RECT 83.660 46.955 86.185 47.110 ;
        RECT 86.985 46.955 89.330 47.140 ;
        RECT 83.660 46.785 89.330 46.955 ;
        RECT 83.660 46.690 86.185 46.785 ;
        RECT 83.840 46.660 86.185 46.690 ;
        RECT 86.985 46.660 89.330 46.785 ;
        RECT 81.940 44.785 82.135 44.795 ;
        RECT 81.940 44.550 82.110 44.785 ;
        RECT 73.810 43.180 75.010 43.760 ;
        RECT 75.610 43.470 80.080 43.760 ;
        RECT 73.010 43.060 75.010 43.180 ;
        RECT 73.010 42.460 77.010 43.060 ;
        RECT 78.040 42.030 78.540 43.470 ;
        RECT 65.945 41.530 78.540 42.030 ;
        RECT 83.840 41.805 84.010 46.660 ;
        RECT 84.350 41.810 84.640 46.660 ;
        RECT 63.865 39.705 64.605 40.485 ;
        RECT 64.080 36.630 64.375 39.705 ;
        RECT 61.480 36.230 63.575 36.260 ;
        RECT 61.480 36.145 63.730 36.230 ;
        RECT 64.710 36.145 64.880 39.120 ;
        RECT 61.480 35.975 64.880 36.145 ;
        RECT 61.480 35.810 63.730 35.975 ;
        RECT 61.480 35.780 63.575 35.810 ;
        RECT 66.375 33.540 66.665 37.890 ;
        RECT 68.465 33.850 68.760 41.530 ;
        RECT 69.410 40.420 70.610 40.620 ;
        RECT 69.410 39.800 71.110 40.420 ;
        RECT 69.410 39.490 70.610 39.800 ;
        RECT 70.555 33.540 70.845 37.890 ;
        RECT 73.010 36.260 73.180 40.860 ;
        RECT 73.520 36.260 73.810 41.090 ;
        RECT 75.610 36.530 75.900 41.530 ;
        RECT 77.700 36.260 77.990 41.090 ;
        RECT 78.330 36.260 78.500 40.920 ;
        RECT 86.440 40.400 86.730 46.350 ;
        RECT 88.530 41.810 88.820 46.660 ;
        RECT 89.160 41.805 89.330 46.660 ;
        RECT 91.490 45.035 91.780 49.380 ;
        RECT 91.780 43.120 92.960 43.400 ;
        RECT 91.280 42.520 92.960 43.120 ;
        RECT 91.780 42.320 92.960 42.520 ;
        RECT 81.730 39.900 86.730 40.400 ;
        RECT 81.730 39.800 82.550 39.900 ;
        RECT 80.230 38.145 80.400 38.380 ;
        RECT 80.205 38.135 80.400 38.145 ;
        RECT 73.010 36.095 75.355 36.260 ;
        RECT 76.155 36.095 78.500 36.260 ;
        RECT 73.010 35.925 78.500 36.095 ;
        RECT 73.010 35.780 75.355 35.925 ;
        RECT 76.155 35.780 78.500 35.925 ;
        RECT 80.170 33.540 80.460 38.135 ;
        RECT 82.260 33.840 82.550 39.800 ;
        RECT 84.410 38.135 84.580 38.380 ;
        RECT 84.350 33.540 84.640 38.135 ;
        RECT 86.440 33.840 86.730 39.900 ;
        RECT 87.480 39.590 88.610 40.590 ;
        RECT 88.590 38.135 88.760 38.380 ;
        RECT 88.530 33.540 88.820 38.135 ;
        RECT 90.980 36.260 91.150 40.675 ;
        RECT 91.490 36.260 91.780 40.670 ;
        RECT 93.580 40.485 93.875 49.075 ;
        RECT 95.670 45.035 95.960 49.380 ;
        RECT 98.760 47.110 100.855 47.140 ;
        RECT 98.605 46.950 100.855 47.110 ;
        RECT 97.455 46.780 100.855 46.950 ;
        RECT 95.445 42.030 95.945 43.180 ;
        RECT 97.455 42.745 97.625 46.780 ;
        RECT 98.605 46.690 100.855 46.780 ;
        RECT 98.760 46.660 100.855 46.690 ;
        RECT 97.960 42.030 98.255 46.295 ;
        RECT 100.055 42.590 100.345 46.660 ;
        RECT 100.685 42.735 100.855 46.660 ;
        RECT 103.020 44.795 103.310 49.380 ;
        RECT 103.080 44.570 103.250 44.795 ;
        RECT 105.110 43.760 105.400 49.090 ;
        RECT 107.200 44.795 107.490 49.380 ;
        RECT 107.260 44.570 107.430 44.795 ;
        RECT 109.290 43.760 109.580 49.090 ;
        RECT 111.380 44.795 111.670 49.380 ;
        RECT 113.340 47.110 115.685 47.140 ;
        RECT 113.160 46.955 115.685 47.110 ;
        RECT 116.485 46.955 118.830 47.140 ;
        RECT 113.160 46.785 118.830 46.955 ;
        RECT 113.160 46.690 115.685 46.785 ;
        RECT 113.340 46.660 115.685 46.690 ;
        RECT 116.485 46.660 118.830 46.785 ;
        RECT 111.440 44.785 111.635 44.795 ;
        RECT 111.440 44.550 111.610 44.785 ;
        RECT 103.310 43.180 104.510 43.760 ;
        RECT 105.110 43.470 109.580 43.760 ;
        RECT 102.510 43.060 104.510 43.180 ;
        RECT 102.510 42.460 106.510 43.060 ;
        RECT 107.540 42.030 108.040 43.470 ;
        RECT 95.445 41.530 108.040 42.030 ;
        RECT 113.340 41.805 113.510 46.660 ;
        RECT 113.850 41.810 114.140 46.660 ;
        RECT 93.365 39.705 94.105 40.485 ;
        RECT 93.580 36.630 93.875 39.705 ;
        RECT 90.980 36.230 93.075 36.260 ;
        RECT 90.980 36.145 93.230 36.230 ;
        RECT 94.210 36.145 94.380 39.120 ;
        RECT 90.980 35.975 94.380 36.145 ;
        RECT 90.980 35.810 93.230 35.975 ;
        RECT 90.980 35.780 93.075 35.810 ;
        RECT 95.875 33.540 96.165 37.890 ;
        RECT 97.965 33.850 98.260 41.530 ;
        RECT 98.910 40.420 100.110 40.620 ;
        RECT 98.910 39.800 100.610 40.420 ;
        RECT 98.910 39.490 100.110 39.800 ;
        RECT 100.055 33.540 100.345 37.890 ;
        RECT 102.510 36.260 102.680 40.860 ;
        RECT 103.020 36.260 103.310 41.090 ;
        RECT 105.110 36.530 105.400 41.530 ;
        RECT 107.200 36.260 107.490 41.090 ;
        RECT 107.830 36.260 108.000 40.920 ;
        RECT 115.940 40.400 116.230 46.350 ;
        RECT 118.030 41.810 118.320 46.660 ;
        RECT 118.660 41.805 118.830 46.660 ;
        RECT 120.990 45.035 121.280 49.380 ;
        RECT 121.280 43.120 122.460 43.400 ;
        RECT 120.780 42.520 122.460 43.120 ;
        RECT 121.280 42.320 122.460 42.520 ;
        RECT 111.230 39.900 116.230 40.400 ;
        RECT 111.230 39.800 112.050 39.900 ;
        RECT 109.730 38.145 109.900 38.380 ;
        RECT 109.705 38.135 109.900 38.145 ;
        RECT 102.510 36.095 104.855 36.260 ;
        RECT 105.655 36.095 108.000 36.260 ;
        RECT 102.510 35.925 108.000 36.095 ;
        RECT 102.510 35.780 104.855 35.925 ;
        RECT 105.655 35.780 108.000 35.925 ;
        RECT 109.670 33.540 109.960 38.135 ;
        RECT 111.760 33.840 112.050 39.800 ;
        RECT 113.910 38.135 114.080 38.380 ;
        RECT 113.850 33.540 114.140 38.135 ;
        RECT 115.940 33.840 116.230 39.900 ;
        RECT 116.980 39.590 118.110 40.590 ;
        RECT 118.090 38.135 118.260 38.380 ;
        RECT 118.030 33.540 118.320 38.135 ;
        RECT 120.480 36.260 120.650 40.675 ;
        RECT 120.990 36.260 121.280 40.670 ;
        RECT 123.080 40.485 123.375 49.075 ;
        RECT 125.170 45.035 125.460 49.380 ;
        RECT 128.260 47.110 130.355 47.140 ;
        RECT 128.105 46.950 130.355 47.110 ;
        RECT 126.955 46.780 130.355 46.950 ;
        RECT 124.945 42.030 125.445 43.180 ;
        RECT 126.955 42.745 127.125 46.780 ;
        RECT 128.105 46.690 130.355 46.780 ;
        RECT 128.260 46.660 130.355 46.690 ;
        RECT 127.460 42.030 127.755 46.295 ;
        RECT 129.555 42.590 129.845 46.660 ;
        RECT 130.185 42.735 130.355 46.660 ;
        RECT 132.520 44.795 132.810 49.380 ;
        RECT 132.580 44.570 132.750 44.795 ;
        RECT 134.610 43.760 134.900 49.090 ;
        RECT 136.700 44.795 136.990 49.380 ;
        RECT 136.760 44.570 136.930 44.795 ;
        RECT 138.790 43.760 139.080 49.090 ;
        RECT 140.880 44.795 141.170 49.380 ;
        RECT 142.840 47.110 145.185 47.140 ;
        RECT 142.660 46.955 145.185 47.110 ;
        RECT 145.985 46.955 148.330 47.140 ;
        RECT 142.660 46.785 148.330 46.955 ;
        RECT 142.660 46.690 145.185 46.785 ;
        RECT 142.840 46.660 145.185 46.690 ;
        RECT 145.985 46.660 148.330 46.785 ;
        RECT 140.940 44.785 141.135 44.795 ;
        RECT 140.940 44.550 141.110 44.785 ;
        RECT 132.810 43.180 134.010 43.760 ;
        RECT 134.610 43.470 139.080 43.760 ;
        RECT 132.010 43.060 134.010 43.180 ;
        RECT 132.010 42.460 136.010 43.060 ;
        RECT 137.040 42.030 137.540 43.470 ;
        RECT 124.945 41.530 137.540 42.030 ;
        RECT 142.840 41.805 143.010 46.660 ;
        RECT 143.350 41.810 143.640 46.660 ;
        RECT 122.865 39.705 123.605 40.485 ;
        RECT 123.080 36.630 123.375 39.705 ;
        RECT 120.480 36.230 122.575 36.260 ;
        RECT 120.480 36.145 122.730 36.230 ;
        RECT 123.710 36.145 123.880 39.120 ;
        RECT 120.480 35.975 123.880 36.145 ;
        RECT 120.480 35.810 122.730 35.975 ;
        RECT 120.480 35.780 122.575 35.810 ;
        RECT 125.375 33.540 125.665 37.890 ;
        RECT 127.465 33.850 127.760 41.530 ;
        RECT 128.410 40.420 129.610 40.620 ;
        RECT 128.410 39.800 130.110 40.420 ;
        RECT 128.410 39.490 129.610 39.800 ;
        RECT 129.555 33.540 129.845 37.890 ;
        RECT 132.010 36.260 132.180 40.860 ;
        RECT 132.520 36.260 132.810 41.090 ;
        RECT 134.610 36.530 134.900 41.530 ;
        RECT 136.700 36.260 136.990 41.090 ;
        RECT 137.330 36.260 137.500 40.920 ;
        RECT 145.440 40.400 145.730 46.350 ;
        RECT 147.530 41.810 147.820 46.660 ;
        RECT 148.160 41.805 148.330 46.660 ;
        RECT 150.490 45.035 150.780 49.380 ;
        RECT 150.780 43.120 151.960 43.400 ;
        RECT 150.280 42.520 151.960 43.120 ;
        RECT 150.780 42.320 151.960 42.520 ;
        RECT 140.730 39.900 145.730 40.400 ;
        RECT 140.730 39.800 141.550 39.900 ;
        RECT 139.230 38.145 139.400 38.380 ;
        RECT 139.205 38.135 139.400 38.145 ;
        RECT 132.010 36.095 134.355 36.260 ;
        RECT 135.155 36.095 137.500 36.260 ;
        RECT 132.010 35.925 137.500 36.095 ;
        RECT 132.010 35.780 134.355 35.925 ;
        RECT 135.155 35.780 137.500 35.925 ;
        RECT 139.170 33.540 139.460 38.135 ;
        RECT 141.260 33.840 141.550 39.800 ;
        RECT 143.410 38.135 143.580 38.380 ;
        RECT 143.350 33.540 143.640 38.135 ;
        RECT 145.440 33.840 145.730 39.900 ;
        RECT 146.480 39.590 147.610 40.590 ;
        RECT 147.590 38.135 147.760 38.380 ;
        RECT 147.530 33.540 147.820 38.135 ;
        RECT 149.980 36.260 150.150 40.675 ;
        RECT 150.490 36.260 150.780 40.670 ;
        RECT 152.580 40.485 152.875 49.075 ;
        RECT 154.670 45.035 154.960 49.380 ;
        RECT 157.760 47.110 159.855 47.140 ;
        RECT 157.605 46.950 159.855 47.110 ;
        RECT 156.455 46.780 159.855 46.950 ;
        RECT 154.445 42.030 154.945 43.180 ;
        RECT 156.455 42.745 156.625 46.780 ;
        RECT 157.605 46.690 159.855 46.780 ;
        RECT 157.760 46.660 159.855 46.690 ;
        RECT 156.960 42.030 157.255 46.295 ;
        RECT 159.055 42.590 159.345 46.660 ;
        RECT 159.685 42.735 159.855 46.660 ;
        RECT 162.020 44.795 162.310 49.380 ;
        RECT 162.080 44.570 162.250 44.795 ;
        RECT 164.110 43.760 164.400 49.090 ;
        RECT 166.200 44.795 166.490 49.380 ;
        RECT 166.260 44.570 166.430 44.795 ;
        RECT 168.290 43.760 168.580 49.090 ;
        RECT 170.380 44.795 170.670 49.380 ;
        RECT 172.340 47.110 174.685 47.140 ;
        RECT 172.160 46.955 174.685 47.110 ;
        RECT 175.485 46.955 177.830 47.140 ;
        RECT 172.160 46.785 177.830 46.955 ;
        RECT 172.160 46.690 174.685 46.785 ;
        RECT 172.340 46.660 174.685 46.690 ;
        RECT 175.485 46.660 177.830 46.785 ;
        RECT 170.440 44.785 170.635 44.795 ;
        RECT 170.440 44.550 170.610 44.785 ;
        RECT 162.310 43.180 163.510 43.760 ;
        RECT 164.110 43.470 168.580 43.760 ;
        RECT 161.510 43.060 163.510 43.180 ;
        RECT 161.510 42.460 165.510 43.060 ;
        RECT 166.540 42.030 167.040 43.470 ;
        RECT 154.445 41.530 167.040 42.030 ;
        RECT 172.340 41.805 172.510 46.660 ;
        RECT 172.850 41.810 173.140 46.660 ;
        RECT 152.365 39.705 153.105 40.485 ;
        RECT 152.580 36.630 152.875 39.705 ;
        RECT 149.980 36.230 152.075 36.260 ;
        RECT 149.980 36.145 152.230 36.230 ;
        RECT 153.210 36.145 153.380 39.120 ;
        RECT 149.980 35.975 153.380 36.145 ;
        RECT 149.980 35.810 152.230 35.975 ;
        RECT 149.980 35.780 152.075 35.810 ;
        RECT 154.875 33.540 155.165 37.890 ;
        RECT 156.965 33.850 157.260 41.530 ;
        RECT 157.910 40.420 159.110 40.620 ;
        RECT 157.910 39.800 159.610 40.420 ;
        RECT 157.910 39.490 159.110 39.800 ;
        RECT 159.055 33.540 159.345 37.890 ;
        RECT 161.510 36.260 161.680 40.860 ;
        RECT 162.020 36.260 162.310 41.090 ;
        RECT 164.110 36.530 164.400 41.530 ;
        RECT 166.200 36.260 166.490 41.090 ;
        RECT 166.830 36.260 167.000 40.920 ;
        RECT 174.940 40.400 175.230 46.350 ;
        RECT 177.030 41.810 177.320 46.660 ;
        RECT 177.660 41.805 177.830 46.660 ;
        RECT 170.230 39.900 175.230 40.400 ;
        RECT 170.230 39.800 171.050 39.900 ;
        RECT 168.730 38.145 168.900 38.380 ;
        RECT 168.705 38.135 168.900 38.145 ;
        RECT 161.510 36.095 163.855 36.260 ;
        RECT 164.655 36.095 167.000 36.260 ;
        RECT 161.510 35.925 167.000 36.095 ;
        RECT 161.510 35.780 163.855 35.925 ;
        RECT 164.655 35.780 167.000 35.925 ;
        RECT 168.670 33.540 168.960 38.135 ;
        RECT 170.760 33.840 171.050 39.800 ;
        RECT 172.910 38.135 173.080 38.380 ;
        RECT 172.850 33.540 173.140 38.135 ;
        RECT 174.940 33.840 175.230 39.900 ;
        RECT 175.980 39.590 177.110 40.590 ;
        RECT 177.090 38.135 177.260 38.380 ;
        RECT 177.030 33.540 177.320 38.135 ;
        RECT 6.865 33.060 9.210 33.540 ;
        RECT 10.010 33.060 12.355 33.540 ;
        RECT 20.660 33.060 23.005 33.540 ;
        RECT 24.060 33.060 26.920 33.540 ;
        RECT 27.985 33.060 30.330 33.540 ;
        RECT 36.365 33.060 38.710 33.540 ;
        RECT 39.510 33.060 41.855 33.540 ;
        RECT 50.160 33.060 52.505 33.540 ;
        RECT 53.560 33.060 56.420 33.540 ;
        RECT 57.485 33.060 59.830 33.540 ;
        RECT 65.865 33.060 68.210 33.540 ;
        RECT 69.010 33.060 71.355 33.540 ;
        RECT 79.660 33.060 82.005 33.540 ;
        RECT 83.060 33.060 85.920 33.540 ;
        RECT 86.985 33.060 89.330 33.540 ;
        RECT 95.365 33.060 97.710 33.540 ;
        RECT 98.510 33.060 100.855 33.540 ;
        RECT 109.160 33.060 111.505 33.540 ;
        RECT 112.560 33.060 115.420 33.540 ;
        RECT 116.485 33.060 118.830 33.540 ;
        RECT 124.865 33.060 127.210 33.540 ;
        RECT 128.010 33.060 130.355 33.540 ;
        RECT 138.660 33.060 141.005 33.540 ;
        RECT 142.060 33.060 144.920 33.540 ;
        RECT 145.985 33.060 148.330 33.540 ;
        RECT 154.365 33.060 156.710 33.540 ;
        RECT 157.510 33.060 159.855 33.540 ;
        RECT 168.160 33.060 170.505 33.540 ;
        RECT 171.560 33.060 174.420 33.540 ;
        RECT 175.485 33.060 177.830 33.540 ;
        RECT 179.510 31.500 180.010 51.000 ;
        RECT 0.430 31.000 180.090 31.500 ;
      LAYER mcon ;
        RECT 36.100 73.100 36.400 73.400 ;
        RECT 36.600 73.100 36.900 73.400 ;
        RECT 37.100 73.100 37.400 73.400 ;
        RECT 37.600 73.100 37.900 73.400 ;
        RECT 72.100 73.100 72.400 73.400 ;
        RECT 72.600 73.100 72.900 73.400 ;
        RECT 73.100 73.100 73.400 73.400 ;
        RECT 73.600 73.100 73.900 73.400 ;
        RECT 108.100 73.100 108.400 73.400 ;
        RECT 108.600 73.100 108.900 73.400 ;
        RECT 109.100 73.100 109.400 73.400 ;
        RECT 109.600 73.100 109.900 73.400 ;
        RECT 144.100 73.100 144.400 73.400 ;
        RECT 144.600 73.100 144.900 73.400 ;
        RECT 145.100 73.100 145.400 73.400 ;
        RECT 145.600 73.100 145.900 73.400 ;
        RECT 3.475 63.135 3.645 63.305 ;
        RECT 3.935 63.135 4.105 63.305 ;
        RECT 4.395 63.135 4.565 63.305 ;
        RECT 4.855 63.135 5.025 63.305 ;
        RECT 5.315 63.135 5.485 63.305 ;
        RECT 7.645 63.135 7.815 63.305 ;
        RECT 8.105 63.135 8.275 63.305 ;
        RECT 8.565 63.135 8.735 63.305 ;
        RECT 2.430 61.850 2.630 62.050 ;
        RECT 6.435 61.775 6.605 61.945 ;
        RECT 3.475 60.415 3.645 60.585 ;
        RECT 3.935 60.415 4.105 60.585 ;
        RECT 4.395 60.415 4.565 60.585 ;
        RECT 4.855 60.415 5.025 60.585 ;
        RECT 5.315 60.415 5.485 60.585 ;
        RECT 7.645 60.415 7.815 60.585 ;
        RECT 8.105 60.415 8.275 60.585 ;
        RECT 8.565 60.415 8.735 60.585 ;
        RECT 18.080 71.170 18.595 71.590 ;
        RECT 18.785 71.170 19.205 71.590 ;
        RECT 19.395 71.170 19.815 71.590 ;
        RECT 20.005 71.170 20.425 71.590 ;
        RECT 21.490 71.170 21.910 71.590 ;
        RECT 22.100 71.170 22.520 71.590 ;
        RECT 22.710 71.170 23.130 71.590 ;
        RECT 23.320 71.170 23.740 71.590 ;
        RECT 23.930 71.170 24.350 71.590 ;
        RECT 25.405 71.170 25.825 71.590 ;
        RECT 26.015 71.170 26.435 71.590 ;
        RECT 26.625 71.170 27.045 71.590 ;
        RECT 27.235 71.170 27.750 71.590 ;
        RECT 36.055 71.170 36.475 71.590 ;
        RECT 36.665 71.170 37.085 71.590 ;
        RECT 37.275 71.170 37.695 71.590 ;
        RECT 37.885 71.170 38.400 71.590 ;
        RECT 39.200 71.170 39.715 71.590 ;
        RECT 39.905 71.170 40.325 71.590 ;
        RECT 40.515 71.170 40.935 71.590 ;
        RECT 41.125 71.170 41.545 71.590 ;
        RECT 47.580 71.170 48.095 71.590 ;
        RECT 48.285 71.170 48.705 71.590 ;
        RECT 48.895 71.170 49.315 71.590 ;
        RECT 49.505 71.170 49.925 71.590 ;
        RECT 50.990 71.170 51.410 71.590 ;
        RECT 51.600 71.170 52.020 71.590 ;
        RECT 52.210 71.170 52.630 71.590 ;
        RECT 52.820 71.170 53.240 71.590 ;
        RECT 53.430 71.170 53.850 71.590 ;
        RECT 54.905 71.170 55.325 71.590 ;
        RECT 55.515 71.170 55.935 71.590 ;
        RECT 56.125 71.170 56.545 71.590 ;
        RECT 56.735 71.170 57.250 71.590 ;
        RECT 65.555 71.170 65.975 71.590 ;
        RECT 66.165 71.170 66.585 71.590 ;
        RECT 66.775 71.170 67.195 71.590 ;
        RECT 67.385 71.170 67.900 71.590 ;
        RECT 68.700 71.170 69.215 71.590 ;
        RECT 69.405 71.170 69.825 71.590 ;
        RECT 70.015 71.170 70.435 71.590 ;
        RECT 70.625 71.170 71.045 71.590 ;
        RECT 77.080 71.170 77.595 71.590 ;
        RECT 77.785 71.170 78.205 71.590 ;
        RECT 78.395 71.170 78.815 71.590 ;
        RECT 79.005 71.170 79.425 71.590 ;
        RECT 80.490 71.170 80.910 71.590 ;
        RECT 81.100 71.170 81.520 71.590 ;
        RECT 81.710 71.170 82.130 71.590 ;
        RECT 82.320 71.170 82.740 71.590 ;
        RECT 82.930 71.170 83.350 71.590 ;
        RECT 84.405 71.170 84.825 71.590 ;
        RECT 85.015 71.170 85.435 71.590 ;
        RECT 85.625 71.170 86.045 71.590 ;
        RECT 86.235 71.170 86.750 71.590 ;
        RECT 95.055 71.170 95.475 71.590 ;
        RECT 95.665 71.170 96.085 71.590 ;
        RECT 96.275 71.170 96.695 71.590 ;
        RECT 96.885 71.170 97.400 71.590 ;
        RECT 98.200 71.170 98.715 71.590 ;
        RECT 98.905 71.170 99.325 71.590 ;
        RECT 99.515 71.170 99.935 71.590 ;
        RECT 100.125 71.170 100.545 71.590 ;
        RECT 106.580 71.170 107.095 71.590 ;
        RECT 107.285 71.170 107.705 71.590 ;
        RECT 107.895 71.170 108.315 71.590 ;
        RECT 108.505 71.170 108.925 71.590 ;
        RECT 109.990 71.170 110.410 71.590 ;
        RECT 110.600 71.170 111.020 71.590 ;
        RECT 111.210 71.170 111.630 71.590 ;
        RECT 111.820 71.170 112.240 71.590 ;
        RECT 112.430 71.170 112.850 71.590 ;
        RECT 113.905 71.170 114.325 71.590 ;
        RECT 114.515 71.170 114.935 71.590 ;
        RECT 115.125 71.170 115.545 71.590 ;
        RECT 115.735 71.170 116.250 71.590 ;
        RECT 124.555 71.170 124.975 71.590 ;
        RECT 125.165 71.170 125.585 71.590 ;
        RECT 125.775 71.170 126.195 71.590 ;
        RECT 126.385 71.170 126.900 71.590 ;
        RECT 127.700 71.170 128.215 71.590 ;
        RECT 128.405 71.170 128.825 71.590 ;
        RECT 129.015 71.170 129.435 71.590 ;
        RECT 129.625 71.170 130.045 71.590 ;
        RECT 136.080 71.170 136.595 71.590 ;
        RECT 136.785 71.170 137.205 71.590 ;
        RECT 137.395 71.170 137.815 71.590 ;
        RECT 138.005 71.170 138.425 71.590 ;
        RECT 139.490 71.170 139.910 71.590 ;
        RECT 140.100 71.170 140.520 71.590 ;
        RECT 140.710 71.170 141.130 71.590 ;
        RECT 141.320 71.170 141.740 71.590 ;
        RECT 141.930 71.170 142.350 71.590 ;
        RECT 143.405 71.170 143.825 71.590 ;
        RECT 144.015 71.170 144.435 71.590 ;
        RECT 144.625 71.170 145.045 71.590 ;
        RECT 145.235 71.170 145.750 71.590 ;
        RECT 154.055 71.170 154.475 71.590 ;
        RECT 154.665 71.170 155.085 71.590 ;
        RECT 155.275 71.170 155.695 71.590 ;
        RECT 155.885 71.170 156.400 71.590 ;
        RECT 157.200 71.170 157.715 71.590 ;
        RECT 157.905 71.170 158.325 71.590 ;
        RECT 158.515 71.170 158.935 71.590 ;
        RECT 159.125 71.170 159.545 71.590 ;
        RECT 18.830 64.120 19.840 65.060 ;
        RECT 28.910 68.450 29.425 68.870 ;
        RECT 29.615 68.450 30.035 68.870 ;
        RECT 30.225 68.450 30.645 68.870 ;
        RECT 30.835 68.450 31.255 68.870 ;
        RECT 32.055 68.450 32.475 68.870 ;
        RECT 32.665 68.450 33.085 68.870 ;
        RECT 33.275 68.450 33.695 68.870 ;
        RECT 33.885 68.450 34.400 68.870 ;
        RECT 24.860 64.280 25.680 64.880 ;
        RECT 36.330 64.290 36.780 64.880 ;
        RECT 36.970 64.290 38.000 64.880 ;
        RECT 44.290 68.450 44.710 68.870 ;
        RECT 44.900 68.450 45.320 68.870 ;
        RECT 45.510 68.450 45.930 68.870 ;
        RECT 42.865 64.225 43.485 64.945 ;
        RECT 30.400 61.620 31.000 62.220 ;
        RECT 31.200 61.620 31.800 62.220 ;
        RECT 32.000 61.620 32.600 62.220 ;
        RECT 32.800 61.530 33.500 62.220 ;
        RECT 33.700 61.530 34.340 62.160 ;
        RECT 18.080 57.570 18.595 57.990 ;
        RECT 18.785 57.570 19.205 57.990 ;
        RECT 19.395 57.570 19.815 57.990 ;
        RECT 20.005 57.570 20.425 57.990 ;
        RECT 21.405 57.570 21.825 57.990 ;
        RECT 22.015 57.570 22.435 57.990 ;
        RECT 22.625 57.570 23.045 57.990 ;
        RECT 23.235 57.570 23.750 57.990 ;
        RECT 36.665 57.570 37.085 57.990 ;
        RECT 37.275 57.570 37.695 57.990 ;
        RECT 37.885 57.570 38.305 57.990 ;
        RECT 40.965 61.560 41.465 62.160 ;
        RECT 48.330 64.120 49.340 65.060 ;
        RECT 58.410 68.450 58.925 68.870 ;
        RECT 59.115 68.450 59.535 68.870 ;
        RECT 59.725 68.450 60.145 68.870 ;
        RECT 60.335 68.450 60.755 68.870 ;
        RECT 61.555 68.450 61.975 68.870 ;
        RECT 62.165 68.450 62.585 68.870 ;
        RECT 62.775 68.450 63.195 68.870 ;
        RECT 63.385 68.450 63.900 68.870 ;
        RECT 54.360 64.280 55.180 64.880 ;
        RECT 44.030 61.610 44.980 62.110 ;
        RECT 45.180 61.610 45.580 62.110 ;
        RECT 65.830 64.290 66.280 64.880 ;
        RECT 66.470 64.290 67.500 64.880 ;
        RECT 73.790 68.450 74.210 68.870 ;
        RECT 74.400 68.450 74.820 68.870 ;
        RECT 75.010 68.450 75.430 68.870 ;
        RECT 72.365 64.225 72.985 64.945 ;
        RECT 59.900 61.620 60.500 62.220 ;
        RECT 60.700 61.620 61.300 62.220 ;
        RECT 61.500 61.620 62.100 62.220 ;
        RECT 62.300 61.530 63.000 62.220 ;
        RECT 63.200 61.530 63.840 62.160 ;
        RECT 47.580 57.570 48.095 57.990 ;
        RECT 48.285 57.570 48.705 57.990 ;
        RECT 48.895 57.570 49.315 57.990 ;
        RECT 49.505 57.570 49.925 57.990 ;
        RECT 50.905 57.570 51.325 57.990 ;
        RECT 51.515 57.570 51.935 57.990 ;
        RECT 52.125 57.570 52.545 57.990 ;
        RECT 52.735 57.570 53.250 57.990 ;
        RECT 66.165 57.570 66.585 57.990 ;
        RECT 66.775 57.570 67.195 57.990 ;
        RECT 67.385 57.570 67.805 57.990 ;
        RECT 70.465 61.560 70.965 62.160 ;
        RECT 77.830 64.120 78.840 65.060 ;
        RECT 87.910 68.450 88.425 68.870 ;
        RECT 88.615 68.450 89.035 68.870 ;
        RECT 89.225 68.450 89.645 68.870 ;
        RECT 89.835 68.450 90.255 68.870 ;
        RECT 91.055 68.450 91.475 68.870 ;
        RECT 91.665 68.450 92.085 68.870 ;
        RECT 92.275 68.450 92.695 68.870 ;
        RECT 92.885 68.450 93.400 68.870 ;
        RECT 83.860 64.280 84.680 64.880 ;
        RECT 73.530 61.610 74.480 62.110 ;
        RECT 74.680 61.610 75.080 62.110 ;
        RECT 95.330 64.290 95.780 64.880 ;
        RECT 95.970 64.290 97.000 64.880 ;
        RECT 103.290 68.450 103.710 68.870 ;
        RECT 103.900 68.450 104.320 68.870 ;
        RECT 104.510 68.450 104.930 68.870 ;
        RECT 101.865 64.225 102.485 64.945 ;
        RECT 89.400 61.620 90.000 62.220 ;
        RECT 90.200 61.620 90.800 62.220 ;
        RECT 91.000 61.620 91.600 62.220 ;
        RECT 91.800 61.530 92.500 62.220 ;
        RECT 92.700 61.530 93.340 62.160 ;
        RECT 77.080 57.570 77.595 57.990 ;
        RECT 77.785 57.570 78.205 57.990 ;
        RECT 78.395 57.570 78.815 57.990 ;
        RECT 79.005 57.570 79.425 57.990 ;
        RECT 80.405 57.570 80.825 57.990 ;
        RECT 81.015 57.570 81.435 57.990 ;
        RECT 81.625 57.570 82.045 57.990 ;
        RECT 82.235 57.570 82.750 57.990 ;
        RECT 95.665 57.570 96.085 57.990 ;
        RECT 96.275 57.570 96.695 57.990 ;
        RECT 96.885 57.570 97.305 57.990 ;
        RECT 99.965 61.560 100.465 62.160 ;
        RECT 107.330 64.120 108.340 65.060 ;
        RECT 117.410 68.450 117.925 68.870 ;
        RECT 118.115 68.450 118.535 68.870 ;
        RECT 118.725 68.450 119.145 68.870 ;
        RECT 119.335 68.450 119.755 68.870 ;
        RECT 120.555 68.450 120.975 68.870 ;
        RECT 121.165 68.450 121.585 68.870 ;
        RECT 121.775 68.450 122.195 68.870 ;
        RECT 122.385 68.450 122.900 68.870 ;
        RECT 113.360 64.280 114.180 64.880 ;
        RECT 103.030 61.610 103.980 62.110 ;
        RECT 104.180 61.610 104.580 62.110 ;
        RECT 124.830 64.290 125.280 64.880 ;
        RECT 125.470 64.290 126.500 64.880 ;
        RECT 132.790 68.450 133.210 68.870 ;
        RECT 133.400 68.450 133.820 68.870 ;
        RECT 134.010 68.450 134.430 68.870 ;
        RECT 131.365 64.225 131.985 64.945 ;
        RECT 118.900 61.620 119.500 62.220 ;
        RECT 119.700 61.620 120.300 62.220 ;
        RECT 120.500 61.620 121.100 62.220 ;
        RECT 121.300 61.530 122.000 62.220 ;
        RECT 122.200 61.530 122.840 62.160 ;
        RECT 106.580 57.570 107.095 57.990 ;
        RECT 107.285 57.570 107.705 57.990 ;
        RECT 107.895 57.570 108.315 57.990 ;
        RECT 108.505 57.570 108.925 57.990 ;
        RECT 109.905 57.570 110.325 57.990 ;
        RECT 110.515 57.570 110.935 57.990 ;
        RECT 111.125 57.570 111.545 57.990 ;
        RECT 111.735 57.570 112.250 57.990 ;
        RECT 125.165 57.570 125.585 57.990 ;
        RECT 125.775 57.570 126.195 57.990 ;
        RECT 126.385 57.570 126.805 57.990 ;
        RECT 129.465 61.560 129.965 62.160 ;
        RECT 136.830 64.120 137.840 65.060 ;
        RECT 146.910 68.450 147.425 68.870 ;
        RECT 147.615 68.450 148.035 68.870 ;
        RECT 148.225 68.450 148.645 68.870 ;
        RECT 148.835 68.450 149.255 68.870 ;
        RECT 150.055 68.450 150.475 68.870 ;
        RECT 150.665 68.450 151.085 68.870 ;
        RECT 151.275 68.450 151.695 68.870 ;
        RECT 151.885 68.450 152.400 68.870 ;
        RECT 142.860 64.280 143.680 64.880 ;
        RECT 132.530 61.610 133.480 62.110 ;
        RECT 133.680 61.610 134.080 62.110 ;
        RECT 154.330 64.290 154.780 64.880 ;
        RECT 154.970 64.290 156.000 64.880 ;
        RECT 162.290 68.450 162.710 68.870 ;
        RECT 162.900 68.450 163.320 68.870 ;
        RECT 163.510 68.450 163.930 68.870 ;
        RECT 160.865 64.225 161.485 64.945 ;
        RECT 148.400 61.620 149.000 62.220 ;
        RECT 149.200 61.620 149.800 62.220 ;
        RECT 150.000 61.620 150.600 62.220 ;
        RECT 150.800 61.530 151.500 62.220 ;
        RECT 151.700 61.530 152.340 62.160 ;
        RECT 136.080 57.570 136.595 57.990 ;
        RECT 136.785 57.570 137.205 57.990 ;
        RECT 137.395 57.570 137.815 57.990 ;
        RECT 138.005 57.570 138.425 57.990 ;
        RECT 139.405 57.570 139.825 57.990 ;
        RECT 140.015 57.570 140.435 57.990 ;
        RECT 140.625 57.570 141.045 57.990 ;
        RECT 141.235 57.570 141.750 57.990 ;
        RECT 154.665 57.570 155.085 57.990 ;
        RECT 155.275 57.570 155.695 57.990 ;
        RECT 155.885 57.570 156.305 57.990 ;
        RECT 158.965 61.560 159.465 62.160 ;
        RECT 162.030 61.610 162.980 62.110 ;
        RECT 163.180 61.610 163.580 62.110 ;
        RECT 24.730 54.850 25.245 55.270 ;
        RECT 25.435 54.850 25.855 55.270 ;
        RECT 26.045 54.850 26.465 55.270 ;
        RECT 26.655 54.850 27.075 55.270 ;
        RECT 28.130 54.850 28.550 55.270 ;
        RECT 28.740 54.850 29.160 55.270 ;
        RECT 29.350 54.850 29.770 55.270 ;
        RECT 29.960 54.850 30.380 55.270 ;
        RECT 30.570 54.850 30.990 55.270 ;
        RECT 32.055 54.850 32.475 55.270 ;
        RECT 32.665 54.850 33.085 55.270 ;
        RECT 33.275 54.850 33.695 55.270 ;
        RECT 33.885 54.850 34.400 55.270 ;
        RECT 41.150 54.850 41.560 55.270 ;
        RECT 41.760 54.850 42.170 55.270 ;
        RECT 42.370 54.850 42.785 55.270 ;
        RECT 44.195 54.850 44.615 55.270 ;
        RECT 44.805 54.850 45.225 55.270 ;
        RECT 45.415 54.850 45.930 55.270 ;
        RECT 54.230 54.850 54.745 55.270 ;
        RECT 54.935 54.850 55.355 55.270 ;
        RECT 55.545 54.850 55.965 55.270 ;
        RECT 56.155 54.850 56.575 55.270 ;
        RECT 57.630 54.850 58.050 55.270 ;
        RECT 58.240 54.850 58.660 55.270 ;
        RECT 58.850 54.850 59.270 55.270 ;
        RECT 59.460 54.850 59.880 55.270 ;
        RECT 60.070 54.850 60.490 55.270 ;
        RECT 61.555 54.850 61.975 55.270 ;
        RECT 62.165 54.850 62.585 55.270 ;
        RECT 62.775 54.850 63.195 55.270 ;
        RECT 63.385 54.850 63.900 55.270 ;
        RECT 70.650 54.850 71.060 55.270 ;
        RECT 71.260 54.850 71.670 55.270 ;
        RECT 71.870 54.850 72.285 55.270 ;
        RECT 73.695 54.850 74.115 55.270 ;
        RECT 74.305 54.850 74.725 55.270 ;
        RECT 74.915 54.850 75.430 55.270 ;
        RECT 83.730 54.850 84.245 55.270 ;
        RECT 84.435 54.850 84.855 55.270 ;
        RECT 85.045 54.850 85.465 55.270 ;
        RECT 85.655 54.850 86.075 55.270 ;
        RECT 87.130 54.850 87.550 55.270 ;
        RECT 87.740 54.850 88.160 55.270 ;
        RECT 88.350 54.850 88.770 55.270 ;
        RECT 88.960 54.850 89.380 55.270 ;
        RECT 89.570 54.850 89.990 55.270 ;
        RECT 91.055 54.850 91.475 55.270 ;
        RECT 91.665 54.850 92.085 55.270 ;
        RECT 92.275 54.850 92.695 55.270 ;
        RECT 92.885 54.850 93.400 55.270 ;
        RECT 100.150 54.850 100.560 55.270 ;
        RECT 100.760 54.850 101.170 55.270 ;
        RECT 101.370 54.850 101.785 55.270 ;
        RECT 103.195 54.850 103.615 55.270 ;
        RECT 103.805 54.850 104.225 55.270 ;
        RECT 104.415 54.850 104.930 55.270 ;
        RECT 113.230 54.850 113.745 55.270 ;
        RECT 113.935 54.850 114.355 55.270 ;
        RECT 114.545 54.850 114.965 55.270 ;
        RECT 115.155 54.850 115.575 55.270 ;
        RECT 116.630 54.850 117.050 55.270 ;
        RECT 117.240 54.850 117.660 55.270 ;
        RECT 117.850 54.850 118.270 55.270 ;
        RECT 118.460 54.850 118.880 55.270 ;
        RECT 119.070 54.850 119.490 55.270 ;
        RECT 120.555 54.850 120.975 55.270 ;
        RECT 121.165 54.850 121.585 55.270 ;
        RECT 121.775 54.850 122.195 55.270 ;
        RECT 122.385 54.850 122.900 55.270 ;
        RECT 129.650 54.850 130.060 55.270 ;
        RECT 130.260 54.850 130.670 55.270 ;
        RECT 130.870 54.850 131.285 55.270 ;
        RECT 132.695 54.850 133.115 55.270 ;
        RECT 133.305 54.850 133.725 55.270 ;
        RECT 133.915 54.850 134.430 55.270 ;
        RECT 142.730 54.850 143.245 55.270 ;
        RECT 143.435 54.850 143.855 55.270 ;
        RECT 144.045 54.850 144.465 55.270 ;
        RECT 144.655 54.850 145.075 55.270 ;
        RECT 146.130 54.850 146.550 55.270 ;
        RECT 146.740 54.850 147.160 55.270 ;
        RECT 147.350 54.850 147.770 55.270 ;
        RECT 147.960 54.850 148.380 55.270 ;
        RECT 148.570 54.850 148.990 55.270 ;
        RECT 150.055 54.850 150.475 55.270 ;
        RECT 150.665 54.850 151.085 55.270 ;
        RECT 151.275 54.850 151.695 55.270 ;
        RECT 151.885 54.850 152.400 55.270 ;
        RECT 159.150 54.850 159.560 55.270 ;
        RECT 159.760 54.850 160.170 55.270 ;
        RECT 160.370 54.850 160.785 55.270 ;
        RECT 162.195 54.850 162.615 55.270 ;
        RECT 162.805 54.850 163.225 55.270 ;
        RECT 163.415 54.850 163.930 55.270 ;
        RECT 172.125 59.485 172.295 59.655 ;
        RECT 172.485 59.485 172.655 59.655 ;
        RECT 172.845 59.485 173.015 59.655 ;
        RECT 173.205 59.485 173.375 59.655 ;
        RECT 173.565 59.485 173.735 59.655 ;
        RECT 175.255 59.025 175.425 59.195 ;
        RECT 175.615 59.025 175.785 59.195 ;
        RECT 175.975 59.025 176.145 59.195 ;
        RECT 176.335 59.025 176.505 59.195 ;
        RECT 176.695 59.025 176.865 59.195 ;
        RECT 172.125 54.965 172.295 55.135 ;
        RECT 172.485 54.965 172.655 55.135 ;
        RECT 172.845 54.965 173.015 55.135 ;
        RECT 173.205 54.965 173.375 55.135 ;
        RECT 173.565 54.965 173.735 55.135 ;
        RECT 175.255 54.505 175.425 54.675 ;
        RECT 175.615 54.505 175.785 54.675 ;
        RECT 175.975 54.505 176.145 54.675 ;
        RECT 176.335 54.505 176.505 54.675 ;
        RECT 176.695 54.505 176.865 54.675 ;
        RECT 3.185 49.410 3.605 49.830 ;
        RECT 3.795 49.410 4.215 49.830 ;
        RECT 4.405 49.410 4.825 49.830 ;
        RECT 6.240 49.410 6.650 49.830 ;
        RECT 6.850 49.410 7.260 49.830 ;
        RECT 7.460 49.410 7.970 49.830 ;
        RECT 14.010 49.410 14.525 49.830 ;
        RECT 14.715 49.410 15.135 49.830 ;
        RECT 15.325 49.410 15.745 49.830 ;
        RECT 15.935 49.410 16.355 49.830 ;
        RECT 17.420 49.410 17.840 49.830 ;
        RECT 18.030 49.410 18.450 49.830 ;
        RECT 18.640 49.410 19.060 49.830 ;
        RECT 19.250 49.410 19.670 49.830 ;
        RECT 19.860 49.410 20.280 49.830 ;
        RECT 21.335 49.410 21.755 49.830 ;
        RECT 21.945 49.410 22.365 49.830 ;
        RECT 22.555 49.410 22.975 49.830 ;
        RECT 23.165 49.410 23.680 49.830 ;
        RECT 32.685 49.410 33.105 49.830 ;
        RECT 33.295 49.410 33.715 49.830 ;
        RECT 33.905 49.410 34.325 49.830 ;
        RECT 35.740 49.410 36.150 49.830 ;
        RECT 36.350 49.410 36.760 49.830 ;
        RECT 36.960 49.410 37.470 49.830 ;
        RECT 43.510 49.410 44.025 49.830 ;
        RECT 44.215 49.410 44.635 49.830 ;
        RECT 44.825 49.410 45.245 49.830 ;
        RECT 45.435 49.410 45.855 49.830 ;
        RECT 46.920 49.410 47.340 49.830 ;
        RECT 47.530 49.410 47.950 49.830 ;
        RECT 48.140 49.410 48.560 49.830 ;
        RECT 48.750 49.410 49.170 49.830 ;
        RECT 49.360 49.410 49.780 49.830 ;
        RECT 50.835 49.410 51.255 49.830 ;
        RECT 51.445 49.410 51.865 49.830 ;
        RECT 52.055 49.410 52.475 49.830 ;
        RECT 52.665 49.410 53.180 49.830 ;
        RECT 62.185 49.410 62.605 49.830 ;
        RECT 62.795 49.410 63.215 49.830 ;
        RECT 63.405 49.410 63.825 49.830 ;
        RECT 65.240 49.410 65.650 49.830 ;
        RECT 65.850 49.410 66.260 49.830 ;
        RECT 66.460 49.410 66.970 49.830 ;
        RECT 73.010 49.410 73.525 49.830 ;
        RECT 73.715 49.410 74.135 49.830 ;
        RECT 74.325 49.410 74.745 49.830 ;
        RECT 74.935 49.410 75.355 49.830 ;
        RECT 76.420 49.410 76.840 49.830 ;
        RECT 77.030 49.410 77.450 49.830 ;
        RECT 77.640 49.410 78.060 49.830 ;
        RECT 78.250 49.410 78.670 49.830 ;
        RECT 78.860 49.410 79.280 49.830 ;
        RECT 80.335 49.410 80.755 49.830 ;
        RECT 80.945 49.410 81.365 49.830 ;
        RECT 81.555 49.410 81.975 49.830 ;
        RECT 82.165 49.410 82.680 49.830 ;
        RECT 91.685 49.410 92.105 49.830 ;
        RECT 92.295 49.410 92.715 49.830 ;
        RECT 92.905 49.410 93.325 49.830 ;
        RECT 94.740 49.410 95.150 49.830 ;
        RECT 95.350 49.410 95.760 49.830 ;
        RECT 95.960 49.410 96.470 49.830 ;
        RECT 102.510 49.410 103.025 49.830 ;
        RECT 103.215 49.410 103.635 49.830 ;
        RECT 103.825 49.410 104.245 49.830 ;
        RECT 104.435 49.410 104.855 49.830 ;
        RECT 105.920 49.410 106.340 49.830 ;
        RECT 106.530 49.410 106.950 49.830 ;
        RECT 107.140 49.410 107.560 49.830 ;
        RECT 107.750 49.410 108.170 49.830 ;
        RECT 108.360 49.410 108.780 49.830 ;
        RECT 109.835 49.410 110.255 49.830 ;
        RECT 110.445 49.410 110.865 49.830 ;
        RECT 111.055 49.410 111.475 49.830 ;
        RECT 111.665 49.410 112.180 49.830 ;
        RECT 121.185 49.410 121.605 49.830 ;
        RECT 121.795 49.410 122.215 49.830 ;
        RECT 122.405 49.410 122.825 49.830 ;
        RECT 124.240 49.410 124.650 49.830 ;
        RECT 124.850 49.410 125.260 49.830 ;
        RECT 125.460 49.410 125.970 49.830 ;
        RECT 132.010 49.410 132.525 49.830 ;
        RECT 132.715 49.410 133.135 49.830 ;
        RECT 133.325 49.410 133.745 49.830 ;
        RECT 133.935 49.410 134.355 49.830 ;
        RECT 135.420 49.410 135.840 49.830 ;
        RECT 136.030 49.410 136.450 49.830 ;
        RECT 136.640 49.410 137.060 49.830 ;
        RECT 137.250 49.410 137.670 49.830 ;
        RECT 137.860 49.410 138.280 49.830 ;
        RECT 139.335 49.410 139.755 49.830 ;
        RECT 139.945 49.410 140.365 49.830 ;
        RECT 140.555 49.410 140.975 49.830 ;
        RECT 141.165 49.410 141.680 49.830 ;
        RECT 150.685 49.410 151.105 49.830 ;
        RECT 151.295 49.410 151.715 49.830 ;
        RECT 151.905 49.410 152.325 49.830 ;
        RECT 153.740 49.410 154.150 49.830 ;
        RECT 154.350 49.410 154.760 49.830 ;
        RECT 154.960 49.410 155.470 49.830 ;
        RECT 161.510 49.410 162.025 49.830 ;
        RECT 162.215 49.410 162.635 49.830 ;
        RECT 162.825 49.410 163.245 49.830 ;
        RECT 163.435 49.410 163.855 49.830 ;
        RECT 164.920 49.410 165.340 49.830 ;
        RECT 165.530 49.410 165.950 49.830 ;
        RECT 166.140 49.410 166.560 49.830 ;
        RECT 166.750 49.410 167.170 49.830 ;
        RECT 167.360 49.410 167.780 49.830 ;
        RECT 168.835 49.410 169.255 49.830 ;
        RECT 169.445 49.410 169.865 49.830 ;
        RECT 170.055 49.410 170.475 49.830 ;
        RECT 170.665 49.410 171.180 49.830 ;
        RECT 2.830 42.570 3.230 43.070 ;
        RECT 3.430 42.570 4.380 43.070 ;
        RECT 6.945 42.520 7.445 43.120 ;
        RECT 10.715 46.690 11.135 47.110 ;
        RECT 11.325 46.690 11.745 47.110 ;
        RECT 11.935 46.690 12.355 47.110 ;
        RECT 25.365 46.690 25.785 47.110 ;
        RECT 25.975 46.690 26.395 47.110 ;
        RECT 26.585 46.690 27.005 47.110 ;
        RECT 27.985 46.690 28.405 47.110 ;
        RECT 28.595 46.690 29.015 47.110 ;
        RECT 29.205 46.690 29.625 47.110 ;
        RECT 29.815 46.690 30.330 47.110 ;
        RECT 14.070 42.520 14.710 43.150 ;
        RECT 14.910 42.460 15.610 43.150 ;
        RECT 15.810 42.460 16.410 43.060 ;
        RECT 16.610 42.460 17.210 43.060 ;
        RECT 17.410 42.460 18.010 43.060 ;
        RECT 4.925 39.735 5.545 40.455 ;
        RECT 3.090 35.810 3.510 36.230 ;
        RECT 3.700 35.810 4.120 36.230 ;
        RECT 4.310 35.810 4.730 36.230 ;
        RECT 10.410 39.800 11.440 40.390 ;
        RECT 11.630 39.800 12.080 40.390 ;
        RECT 32.330 42.570 32.730 43.070 ;
        RECT 32.930 42.570 33.880 43.070 ;
        RECT 14.010 35.810 14.525 36.230 ;
        RECT 14.715 35.810 15.135 36.230 ;
        RECT 15.325 35.810 15.745 36.230 ;
        RECT 15.935 35.810 16.355 36.230 ;
        RECT 17.155 35.810 17.575 36.230 ;
        RECT 17.765 35.810 18.185 36.230 ;
        RECT 18.375 35.810 18.795 36.230 ;
        RECT 18.985 35.810 19.500 36.230 ;
        RECT 28.570 39.620 29.580 40.560 ;
        RECT 36.445 42.520 36.945 43.120 ;
        RECT 40.215 46.690 40.635 47.110 ;
        RECT 40.825 46.690 41.245 47.110 ;
        RECT 41.435 46.690 41.855 47.110 ;
        RECT 54.865 46.690 55.285 47.110 ;
        RECT 55.475 46.690 55.895 47.110 ;
        RECT 56.085 46.690 56.505 47.110 ;
        RECT 57.485 46.690 57.905 47.110 ;
        RECT 58.095 46.690 58.515 47.110 ;
        RECT 58.705 46.690 59.125 47.110 ;
        RECT 59.315 46.690 59.830 47.110 ;
        RECT 43.570 42.520 44.210 43.150 ;
        RECT 44.410 42.460 45.110 43.150 ;
        RECT 45.310 42.460 45.910 43.060 ;
        RECT 46.110 42.460 46.710 43.060 ;
        RECT 46.910 42.460 47.510 43.060 ;
        RECT 34.425 39.735 35.045 40.455 ;
        RECT 32.590 35.810 33.010 36.230 ;
        RECT 33.200 35.810 33.620 36.230 ;
        RECT 33.810 35.810 34.230 36.230 ;
        RECT 39.910 39.800 40.940 40.390 ;
        RECT 41.130 39.800 41.580 40.390 ;
        RECT 61.830 42.570 62.230 43.070 ;
        RECT 62.430 42.570 63.380 43.070 ;
        RECT 43.510 35.810 44.025 36.230 ;
        RECT 44.215 35.810 44.635 36.230 ;
        RECT 44.825 35.810 45.245 36.230 ;
        RECT 45.435 35.810 45.855 36.230 ;
        RECT 46.655 35.810 47.075 36.230 ;
        RECT 47.265 35.810 47.685 36.230 ;
        RECT 47.875 35.810 48.295 36.230 ;
        RECT 48.485 35.810 49.000 36.230 ;
        RECT 58.070 39.620 59.080 40.560 ;
        RECT 65.945 42.520 66.445 43.120 ;
        RECT 69.715 46.690 70.135 47.110 ;
        RECT 70.325 46.690 70.745 47.110 ;
        RECT 70.935 46.690 71.355 47.110 ;
        RECT 84.365 46.690 84.785 47.110 ;
        RECT 84.975 46.690 85.395 47.110 ;
        RECT 85.585 46.690 86.005 47.110 ;
        RECT 86.985 46.690 87.405 47.110 ;
        RECT 87.595 46.690 88.015 47.110 ;
        RECT 88.205 46.690 88.625 47.110 ;
        RECT 88.815 46.690 89.330 47.110 ;
        RECT 73.070 42.520 73.710 43.150 ;
        RECT 73.910 42.460 74.610 43.150 ;
        RECT 74.810 42.460 75.410 43.060 ;
        RECT 75.610 42.460 76.210 43.060 ;
        RECT 76.410 42.460 77.010 43.060 ;
        RECT 63.925 39.735 64.545 40.455 ;
        RECT 62.090 35.810 62.510 36.230 ;
        RECT 62.700 35.810 63.120 36.230 ;
        RECT 63.310 35.810 63.730 36.230 ;
        RECT 69.410 39.800 70.440 40.390 ;
        RECT 70.630 39.800 71.080 40.390 ;
        RECT 91.330 42.570 91.730 43.070 ;
        RECT 91.930 42.570 92.880 43.070 ;
        RECT 73.010 35.810 73.525 36.230 ;
        RECT 73.715 35.810 74.135 36.230 ;
        RECT 74.325 35.810 74.745 36.230 ;
        RECT 74.935 35.810 75.355 36.230 ;
        RECT 76.155 35.810 76.575 36.230 ;
        RECT 76.765 35.810 77.185 36.230 ;
        RECT 77.375 35.810 77.795 36.230 ;
        RECT 77.985 35.810 78.500 36.230 ;
        RECT 87.570 39.620 88.580 40.560 ;
        RECT 95.445 42.520 95.945 43.120 ;
        RECT 99.215 46.690 99.635 47.110 ;
        RECT 99.825 46.690 100.245 47.110 ;
        RECT 100.435 46.690 100.855 47.110 ;
        RECT 113.865 46.690 114.285 47.110 ;
        RECT 114.475 46.690 114.895 47.110 ;
        RECT 115.085 46.690 115.505 47.110 ;
        RECT 116.485 46.690 116.905 47.110 ;
        RECT 117.095 46.690 117.515 47.110 ;
        RECT 117.705 46.690 118.125 47.110 ;
        RECT 118.315 46.690 118.830 47.110 ;
        RECT 102.570 42.520 103.210 43.150 ;
        RECT 103.410 42.460 104.110 43.150 ;
        RECT 104.310 42.460 104.910 43.060 ;
        RECT 105.110 42.460 105.710 43.060 ;
        RECT 105.910 42.460 106.510 43.060 ;
        RECT 93.425 39.735 94.045 40.455 ;
        RECT 91.590 35.810 92.010 36.230 ;
        RECT 92.200 35.810 92.620 36.230 ;
        RECT 92.810 35.810 93.230 36.230 ;
        RECT 98.910 39.800 99.940 40.390 ;
        RECT 100.130 39.800 100.580 40.390 ;
        RECT 120.830 42.570 121.230 43.070 ;
        RECT 121.430 42.570 122.380 43.070 ;
        RECT 102.510 35.810 103.025 36.230 ;
        RECT 103.215 35.810 103.635 36.230 ;
        RECT 103.825 35.810 104.245 36.230 ;
        RECT 104.435 35.810 104.855 36.230 ;
        RECT 105.655 35.810 106.075 36.230 ;
        RECT 106.265 35.810 106.685 36.230 ;
        RECT 106.875 35.810 107.295 36.230 ;
        RECT 107.485 35.810 108.000 36.230 ;
        RECT 117.070 39.620 118.080 40.560 ;
        RECT 124.945 42.520 125.445 43.120 ;
        RECT 128.715 46.690 129.135 47.110 ;
        RECT 129.325 46.690 129.745 47.110 ;
        RECT 129.935 46.690 130.355 47.110 ;
        RECT 143.365 46.690 143.785 47.110 ;
        RECT 143.975 46.690 144.395 47.110 ;
        RECT 144.585 46.690 145.005 47.110 ;
        RECT 145.985 46.690 146.405 47.110 ;
        RECT 146.595 46.690 147.015 47.110 ;
        RECT 147.205 46.690 147.625 47.110 ;
        RECT 147.815 46.690 148.330 47.110 ;
        RECT 132.070 42.520 132.710 43.150 ;
        RECT 132.910 42.460 133.610 43.150 ;
        RECT 133.810 42.460 134.410 43.060 ;
        RECT 134.610 42.460 135.210 43.060 ;
        RECT 135.410 42.460 136.010 43.060 ;
        RECT 122.925 39.735 123.545 40.455 ;
        RECT 121.090 35.810 121.510 36.230 ;
        RECT 121.700 35.810 122.120 36.230 ;
        RECT 122.310 35.810 122.730 36.230 ;
        RECT 128.410 39.800 129.440 40.390 ;
        RECT 129.630 39.800 130.080 40.390 ;
        RECT 150.330 42.570 150.730 43.070 ;
        RECT 150.930 42.570 151.880 43.070 ;
        RECT 132.010 35.810 132.525 36.230 ;
        RECT 132.715 35.810 133.135 36.230 ;
        RECT 133.325 35.810 133.745 36.230 ;
        RECT 133.935 35.810 134.355 36.230 ;
        RECT 135.155 35.810 135.575 36.230 ;
        RECT 135.765 35.810 136.185 36.230 ;
        RECT 136.375 35.810 136.795 36.230 ;
        RECT 136.985 35.810 137.500 36.230 ;
        RECT 146.570 39.620 147.580 40.560 ;
        RECT 154.445 42.520 154.945 43.120 ;
        RECT 158.215 46.690 158.635 47.110 ;
        RECT 158.825 46.690 159.245 47.110 ;
        RECT 159.435 46.690 159.855 47.110 ;
        RECT 172.865 46.690 173.285 47.110 ;
        RECT 173.475 46.690 173.895 47.110 ;
        RECT 174.085 46.690 174.505 47.110 ;
        RECT 175.485 46.690 175.905 47.110 ;
        RECT 176.095 46.690 176.515 47.110 ;
        RECT 176.705 46.690 177.125 47.110 ;
        RECT 177.315 46.690 177.830 47.110 ;
        RECT 161.570 42.520 162.210 43.150 ;
        RECT 162.410 42.460 163.110 43.150 ;
        RECT 163.310 42.460 163.910 43.060 ;
        RECT 164.110 42.460 164.710 43.060 ;
        RECT 164.910 42.460 165.510 43.060 ;
        RECT 152.425 39.735 153.045 40.455 ;
        RECT 150.590 35.810 151.010 36.230 ;
        RECT 151.200 35.810 151.620 36.230 ;
        RECT 151.810 35.810 152.230 36.230 ;
        RECT 157.910 39.800 158.940 40.390 ;
        RECT 159.130 39.800 159.580 40.390 ;
        RECT 161.510 35.810 162.025 36.230 ;
        RECT 162.215 35.810 162.635 36.230 ;
        RECT 162.825 35.810 163.245 36.230 ;
        RECT 163.435 35.810 163.855 36.230 ;
        RECT 164.655 35.810 165.075 36.230 ;
        RECT 165.265 35.810 165.685 36.230 ;
        RECT 165.875 35.810 166.295 36.230 ;
        RECT 166.485 35.810 167.000 36.230 ;
        RECT 176.070 39.620 177.080 40.560 ;
        RECT 6.865 33.090 7.285 33.510 ;
        RECT 7.475 33.090 7.895 33.510 ;
        RECT 8.085 33.090 8.505 33.510 ;
        RECT 8.695 33.090 9.210 33.510 ;
        RECT 10.010 33.090 10.525 33.510 ;
        RECT 10.715 33.090 11.135 33.510 ;
        RECT 11.325 33.090 11.745 33.510 ;
        RECT 11.935 33.090 12.355 33.510 ;
        RECT 20.660 33.090 21.175 33.510 ;
        RECT 21.365 33.090 21.785 33.510 ;
        RECT 21.975 33.090 22.395 33.510 ;
        RECT 22.585 33.090 23.005 33.510 ;
        RECT 24.060 33.090 24.480 33.510 ;
        RECT 24.670 33.090 25.090 33.510 ;
        RECT 25.280 33.090 25.700 33.510 ;
        RECT 25.890 33.090 26.310 33.510 ;
        RECT 26.500 33.090 26.920 33.510 ;
        RECT 27.985 33.090 28.405 33.510 ;
        RECT 28.595 33.090 29.015 33.510 ;
        RECT 29.205 33.090 29.625 33.510 ;
        RECT 29.815 33.090 30.330 33.510 ;
        RECT 36.365 33.090 36.785 33.510 ;
        RECT 36.975 33.090 37.395 33.510 ;
        RECT 37.585 33.090 38.005 33.510 ;
        RECT 38.195 33.090 38.710 33.510 ;
        RECT 39.510 33.090 40.025 33.510 ;
        RECT 40.215 33.090 40.635 33.510 ;
        RECT 40.825 33.090 41.245 33.510 ;
        RECT 41.435 33.090 41.855 33.510 ;
        RECT 50.160 33.090 50.675 33.510 ;
        RECT 50.865 33.090 51.285 33.510 ;
        RECT 51.475 33.090 51.895 33.510 ;
        RECT 52.085 33.090 52.505 33.510 ;
        RECT 53.560 33.090 53.980 33.510 ;
        RECT 54.170 33.090 54.590 33.510 ;
        RECT 54.780 33.090 55.200 33.510 ;
        RECT 55.390 33.090 55.810 33.510 ;
        RECT 56.000 33.090 56.420 33.510 ;
        RECT 57.485 33.090 57.905 33.510 ;
        RECT 58.095 33.090 58.515 33.510 ;
        RECT 58.705 33.090 59.125 33.510 ;
        RECT 59.315 33.090 59.830 33.510 ;
        RECT 65.865 33.090 66.285 33.510 ;
        RECT 66.475 33.090 66.895 33.510 ;
        RECT 67.085 33.090 67.505 33.510 ;
        RECT 67.695 33.090 68.210 33.510 ;
        RECT 69.010 33.090 69.525 33.510 ;
        RECT 69.715 33.090 70.135 33.510 ;
        RECT 70.325 33.090 70.745 33.510 ;
        RECT 70.935 33.090 71.355 33.510 ;
        RECT 79.660 33.090 80.175 33.510 ;
        RECT 80.365 33.090 80.785 33.510 ;
        RECT 80.975 33.090 81.395 33.510 ;
        RECT 81.585 33.090 82.005 33.510 ;
        RECT 83.060 33.090 83.480 33.510 ;
        RECT 83.670 33.090 84.090 33.510 ;
        RECT 84.280 33.090 84.700 33.510 ;
        RECT 84.890 33.090 85.310 33.510 ;
        RECT 85.500 33.090 85.920 33.510 ;
        RECT 86.985 33.090 87.405 33.510 ;
        RECT 87.595 33.090 88.015 33.510 ;
        RECT 88.205 33.090 88.625 33.510 ;
        RECT 88.815 33.090 89.330 33.510 ;
        RECT 95.365 33.090 95.785 33.510 ;
        RECT 95.975 33.090 96.395 33.510 ;
        RECT 96.585 33.090 97.005 33.510 ;
        RECT 97.195 33.090 97.710 33.510 ;
        RECT 98.510 33.090 99.025 33.510 ;
        RECT 99.215 33.090 99.635 33.510 ;
        RECT 99.825 33.090 100.245 33.510 ;
        RECT 100.435 33.090 100.855 33.510 ;
        RECT 109.160 33.090 109.675 33.510 ;
        RECT 109.865 33.090 110.285 33.510 ;
        RECT 110.475 33.090 110.895 33.510 ;
        RECT 111.085 33.090 111.505 33.510 ;
        RECT 112.560 33.090 112.980 33.510 ;
        RECT 113.170 33.090 113.590 33.510 ;
        RECT 113.780 33.090 114.200 33.510 ;
        RECT 114.390 33.090 114.810 33.510 ;
        RECT 115.000 33.090 115.420 33.510 ;
        RECT 116.485 33.090 116.905 33.510 ;
        RECT 117.095 33.090 117.515 33.510 ;
        RECT 117.705 33.090 118.125 33.510 ;
        RECT 118.315 33.090 118.830 33.510 ;
        RECT 124.865 33.090 125.285 33.510 ;
        RECT 125.475 33.090 125.895 33.510 ;
        RECT 126.085 33.090 126.505 33.510 ;
        RECT 126.695 33.090 127.210 33.510 ;
        RECT 128.010 33.090 128.525 33.510 ;
        RECT 128.715 33.090 129.135 33.510 ;
        RECT 129.325 33.090 129.745 33.510 ;
        RECT 129.935 33.090 130.355 33.510 ;
        RECT 138.660 33.090 139.175 33.510 ;
        RECT 139.365 33.090 139.785 33.510 ;
        RECT 139.975 33.090 140.395 33.510 ;
        RECT 140.585 33.090 141.005 33.510 ;
        RECT 142.060 33.090 142.480 33.510 ;
        RECT 142.670 33.090 143.090 33.510 ;
        RECT 143.280 33.090 143.700 33.510 ;
        RECT 143.890 33.090 144.310 33.510 ;
        RECT 144.500 33.090 144.920 33.510 ;
        RECT 145.985 33.090 146.405 33.510 ;
        RECT 146.595 33.090 147.015 33.510 ;
        RECT 147.205 33.090 147.625 33.510 ;
        RECT 147.815 33.090 148.330 33.510 ;
        RECT 154.365 33.090 154.785 33.510 ;
        RECT 154.975 33.090 155.395 33.510 ;
        RECT 155.585 33.090 156.005 33.510 ;
        RECT 156.195 33.090 156.710 33.510 ;
        RECT 157.510 33.090 158.025 33.510 ;
        RECT 158.215 33.090 158.635 33.510 ;
        RECT 158.825 33.090 159.245 33.510 ;
        RECT 159.435 33.090 159.855 33.510 ;
        RECT 168.160 33.090 168.675 33.510 ;
        RECT 168.865 33.090 169.285 33.510 ;
        RECT 169.475 33.090 169.895 33.510 ;
        RECT 170.085 33.090 170.505 33.510 ;
        RECT 171.560 33.090 171.980 33.510 ;
        RECT 172.170 33.090 172.590 33.510 ;
        RECT 172.780 33.090 173.200 33.510 ;
        RECT 173.390 33.090 173.810 33.510 ;
        RECT 174.000 33.090 174.420 33.510 ;
        RECT 175.485 33.090 175.905 33.510 ;
        RECT 176.095 33.090 176.515 33.510 ;
        RECT 176.705 33.090 177.125 33.510 ;
        RECT 177.315 33.090 177.830 33.510 ;
        RECT 36.100 31.100 36.400 31.400 ;
        RECT 36.600 31.100 36.900 31.400 ;
        RECT 37.100 31.100 37.400 31.400 ;
        RECT 37.600 31.100 37.900 31.400 ;
        RECT 72.100 31.100 72.400 31.400 ;
        RECT 72.600 31.100 72.900 31.400 ;
        RECT 73.100 31.100 73.400 31.400 ;
        RECT 73.600 31.100 73.900 31.400 ;
        RECT 108.100 31.100 108.400 31.400 ;
        RECT 108.600 31.100 108.900 31.400 ;
        RECT 109.100 31.100 109.400 31.400 ;
        RECT 109.600 31.100 109.900 31.400 ;
        RECT 144.100 31.100 144.400 31.400 ;
        RECT 144.600 31.100 144.900 31.400 ;
        RECT 145.100 31.100 145.400 31.400 ;
        RECT 145.600 31.100 145.900 31.400 ;
      LAYER met1 ;
        RECT 36.000 73.000 38.000 73.500 ;
        RECT 72.000 73.000 74.000 73.500 ;
        RECT 108.000 73.000 110.000 73.500 ;
        RECT 144.000 73.000 146.000 73.500 ;
        RECT 15.790 71.140 173.000 71.620 ;
        RECT 15.510 68.420 164.900 68.900 ;
        RECT 18.800 64.915 19.930 65.140 ;
        RECT 42.805 64.915 43.545 64.975 ;
        RECT 48.300 64.915 49.430 65.140 ;
        RECT 72.305 64.915 73.045 64.975 ;
        RECT 77.800 64.915 78.930 65.140 ;
        RECT 101.805 64.915 102.545 64.975 ;
        RECT 107.300 64.915 108.430 65.140 ;
        RECT 131.305 64.915 132.045 64.975 ;
        RECT 136.800 64.915 137.930 65.140 ;
        RECT 160.805 64.915 161.545 64.975 ;
        RECT 17.350 64.255 19.930 64.915 ;
        RECT 34.570 64.910 49.430 64.915 ;
        RECT 64.070 64.910 78.930 64.915 ;
        RECT 93.570 64.910 108.430 64.915 ;
        RECT 123.070 64.910 137.930 64.915 ;
        RECT 152.570 64.910 164.950 64.915 ;
        RECT 18.800 64.040 19.930 64.255 ;
        RECT 24.800 64.255 49.430 64.910 ;
        RECT 24.800 64.250 38.060 64.255 ;
        RECT 42.805 64.195 43.545 64.255 ;
        RECT 48.300 64.040 49.430 64.255 ;
        RECT 54.300 64.255 78.930 64.910 ;
        RECT 54.300 64.250 67.560 64.255 ;
        RECT 72.305 64.195 73.045 64.255 ;
        RECT 77.800 64.040 78.930 64.255 ;
        RECT 83.800 64.255 108.430 64.910 ;
        RECT 83.800 64.250 97.060 64.255 ;
        RECT 101.805 64.195 102.545 64.255 ;
        RECT 107.300 64.040 108.430 64.255 ;
        RECT 113.300 64.255 137.930 64.910 ;
        RECT 113.300 64.250 126.560 64.255 ;
        RECT 131.305 64.195 132.045 64.255 ;
        RECT 136.800 64.040 137.930 64.255 ;
        RECT 142.800 64.255 164.950 64.910 ;
        RECT 142.800 64.250 156.060 64.255 ;
        RECT 160.805 64.195 161.545 64.255 ;
        RECT 3.330 62.980 20.000 63.460 ;
        RECT 30.300 62.220 33.600 62.250 ;
        RECT 59.800 62.220 63.100 62.250 ;
        RECT 89.300 62.220 92.600 62.250 ;
        RECT 118.800 62.220 122.100 62.250 ;
        RECT 148.300 62.220 151.600 62.250 ;
        RECT 30.300 62.160 34.400 62.220 ;
        RECT 2.370 61.800 2.710 62.100 ;
        RECT 6.310 62.010 6.730 62.040 ;
        RECT 16.510 62.010 34.400 62.160 ;
        RECT 6.310 61.710 34.400 62.010 ;
        RECT 6.310 61.680 6.730 61.710 ;
        RECT 16.510 61.560 34.400 61.710 ;
        RECT 30.300 61.500 34.400 61.560 ;
        RECT 40.935 62.160 41.495 62.220 ;
        RECT 59.800 62.160 63.900 62.220 ;
        RECT 40.935 61.560 63.900 62.160 ;
        RECT 40.935 61.500 41.495 61.560 ;
        RECT 59.800 61.500 63.900 61.560 ;
        RECT 70.435 62.160 70.995 62.220 ;
        RECT 89.300 62.160 93.400 62.220 ;
        RECT 70.435 61.560 93.400 62.160 ;
        RECT 70.435 61.500 70.995 61.560 ;
        RECT 89.300 61.500 93.400 61.560 ;
        RECT 99.935 62.160 100.495 62.220 ;
        RECT 118.800 62.160 122.900 62.220 ;
        RECT 99.935 61.560 122.900 62.160 ;
        RECT 99.935 61.500 100.495 61.560 ;
        RECT 118.800 61.500 122.900 61.560 ;
        RECT 129.435 62.160 129.995 62.220 ;
        RECT 148.300 62.160 152.400 62.220 ;
        RECT 129.435 61.560 152.400 62.160 ;
        RECT 129.435 61.500 129.995 61.560 ;
        RECT 148.300 61.500 152.400 61.560 ;
        RECT 158.935 62.160 159.495 62.220 ;
        RECT 158.935 61.560 164.950 62.160 ;
        RECT 158.935 61.500 159.495 61.560 ;
        RECT 0.000 60.260 9.475 60.740 ;
        RECT 171.100 60.260 182.000 60.740 ;
        RECT 171.950 59.440 173.910 60.260 ;
        RECT 175.030 58.980 177.090 59.240 ;
        RECT 14.515 57.540 171.950 58.020 ;
        RECT 162.000 57.535 164.000 57.540 ;
        RECT 17.400 55.290 164.900 55.300 ;
        RECT 16.510 54.810 177.040 55.290 ;
        RECT 175.080 54.460 177.040 54.810 ;
        RECT 1.510 49.380 179.950 49.860 ;
        RECT 0.000 46.660 178.955 47.140 ;
        RECT 6.915 43.120 7.475 43.180 ;
        RECT 1.510 42.520 7.475 43.120 ;
        RECT 6.915 42.460 7.475 42.520 ;
        RECT 14.010 43.120 18.110 43.180 ;
        RECT 36.415 43.120 36.975 43.180 ;
        RECT 14.010 42.520 36.975 43.120 ;
        RECT 14.010 42.460 18.110 42.520 ;
        RECT 36.415 42.460 36.975 42.520 ;
        RECT 43.510 43.120 47.610 43.180 ;
        RECT 65.915 43.120 66.475 43.180 ;
        RECT 43.510 42.520 66.475 43.120 ;
        RECT 43.510 42.460 47.610 42.520 ;
        RECT 65.915 42.460 66.475 42.520 ;
        RECT 73.010 43.120 77.110 43.180 ;
        RECT 95.415 43.120 95.975 43.180 ;
        RECT 73.010 42.520 95.975 43.120 ;
        RECT 73.010 42.460 77.110 42.520 ;
        RECT 95.415 42.460 95.975 42.520 ;
        RECT 102.510 43.120 106.610 43.180 ;
        RECT 124.915 43.120 125.475 43.180 ;
        RECT 102.510 42.520 125.475 43.120 ;
        RECT 102.510 42.460 106.610 42.520 ;
        RECT 124.915 42.460 125.475 42.520 ;
        RECT 132.010 43.120 136.110 43.180 ;
        RECT 154.415 43.120 154.975 43.180 ;
        RECT 132.010 42.520 154.975 43.120 ;
        RECT 132.010 42.460 136.110 42.520 ;
        RECT 154.415 42.460 154.975 42.520 ;
        RECT 161.510 43.120 165.610 43.180 ;
        RECT 161.510 42.520 178.510 43.120 ;
        RECT 161.510 42.460 165.610 42.520 ;
        RECT 14.810 42.430 18.110 42.460 ;
        RECT 44.310 42.430 47.610 42.460 ;
        RECT 73.810 42.430 77.110 42.460 ;
        RECT 103.310 42.430 106.610 42.460 ;
        RECT 132.810 42.430 136.110 42.460 ;
        RECT 162.310 42.430 165.610 42.460 ;
        RECT 4.865 40.425 5.605 40.485 ;
        RECT 10.350 40.425 23.610 40.430 ;
        RECT 1.510 39.770 23.610 40.425 ;
        RECT 28.480 40.425 29.610 40.640 ;
        RECT 34.365 40.425 35.105 40.485 ;
        RECT 39.850 40.425 53.110 40.430 ;
        RECT 28.480 39.770 53.110 40.425 ;
        RECT 57.980 40.425 59.110 40.640 ;
        RECT 63.865 40.425 64.605 40.485 ;
        RECT 69.350 40.425 82.610 40.430 ;
        RECT 57.980 39.770 82.610 40.425 ;
        RECT 87.480 40.425 88.610 40.640 ;
        RECT 93.365 40.425 94.105 40.485 ;
        RECT 98.850 40.425 112.110 40.430 ;
        RECT 87.480 39.770 112.110 40.425 ;
        RECT 116.980 40.425 118.110 40.640 ;
        RECT 122.865 40.425 123.605 40.485 ;
        RECT 128.350 40.425 141.610 40.430 ;
        RECT 116.980 39.770 141.610 40.425 ;
        RECT 146.480 40.425 147.610 40.640 ;
        RECT 152.365 40.425 153.105 40.485 ;
        RECT 157.850 40.425 171.110 40.430 ;
        RECT 146.480 39.770 171.110 40.425 ;
        RECT 175.980 40.425 177.110 40.640 ;
        RECT 175.980 40.395 178.510 40.425 ;
        RECT 172.150 39.795 178.510 40.395 ;
        RECT 1.510 39.765 13.840 39.770 ;
        RECT 28.480 39.765 43.340 39.770 ;
        RECT 57.980 39.765 72.840 39.770 ;
        RECT 87.480 39.765 102.340 39.770 ;
        RECT 116.980 39.765 131.840 39.770 ;
        RECT 146.480 39.765 161.340 39.770 ;
        RECT 175.980 39.765 178.510 39.795 ;
        RECT 4.865 39.705 5.605 39.765 ;
        RECT 28.480 39.540 29.610 39.765 ;
        RECT 34.365 39.705 35.105 39.765 ;
        RECT 57.980 39.540 59.110 39.765 ;
        RECT 63.865 39.705 64.605 39.765 ;
        RECT 87.480 39.540 88.610 39.765 ;
        RECT 93.365 39.705 94.105 39.765 ;
        RECT 116.980 39.540 118.110 39.765 ;
        RECT 122.865 39.705 123.605 39.765 ;
        RECT 146.480 39.540 147.610 39.765 ;
        RECT 152.365 39.705 153.105 39.765 ;
        RECT 175.980 39.540 177.110 39.765 ;
        RECT 0.000 35.780 178.950 36.260 ;
        RECT 1.510 33.060 179.950 33.540 ;
        RECT 36.000 31.060 38.000 31.500 ;
        RECT 36.000 31.000 37.640 31.060 ;
        RECT 72.000 31.000 74.000 31.500 ;
        RECT 108.000 31.000 110.000 31.500 ;
        RECT 144.000 31.000 146.000 31.500 ;
      LAYER via ;
        RECT 36.130 73.100 36.430 73.400 ;
        RECT 36.490 73.100 36.790 73.400 ;
        RECT 36.850 73.100 37.150 73.400 ;
        RECT 37.210 73.100 37.510 73.400 ;
        RECT 37.570 73.100 37.870 73.400 ;
        RECT 72.130 73.100 72.430 73.400 ;
        RECT 72.490 73.100 72.790 73.400 ;
        RECT 72.850 73.100 73.150 73.400 ;
        RECT 73.210 73.100 73.510 73.400 ;
        RECT 73.570 73.100 73.870 73.400 ;
        RECT 108.130 73.100 108.430 73.400 ;
        RECT 108.490 73.100 108.790 73.400 ;
        RECT 108.850 73.100 109.150 73.400 ;
        RECT 109.210 73.100 109.510 73.400 ;
        RECT 109.570 73.100 109.870 73.400 ;
        RECT 144.130 73.100 144.430 73.400 ;
        RECT 144.490 73.100 144.790 73.400 ;
        RECT 144.850 73.100 145.150 73.400 ;
        RECT 145.210 73.100 145.510 73.400 ;
        RECT 145.570 73.100 145.870 73.400 ;
        RECT 38.510 71.240 38.770 71.500 ;
        RECT 38.880 71.240 39.140 71.500 ;
        RECT 39.250 71.240 39.510 71.500 ;
        RECT 69.510 71.240 69.770 71.500 ;
        RECT 69.880 71.240 70.140 71.500 ;
        RECT 70.250 71.240 70.510 71.500 ;
        RECT 111.510 71.240 111.770 71.500 ;
        RECT 111.880 71.240 112.140 71.500 ;
        RECT 112.250 71.240 112.510 71.500 ;
        RECT 142.510 71.240 142.770 71.500 ;
        RECT 142.880 71.240 143.140 71.500 ;
        RECT 143.250 71.240 143.510 71.500 ;
        RECT 172.000 71.250 172.260 71.510 ;
        RECT 172.320 71.250 172.580 71.510 ;
        RECT 172.640 71.250 172.900 71.510 ;
        RECT 18.130 68.510 18.430 68.810 ;
        RECT 18.490 68.510 18.790 68.810 ;
        RECT 18.850 68.510 19.150 68.810 ;
        RECT 19.210 68.510 19.510 68.810 ;
        RECT 19.570 68.510 19.870 68.810 ;
        RECT 54.130 68.510 54.430 68.810 ;
        RECT 54.490 68.510 54.790 68.810 ;
        RECT 54.850 68.510 55.150 68.810 ;
        RECT 55.210 68.510 55.510 68.810 ;
        RECT 55.570 68.510 55.870 68.810 ;
        RECT 90.130 68.510 90.430 68.810 ;
        RECT 90.490 68.510 90.790 68.810 ;
        RECT 90.850 68.510 91.150 68.810 ;
        RECT 91.210 68.510 91.510 68.810 ;
        RECT 91.570 68.510 91.870 68.810 ;
        RECT 126.130 68.510 126.430 68.810 ;
        RECT 126.490 68.510 126.790 68.810 ;
        RECT 126.850 68.510 127.150 68.810 ;
        RECT 127.210 68.510 127.510 68.810 ;
        RECT 127.570 68.510 127.870 68.810 ;
        RECT 162.130 68.510 162.430 68.810 ;
        RECT 162.490 68.510 162.790 68.810 ;
        RECT 162.850 68.510 163.150 68.810 ;
        RECT 163.210 68.510 163.510 68.810 ;
        RECT 163.570 68.510 163.870 68.810 ;
        RECT 17.555 64.295 18.135 64.875 ;
        RECT 163.990 64.295 164.890 64.875 ;
        RECT 18.130 63.070 18.430 63.370 ;
        RECT 18.490 63.070 18.790 63.370 ;
        RECT 18.850 63.070 19.150 63.370 ;
        RECT 19.210 63.070 19.510 63.370 ;
        RECT 19.570 63.070 19.870 63.370 ;
        RECT 2.400 61.820 2.660 62.080 ;
        RECT 17.435 61.570 18.335 62.150 ;
        RECT 46.290 61.700 46.610 62.020 ;
        RECT 46.770 61.710 47.090 62.030 ;
        RECT 75.730 61.700 76.050 62.020 ;
        RECT 76.210 61.710 76.530 62.030 ;
        RECT 105.170 61.700 105.490 62.020 ;
        RECT 105.650 61.710 105.970 62.030 ;
        RECT 134.610 61.700 134.930 62.020 ;
        RECT 135.090 61.710 135.410 62.030 ;
        RECT 163.980 61.570 164.880 62.150 ;
        RECT 0.130 60.350 0.430 60.650 ;
        RECT 0.490 60.350 0.790 60.650 ;
        RECT 0.850 60.350 1.150 60.650 ;
        RECT 1.210 60.350 1.510 60.650 ;
        RECT 1.570 60.350 1.870 60.650 ;
        RECT 180.130 60.350 180.430 60.650 ;
        RECT 180.490 60.350 180.790 60.650 ;
        RECT 180.850 60.350 181.150 60.650 ;
        RECT 181.210 60.350 181.510 60.650 ;
        RECT 181.570 60.350 181.870 60.650 ;
        RECT 175.130 58.980 175.390 59.240 ;
        RECT 175.450 58.980 175.710 59.240 ;
        RECT 175.770 58.980 176.030 59.240 ;
        RECT 176.090 58.980 176.350 59.240 ;
        RECT 176.410 58.980 176.670 59.240 ;
        RECT 176.730 58.980 176.990 59.240 ;
        RECT 18.130 57.630 18.430 57.930 ;
        RECT 18.490 57.630 18.790 57.930 ;
        RECT 18.850 57.630 19.150 57.930 ;
        RECT 19.210 57.630 19.510 57.930 ;
        RECT 19.570 57.630 19.870 57.930 ;
        RECT 54.130 57.630 54.430 57.930 ;
        RECT 54.490 57.630 54.790 57.930 ;
        RECT 54.850 57.630 55.150 57.930 ;
        RECT 55.210 57.630 55.510 57.930 ;
        RECT 55.570 57.630 55.870 57.930 ;
        RECT 90.130 57.630 90.430 57.930 ;
        RECT 90.490 57.630 90.790 57.930 ;
        RECT 90.850 57.630 91.150 57.930 ;
        RECT 91.210 57.630 91.510 57.930 ;
        RECT 91.570 57.630 91.870 57.930 ;
        RECT 126.130 57.630 126.430 57.930 ;
        RECT 126.490 57.630 126.790 57.930 ;
        RECT 126.850 57.630 127.150 57.930 ;
        RECT 127.210 57.630 127.510 57.930 ;
        RECT 127.570 57.630 127.870 57.930 ;
        RECT 162.130 57.625 162.430 57.925 ;
        RECT 162.490 57.625 162.790 57.925 ;
        RECT 162.850 57.625 163.150 57.925 ;
        RECT 163.210 57.625 163.510 57.925 ;
        RECT 163.570 57.625 163.870 57.925 ;
        RECT 38.510 54.920 38.770 55.180 ;
        RECT 38.880 54.920 39.140 55.180 ;
        RECT 39.250 54.920 39.510 55.180 ;
        RECT 69.510 54.920 69.770 55.180 ;
        RECT 69.880 54.920 70.140 55.180 ;
        RECT 70.250 54.920 70.510 55.180 ;
        RECT 111.510 54.920 111.770 55.180 ;
        RECT 111.880 54.920 112.140 55.180 ;
        RECT 112.250 54.920 112.510 55.180 ;
        RECT 142.510 54.920 142.770 55.180 ;
        RECT 142.880 54.920 143.140 55.180 ;
        RECT 143.250 54.920 143.510 55.180 ;
        RECT 171.980 54.950 172.240 55.210 ;
        RECT 172.340 54.950 172.600 55.210 ;
        RECT 172.700 54.950 172.960 55.210 ;
        RECT 173.060 54.950 173.320 55.210 ;
        RECT 173.430 54.950 173.690 55.210 ;
        RECT 173.790 54.950 174.050 55.210 ;
        RECT 174.170 54.950 174.430 55.210 ;
        RECT 174.545 54.950 174.805 55.210 ;
        RECT 174.925 54.950 175.185 55.210 ;
        RECT 175.300 54.950 175.560 55.210 ;
        RECT 175.675 54.950 175.935 55.210 ;
        RECT 176.045 54.950 176.305 55.210 ;
        RECT 176.425 54.950 176.685 55.210 ;
        RECT 38.510 49.480 38.770 49.740 ;
        RECT 38.880 49.480 39.140 49.740 ;
        RECT 39.250 49.480 39.510 49.740 ;
        RECT 69.510 49.480 69.770 49.740 ;
        RECT 69.880 49.480 70.140 49.740 ;
        RECT 70.250 49.480 70.510 49.740 ;
        RECT 111.510 49.480 111.770 49.740 ;
        RECT 111.880 49.480 112.140 49.740 ;
        RECT 112.250 49.480 112.510 49.740 ;
        RECT 142.510 49.480 142.770 49.740 ;
        RECT 142.880 49.480 143.140 49.740 ;
        RECT 143.250 49.480 143.510 49.740 ;
        RECT 178.975 49.490 179.235 49.750 ;
        RECT 179.295 49.490 179.555 49.750 ;
        RECT 179.615 49.490 179.875 49.750 ;
        RECT 18.130 46.750 18.430 47.050 ;
        RECT 18.490 46.750 18.790 47.050 ;
        RECT 18.850 46.750 19.150 47.050 ;
        RECT 19.210 46.750 19.510 47.050 ;
        RECT 19.570 46.750 19.870 47.050 ;
        RECT 54.130 46.750 54.430 47.050 ;
        RECT 54.490 46.750 54.790 47.050 ;
        RECT 54.850 46.750 55.150 47.050 ;
        RECT 55.210 46.750 55.510 47.050 ;
        RECT 55.570 46.750 55.870 47.050 ;
        RECT 90.130 46.750 90.430 47.050 ;
        RECT 90.490 46.750 90.790 47.050 ;
        RECT 90.850 46.750 91.150 47.050 ;
        RECT 91.210 46.750 91.510 47.050 ;
        RECT 91.570 46.750 91.870 47.050 ;
        RECT 126.130 46.750 126.430 47.050 ;
        RECT 126.490 46.750 126.790 47.050 ;
        RECT 126.850 46.750 127.150 47.050 ;
        RECT 127.210 46.750 127.510 47.050 ;
        RECT 127.570 46.750 127.870 47.050 ;
        RECT 162.130 46.750 162.430 47.050 ;
        RECT 162.490 46.750 162.790 47.050 ;
        RECT 162.850 46.750 163.150 47.050 ;
        RECT 163.210 46.750 163.510 47.050 ;
        RECT 163.570 46.750 163.870 47.050 ;
        RECT 6.275 42.530 6.855 43.110 ;
        RECT 30.650 42.620 30.970 42.940 ;
        RECT 31.130 42.630 31.450 42.950 ;
        RECT 60.090 42.620 60.410 42.940 ;
        RECT 60.570 42.630 60.890 42.950 ;
        RECT 89.530 42.620 89.850 42.940 ;
        RECT 90.010 42.630 90.330 42.950 ;
        RECT 119.430 42.620 119.750 42.940 ;
        RECT 119.910 42.630 120.230 42.950 ;
        RECT 148.870 42.620 149.190 42.940 ;
        RECT 149.350 42.630 149.670 42.950 ;
        RECT 165.660 42.530 166.240 43.110 ;
        RECT 166.380 42.530 166.960 43.110 ;
        RECT 3.565 39.805 4.145 40.385 ;
        RECT 172.270 39.805 172.850 40.385 ;
        RECT 18.130 35.870 18.430 36.170 ;
        RECT 18.490 35.870 18.790 36.170 ;
        RECT 18.850 35.870 19.150 36.170 ;
        RECT 19.210 35.870 19.510 36.170 ;
        RECT 19.570 35.870 19.870 36.170 ;
        RECT 54.130 35.870 54.430 36.170 ;
        RECT 54.490 35.870 54.790 36.170 ;
        RECT 54.850 35.870 55.150 36.170 ;
        RECT 55.210 35.870 55.510 36.170 ;
        RECT 55.570 35.870 55.870 36.170 ;
        RECT 126.130 35.870 126.430 36.170 ;
        RECT 126.490 35.870 126.790 36.170 ;
        RECT 126.850 35.870 127.150 36.170 ;
        RECT 127.210 35.870 127.510 36.170 ;
        RECT 127.570 35.870 127.870 36.170 ;
        RECT 162.130 35.870 162.430 36.170 ;
        RECT 162.490 35.870 162.790 36.170 ;
        RECT 162.850 35.870 163.150 36.170 ;
        RECT 163.210 35.870 163.510 36.170 ;
        RECT 163.570 35.870 163.870 36.170 ;
        RECT 38.510 33.160 38.770 33.420 ;
        RECT 38.880 33.160 39.140 33.420 ;
        RECT 39.250 33.160 39.510 33.420 ;
        RECT 69.510 33.160 69.770 33.420 ;
        RECT 69.880 33.160 70.140 33.420 ;
        RECT 70.250 33.160 70.510 33.420 ;
        RECT 111.510 33.160 111.770 33.420 ;
        RECT 111.880 33.160 112.140 33.420 ;
        RECT 112.250 33.160 112.510 33.420 ;
        RECT 142.510 33.160 142.770 33.420 ;
        RECT 142.880 33.160 143.140 33.420 ;
        RECT 143.250 33.160 143.510 33.420 ;
        RECT 178.985 33.170 179.245 33.430 ;
        RECT 179.305 33.170 179.565 33.430 ;
        RECT 179.625 33.170 179.885 33.430 ;
        RECT 36.130 31.100 36.430 31.400 ;
        RECT 36.490 31.100 36.790 31.400 ;
        RECT 36.850 31.100 37.150 31.400 ;
        RECT 37.210 31.100 37.510 31.400 ;
        RECT 37.570 31.100 37.870 31.400 ;
        RECT 72.130 31.100 72.430 31.400 ;
        RECT 72.490 31.100 72.790 31.400 ;
        RECT 72.850 31.100 73.150 31.400 ;
        RECT 73.210 31.100 73.510 31.400 ;
        RECT 73.570 31.100 73.870 31.400 ;
        RECT 108.130 31.100 108.430 31.400 ;
        RECT 108.490 31.100 108.790 31.400 ;
        RECT 108.850 31.100 109.150 31.400 ;
        RECT 109.210 31.100 109.510 31.400 ;
        RECT 109.570 31.100 109.870 31.400 ;
        RECT 144.130 31.100 144.430 31.400 ;
        RECT 144.490 31.100 144.790 31.400 ;
        RECT 144.850 31.100 145.150 31.400 ;
        RECT 145.210 31.100 145.510 31.400 ;
        RECT 145.570 31.100 145.870 31.400 ;
      LAYER met2 ;
        RECT 36.000 73.000 38.000 73.500 ;
        RECT 72.000 73.000 74.000 73.500 ;
        RECT 108.000 73.000 110.000 73.500 ;
        RECT 144.000 73.000 146.000 73.500 ;
        RECT 38.510 71.170 39.510 71.570 ;
        RECT 69.510 71.170 70.510 71.570 ;
        RECT 111.510 71.170 112.510 71.570 ;
        RECT 142.510 71.170 143.510 71.570 ;
        RECT 18.000 68.420 20.000 68.900 ;
        RECT 54.000 68.420 56.000 68.900 ;
        RECT 90.000 68.420 92.000 68.900 ;
        RECT 126.000 68.420 128.000 68.900 ;
        RECT 162.000 68.420 164.000 68.900 ;
        RECT 17.400 64.935 18.295 64.965 ;
        RECT 13.930 64.235 18.295 64.935 ;
        RECT 2.330 61.800 2.730 62.100 ;
        RECT 0.000 60.260 2.000 60.740 ;
        RECT 13.930 53.350 14.630 64.235 ;
        RECT 17.400 64.205 18.295 64.235 ;
        RECT 163.980 64.935 164.900 64.965 ;
        RECT 163.980 64.235 169.000 64.935 ;
        RECT 163.980 64.205 164.900 64.235 ;
        RECT 18.000 62.980 20.000 63.460 ;
        RECT 18.000 57.540 20.000 58.020 ;
        RECT 54.000 57.540 56.000 58.020 ;
        RECT 90.000 57.540 92.000 58.020 ;
        RECT 126.000 57.540 128.000 58.020 ;
        RECT 162.000 57.535 164.000 58.020 ;
        RECT 38.510 54.850 39.510 55.250 ;
        RECT 69.510 54.850 70.510 55.250 ;
        RECT 111.510 54.850 112.510 55.250 ;
        RECT 142.510 54.850 143.510 55.250 ;
        RECT 3.510 52.650 14.630 53.350 ;
        RECT 3.510 51.835 4.210 52.650 ;
        RECT 3.505 46.265 4.210 51.835 ;
        RECT 168.300 50.935 169.000 64.235 ;
        RECT 171.950 55.540 172.950 71.670 ;
        RECT 180.000 60.260 182.000 60.740 ;
        RECT 171.950 54.540 179.950 55.540 ;
        RECT 178.950 54.000 179.945 54.540 ;
        RECT 168.300 50.235 172.910 50.935 ;
        RECT 38.510 49.410 39.510 49.810 ;
        RECT 69.510 49.410 70.510 49.810 ;
        RECT 111.510 49.410 112.510 49.810 ;
        RECT 142.510 49.410 143.510 49.810 ;
        RECT 18.000 46.660 20.000 47.140 ;
        RECT 54.000 46.660 56.000 47.140 ;
        RECT 90.000 46.660 92.000 47.140 ;
        RECT 126.000 46.660 128.000 47.140 ;
        RECT 162.000 46.660 164.000 47.140 ;
        RECT 3.505 39.715 4.205 46.265 ;
        RECT 172.210 39.745 172.910 50.235 ;
        RECT 18.000 35.780 20.000 36.260 ;
        RECT 54.000 35.780 56.000 36.260 ;
        RECT 126.000 35.780 128.000 36.260 ;
        RECT 162.000 35.780 164.000 36.260 ;
        RECT 38.510 33.090 39.510 33.490 ;
        RECT 69.510 33.090 70.510 33.490 ;
        RECT 111.510 33.090 112.510 33.490 ;
        RECT 142.510 33.090 143.510 33.490 ;
        RECT 178.950 33.010 179.950 54.000 ;
        RECT 36.000 31.060 38.000 31.500 ;
        RECT 36.000 31.000 37.640 31.060 ;
        RECT 72.000 31.000 74.000 31.500 ;
        RECT 108.000 31.000 110.000 31.500 ;
        RECT 144.000 31.000 146.000 31.500 ;
      LAYER via2 ;
        RECT 36.180 73.090 36.500 73.410 ;
        RECT 36.620 73.090 36.940 73.410 ;
        RECT 37.060 73.090 37.380 73.410 ;
        RECT 37.500 73.090 37.820 73.410 ;
        RECT 72.180 73.090 72.500 73.410 ;
        RECT 72.620 73.090 72.940 73.410 ;
        RECT 73.060 73.090 73.380 73.410 ;
        RECT 73.500 73.090 73.820 73.410 ;
        RECT 108.180 73.090 108.500 73.410 ;
        RECT 108.620 73.090 108.940 73.410 ;
        RECT 109.060 73.090 109.380 73.410 ;
        RECT 109.500 73.090 109.820 73.410 ;
        RECT 144.180 73.090 144.500 73.410 ;
        RECT 144.620 73.090 144.940 73.410 ;
        RECT 145.060 73.090 145.380 73.410 ;
        RECT 145.500 73.090 145.820 73.410 ;
        RECT 38.610 71.220 38.910 71.520 ;
        RECT 39.110 71.220 39.410 71.520 ;
        RECT 69.610 71.220 69.910 71.520 ;
        RECT 70.110 71.220 70.410 71.520 ;
        RECT 111.610 71.220 111.910 71.520 ;
        RECT 112.110 71.220 112.410 71.520 ;
        RECT 142.610 71.220 142.910 71.520 ;
        RECT 143.110 71.220 143.410 71.520 ;
        RECT 18.180 68.500 18.500 68.820 ;
        RECT 18.620 68.500 18.940 68.820 ;
        RECT 19.060 68.500 19.380 68.820 ;
        RECT 19.500 68.500 19.820 68.820 ;
        RECT 54.180 68.500 54.500 68.820 ;
        RECT 54.620 68.500 54.940 68.820 ;
        RECT 55.060 68.500 55.380 68.820 ;
        RECT 55.500 68.500 55.820 68.820 ;
        RECT 90.180 68.500 90.500 68.820 ;
        RECT 90.620 68.500 90.940 68.820 ;
        RECT 91.060 68.500 91.380 68.820 ;
        RECT 91.500 68.500 91.820 68.820 ;
        RECT 126.180 68.500 126.500 68.820 ;
        RECT 126.620 68.500 126.940 68.820 ;
        RECT 127.060 68.500 127.380 68.820 ;
        RECT 127.500 68.500 127.820 68.820 ;
        RECT 162.180 68.500 162.500 68.820 ;
        RECT 162.620 68.500 162.940 68.820 ;
        RECT 163.060 68.500 163.380 68.820 ;
        RECT 163.500 68.500 163.820 68.820 ;
        RECT 2.380 61.800 2.680 62.100 ;
        RECT 0.180 60.340 0.500 60.660 ;
        RECT 0.620 60.340 0.940 60.660 ;
        RECT 1.060 60.340 1.380 60.660 ;
        RECT 1.500 60.340 1.820 60.660 ;
        RECT 18.180 63.060 18.500 63.380 ;
        RECT 18.620 63.060 18.940 63.380 ;
        RECT 19.060 63.060 19.380 63.380 ;
        RECT 19.500 63.060 19.820 63.380 ;
        RECT 18.180 57.620 18.500 57.940 ;
        RECT 18.620 57.620 18.940 57.940 ;
        RECT 19.060 57.620 19.380 57.940 ;
        RECT 19.500 57.620 19.820 57.940 ;
        RECT 54.180 57.620 54.500 57.940 ;
        RECT 54.620 57.620 54.940 57.940 ;
        RECT 55.060 57.620 55.380 57.940 ;
        RECT 55.500 57.620 55.820 57.940 ;
        RECT 90.180 57.620 90.500 57.940 ;
        RECT 90.620 57.620 90.940 57.940 ;
        RECT 91.060 57.620 91.380 57.940 ;
        RECT 91.500 57.620 91.820 57.940 ;
        RECT 126.180 57.620 126.500 57.940 ;
        RECT 126.620 57.620 126.940 57.940 ;
        RECT 127.060 57.620 127.380 57.940 ;
        RECT 127.500 57.620 127.820 57.940 ;
        RECT 162.180 57.615 162.500 57.935 ;
        RECT 162.620 57.615 162.940 57.935 ;
        RECT 163.060 57.615 163.380 57.935 ;
        RECT 163.500 57.615 163.820 57.935 ;
        RECT 38.610 54.900 38.910 55.200 ;
        RECT 39.110 54.900 39.410 55.200 ;
        RECT 69.610 54.900 69.910 55.200 ;
        RECT 70.110 54.900 70.410 55.200 ;
        RECT 111.610 54.900 111.910 55.200 ;
        RECT 112.110 54.900 112.410 55.200 ;
        RECT 142.610 54.900 142.910 55.200 ;
        RECT 143.110 54.900 143.410 55.200 ;
        RECT 180.180 60.340 180.500 60.660 ;
        RECT 180.620 60.340 180.940 60.660 ;
        RECT 181.060 60.340 181.380 60.660 ;
        RECT 181.500 60.340 181.820 60.660 ;
        RECT 179.260 52.400 179.660 52.800 ;
        RECT 179.260 51.870 179.660 52.270 ;
        RECT 38.610 49.460 38.910 49.760 ;
        RECT 39.110 49.460 39.410 49.760 ;
        RECT 69.610 49.460 69.910 49.760 ;
        RECT 70.110 49.460 70.410 49.760 ;
        RECT 111.610 49.460 111.910 49.760 ;
        RECT 112.110 49.460 112.410 49.760 ;
        RECT 142.610 49.460 142.910 49.760 ;
        RECT 143.110 49.460 143.410 49.760 ;
        RECT 18.180 46.740 18.500 47.060 ;
        RECT 18.620 46.740 18.940 47.060 ;
        RECT 19.060 46.740 19.380 47.060 ;
        RECT 19.500 46.740 19.820 47.060 ;
        RECT 54.180 46.740 54.500 47.060 ;
        RECT 54.620 46.740 54.940 47.060 ;
        RECT 55.060 46.740 55.380 47.060 ;
        RECT 55.500 46.740 55.820 47.060 ;
        RECT 90.180 46.740 90.500 47.060 ;
        RECT 90.620 46.740 90.940 47.060 ;
        RECT 91.060 46.740 91.380 47.060 ;
        RECT 91.500 46.740 91.820 47.060 ;
        RECT 126.180 46.740 126.500 47.060 ;
        RECT 126.620 46.740 126.940 47.060 ;
        RECT 127.060 46.740 127.380 47.060 ;
        RECT 127.500 46.740 127.820 47.060 ;
        RECT 162.180 46.740 162.500 47.060 ;
        RECT 162.620 46.740 162.940 47.060 ;
        RECT 163.060 46.740 163.380 47.060 ;
        RECT 163.500 46.740 163.820 47.060 ;
        RECT 18.180 35.860 18.500 36.180 ;
        RECT 18.620 35.860 18.940 36.180 ;
        RECT 19.060 35.860 19.380 36.180 ;
        RECT 19.500 35.860 19.820 36.180 ;
        RECT 54.180 35.860 54.500 36.180 ;
        RECT 54.620 35.860 54.940 36.180 ;
        RECT 55.060 35.860 55.380 36.180 ;
        RECT 55.500 35.860 55.820 36.180 ;
        RECT 126.180 35.860 126.500 36.180 ;
        RECT 126.620 35.860 126.940 36.180 ;
        RECT 127.060 35.860 127.380 36.180 ;
        RECT 127.500 35.860 127.820 36.180 ;
        RECT 162.180 35.860 162.500 36.180 ;
        RECT 162.620 35.860 162.940 36.180 ;
        RECT 163.060 35.860 163.380 36.180 ;
        RECT 163.500 35.860 163.820 36.180 ;
        RECT 38.610 33.140 38.910 33.440 ;
        RECT 39.110 33.140 39.410 33.440 ;
        RECT 69.610 33.140 69.910 33.440 ;
        RECT 70.110 33.140 70.410 33.440 ;
        RECT 111.610 33.140 111.910 33.440 ;
        RECT 112.110 33.140 112.410 33.440 ;
        RECT 142.610 33.140 142.910 33.440 ;
        RECT 143.110 33.140 143.410 33.440 ;
        RECT 36.180 31.090 36.500 31.410 ;
        RECT 36.620 31.090 36.940 31.410 ;
        RECT 37.060 31.090 37.380 31.410 ;
        RECT 37.500 31.090 37.820 31.410 ;
        RECT 72.180 31.090 72.500 31.410 ;
        RECT 72.620 31.090 72.940 31.410 ;
        RECT 73.060 31.090 73.380 31.410 ;
        RECT 73.500 31.090 73.820 31.410 ;
        RECT 108.180 31.090 108.500 31.410 ;
        RECT 108.620 31.090 108.940 31.410 ;
        RECT 109.060 31.090 109.380 31.410 ;
        RECT 109.500 31.090 109.820 31.410 ;
        RECT 144.180 31.090 144.500 31.410 ;
        RECT 144.620 31.090 144.940 31.410 ;
        RECT 145.060 31.090 145.380 31.410 ;
        RECT 145.500 31.090 145.820 31.410 ;
      LAYER met3 ;
        RECT 5.000 103.000 177.000 105.000 ;
        RECT 0.000 99.000 182.000 101.000 ;
        RECT 36.000 73.000 38.000 73.500 ;
        RECT 72.000 73.000 74.000 73.500 ;
        RECT 108.000 73.000 110.000 73.500 ;
        RECT 144.000 73.000 146.000 73.500 ;
        RECT 18.000 68.420 20.000 68.900 ;
        RECT 18.000 62.980 20.000 63.460 ;
        RECT 0.000 60.260 2.000 60.740 ;
        RECT 18.000 57.540 20.000 58.020 ;
        RECT 38.510 52.910 39.510 71.620 ;
        RECT 54.000 68.420 56.000 68.900 ;
        RECT 54.000 57.540 56.000 58.020 ;
        RECT 69.510 52.910 70.510 71.620 ;
        RECT 90.000 68.420 92.000 68.900 ;
        RECT 90.000 57.540 92.000 58.020 ;
        RECT 111.510 52.910 112.510 71.620 ;
        RECT 126.000 68.420 128.000 68.900 ;
        RECT 126.000 57.540 128.000 58.020 ;
        RECT 142.510 52.910 143.510 71.620 ;
        RECT 162.000 68.420 164.000 68.900 ;
        RECT 180.000 60.260 182.000 60.740 ;
        RECT 162.000 57.535 164.000 58.020 ;
        RECT 38.510 51.760 179.950 52.910 ;
        RECT 18.000 46.660 20.000 47.140 ;
        RECT 18.000 35.780 20.000 36.260 ;
        RECT 38.510 33.060 39.510 51.760 ;
        RECT 54.000 46.660 56.000 47.140 ;
        RECT 54.000 35.780 56.000 36.260 ;
        RECT 69.510 33.060 70.510 51.760 ;
        RECT 90.000 46.660 92.000 47.140 ;
        RECT 111.510 33.060 112.510 51.760 ;
        RECT 126.000 46.660 128.000 47.140 ;
        RECT 126.000 35.780 128.000 36.260 ;
        RECT 142.510 33.060 143.510 51.760 ;
        RECT 162.000 46.660 164.000 47.140 ;
        RECT 162.000 35.780 164.000 36.260 ;
        RECT 36.000 31.060 38.000 31.500 ;
        RECT 36.000 31.000 37.640 31.060 ;
        RECT 72.000 31.000 74.000 31.500 ;
        RECT 108.000 31.000 110.000 31.500 ;
        RECT 144.000 31.000 146.000 31.500 ;
        RECT 0.000 4.000 182.000 6.000 ;
        RECT 5.000 0.000 177.000 2.000 ;
      LAYER via3 ;
        RECT 5.200 104.400 5.600 104.800 ;
        RECT 5.800 104.400 6.200 104.800 ;
        RECT 6.400 104.400 6.800 104.800 ;
        RECT 18.200 104.400 18.600 104.800 ;
        RECT 18.800 104.400 19.200 104.800 ;
        RECT 19.400 104.400 19.800 104.800 ;
        RECT 54.200 104.400 54.600 104.800 ;
        RECT 54.800 104.400 55.200 104.800 ;
        RECT 55.400 104.400 55.800 104.800 ;
        RECT 90.200 104.400 90.600 104.800 ;
        RECT 90.800 104.400 91.200 104.800 ;
        RECT 91.400 104.400 91.800 104.800 ;
        RECT 126.200 104.400 126.600 104.800 ;
        RECT 126.800 104.400 127.200 104.800 ;
        RECT 127.400 104.400 127.800 104.800 ;
        RECT 162.200 104.400 162.600 104.800 ;
        RECT 162.800 104.400 163.200 104.800 ;
        RECT 163.400 104.400 163.800 104.800 ;
        RECT 175.200 104.400 175.600 104.800 ;
        RECT 175.800 104.400 176.200 104.800 ;
        RECT 176.400 104.400 176.800 104.800 ;
        RECT 5.200 103.800 5.600 104.200 ;
        RECT 5.800 103.800 6.200 104.200 ;
        RECT 6.400 103.800 6.800 104.200 ;
        RECT 18.200 103.800 18.600 104.200 ;
        RECT 18.800 103.800 19.200 104.200 ;
        RECT 19.400 103.800 19.800 104.200 ;
        RECT 54.200 103.800 54.600 104.200 ;
        RECT 54.800 103.800 55.200 104.200 ;
        RECT 55.400 103.800 55.800 104.200 ;
        RECT 90.200 103.800 90.600 104.200 ;
        RECT 90.800 103.800 91.200 104.200 ;
        RECT 91.400 103.800 91.800 104.200 ;
        RECT 126.200 103.800 126.600 104.200 ;
        RECT 126.800 103.800 127.200 104.200 ;
        RECT 127.400 103.800 127.800 104.200 ;
        RECT 162.200 103.800 162.600 104.200 ;
        RECT 162.800 103.800 163.200 104.200 ;
        RECT 163.400 103.800 163.800 104.200 ;
        RECT 175.200 103.800 175.600 104.200 ;
        RECT 175.800 103.800 176.200 104.200 ;
        RECT 176.400 103.800 176.800 104.200 ;
        RECT 5.200 103.200 5.600 103.600 ;
        RECT 5.800 103.200 6.200 103.600 ;
        RECT 6.400 103.200 6.800 103.600 ;
        RECT 18.200 103.200 18.600 103.600 ;
        RECT 18.800 103.200 19.200 103.600 ;
        RECT 19.400 103.200 19.800 103.600 ;
        RECT 54.200 103.200 54.600 103.600 ;
        RECT 54.800 103.200 55.200 103.600 ;
        RECT 55.400 103.200 55.800 103.600 ;
        RECT 90.200 103.200 90.600 103.600 ;
        RECT 90.800 103.200 91.200 103.600 ;
        RECT 91.400 103.200 91.800 103.600 ;
        RECT 126.200 103.200 126.600 103.600 ;
        RECT 126.800 103.200 127.200 103.600 ;
        RECT 127.400 103.200 127.800 103.600 ;
        RECT 162.200 103.200 162.600 103.600 ;
        RECT 162.800 103.200 163.200 103.600 ;
        RECT 163.400 103.200 163.800 103.600 ;
        RECT 175.200 103.200 175.600 103.600 ;
        RECT 175.800 103.200 176.200 103.600 ;
        RECT 176.400 103.200 176.800 103.600 ;
        RECT 0.200 100.400 0.600 100.800 ;
        RECT 0.800 100.400 1.200 100.800 ;
        RECT 1.400 100.400 1.800 100.800 ;
        RECT 36.200 100.400 36.600 100.800 ;
        RECT 36.800 100.400 37.200 100.800 ;
        RECT 37.400 100.400 37.800 100.800 ;
        RECT 72.200 100.400 72.600 100.800 ;
        RECT 72.800 100.400 73.200 100.800 ;
        RECT 73.400 100.400 73.800 100.800 ;
        RECT 108.200 100.400 108.600 100.800 ;
        RECT 108.800 100.400 109.200 100.800 ;
        RECT 109.400 100.400 109.800 100.800 ;
        RECT 144.200 100.400 144.600 100.800 ;
        RECT 144.800 100.400 145.200 100.800 ;
        RECT 145.400 100.400 145.800 100.800 ;
        RECT 180.200 100.400 180.600 100.800 ;
        RECT 180.800 100.400 181.200 100.800 ;
        RECT 181.400 100.400 181.800 100.800 ;
        RECT 0.200 99.800 0.600 100.200 ;
        RECT 0.800 99.800 1.200 100.200 ;
        RECT 1.400 99.800 1.800 100.200 ;
        RECT 36.200 99.800 36.600 100.200 ;
        RECT 36.800 99.800 37.200 100.200 ;
        RECT 37.400 99.800 37.800 100.200 ;
        RECT 72.200 99.800 72.600 100.200 ;
        RECT 72.800 99.800 73.200 100.200 ;
        RECT 73.400 99.800 73.800 100.200 ;
        RECT 108.200 99.800 108.600 100.200 ;
        RECT 108.800 99.800 109.200 100.200 ;
        RECT 109.400 99.800 109.800 100.200 ;
        RECT 144.200 99.800 144.600 100.200 ;
        RECT 144.800 99.800 145.200 100.200 ;
        RECT 145.400 99.800 145.800 100.200 ;
        RECT 180.200 99.800 180.600 100.200 ;
        RECT 180.800 99.800 181.200 100.200 ;
        RECT 181.400 99.800 181.800 100.200 ;
        RECT 0.200 99.200 0.600 99.600 ;
        RECT 0.800 99.200 1.200 99.600 ;
        RECT 1.400 99.200 1.800 99.600 ;
        RECT 36.200 99.200 36.600 99.600 ;
        RECT 36.800 99.200 37.200 99.600 ;
        RECT 37.400 99.200 37.800 99.600 ;
        RECT 72.200 99.200 72.600 99.600 ;
        RECT 72.800 99.200 73.200 99.600 ;
        RECT 73.400 99.200 73.800 99.600 ;
        RECT 108.200 99.200 108.600 99.600 ;
        RECT 108.800 99.200 109.200 99.600 ;
        RECT 109.400 99.200 109.800 99.600 ;
        RECT 144.200 99.200 144.600 99.600 ;
        RECT 144.800 99.200 145.200 99.600 ;
        RECT 145.400 99.200 145.800 99.600 ;
        RECT 180.200 99.200 180.600 99.600 ;
        RECT 180.800 99.200 181.200 99.600 ;
        RECT 181.400 99.200 181.800 99.600 ;
        RECT 36.160 73.070 36.520 73.435 ;
        RECT 36.600 73.070 36.960 73.435 ;
        RECT 37.040 73.070 37.400 73.435 ;
        RECT 37.480 73.070 37.840 73.435 ;
        RECT 72.160 73.070 72.520 73.435 ;
        RECT 72.600 73.070 72.960 73.435 ;
        RECT 73.040 73.070 73.400 73.435 ;
        RECT 73.480 73.070 73.840 73.435 ;
        RECT 108.160 73.070 108.520 73.435 ;
        RECT 108.600 73.070 108.960 73.435 ;
        RECT 109.040 73.070 109.400 73.435 ;
        RECT 109.480 73.070 109.840 73.435 ;
        RECT 144.160 73.070 144.520 73.435 ;
        RECT 144.600 73.070 144.960 73.435 ;
        RECT 145.040 73.070 145.400 73.435 ;
        RECT 145.480 73.070 145.840 73.435 ;
        RECT 18.160 68.480 18.520 68.840 ;
        RECT 18.600 68.480 18.960 68.840 ;
        RECT 19.040 68.480 19.400 68.840 ;
        RECT 19.480 68.480 19.840 68.840 ;
        RECT 18.160 63.040 18.520 63.400 ;
        RECT 18.600 63.040 18.960 63.400 ;
        RECT 19.040 63.040 19.400 63.400 ;
        RECT 19.480 63.040 19.840 63.400 ;
        RECT 0.160 60.320 0.520 60.685 ;
        RECT 0.600 60.320 0.960 60.685 ;
        RECT 1.040 60.320 1.400 60.685 ;
        RECT 1.480 60.320 1.840 60.685 ;
        RECT 18.160 57.600 18.520 57.960 ;
        RECT 18.600 57.600 18.960 57.960 ;
        RECT 19.040 57.600 19.400 57.960 ;
        RECT 19.480 57.600 19.840 57.960 ;
        RECT 54.160 68.480 54.520 68.840 ;
        RECT 54.600 68.480 54.960 68.840 ;
        RECT 55.040 68.480 55.400 68.840 ;
        RECT 55.480 68.480 55.840 68.840 ;
        RECT 54.160 57.600 54.520 57.960 ;
        RECT 54.600 57.600 54.960 57.960 ;
        RECT 55.040 57.600 55.400 57.960 ;
        RECT 55.480 57.600 55.840 57.960 ;
        RECT 90.160 68.480 90.520 68.840 ;
        RECT 90.600 68.480 90.960 68.840 ;
        RECT 91.040 68.480 91.400 68.840 ;
        RECT 91.480 68.480 91.840 68.840 ;
        RECT 90.160 57.600 90.520 57.960 ;
        RECT 90.600 57.600 90.960 57.960 ;
        RECT 91.040 57.600 91.400 57.960 ;
        RECT 91.480 57.600 91.840 57.960 ;
        RECT 126.160 68.480 126.520 68.840 ;
        RECT 126.600 68.480 126.960 68.840 ;
        RECT 127.040 68.480 127.400 68.840 ;
        RECT 127.480 68.480 127.840 68.840 ;
        RECT 126.160 57.600 126.520 57.960 ;
        RECT 126.600 57.600 126.960 57.960 ;
        RECT 127.040 57.600 127.400 57.960 ;
        RECT 127.480 57.600 127.840 57.960 ;
        RECT 162.160 68.480 162.520 68.840 ;
        RECT 162.600 68.480 162.960 68.840 ;
        RECT 163.040 68.480 163.400 68.840 ;
        RECT 163.480 68.480 163.840 68.840 ;
        RECT 180.160 60.320 180.520 60.685 ;
        RECT 180.600 60.320 180.960 60.685 ;
        RECT 181.040 60.320 181.400 60.685 ;
        RECT 181.480 60.320 181.840 60.685 ;
        RECT 162.160 57.595 162.520 57.960 ;
        RECT 162.600 57.595 162.960 57.960 ;
        RECT 163.040 57.595 163.400 57.960 ;
        RECT 163.480 57.595 163.840 57.960 ;
        RECT 18.160 46.720 18.520 47.085 ;
        RECT 18.600 46.720 18.960 47.085 ;
        RECT 19.040 46.720 19.400 47.085 ;
        RECT 19.480 46.720 19.840 47.085 ;
        RECT 18.160 35.840 18.520 36.205 ;
        RECT 18.600 35.840 18.960 36.205 ;
        RECT 19.040 35.840 19.400 36.205 ;
        RECT 19.480 35.840 19.840 36.205 ;
        RECT 54.160 46.720 54.520 47.085 ;
        RECT 54.600 46.720 54.960 47.085 ;
        RECT 55.040 46.720 55.400 47.085 ;
        RECT 55.480 46.720 55.840 47.085 ;
        RECT 54.160 35.840 54.520 36.205 ;
        RECT 54.600 35.840 54.960 36.205 ;
        RECT 55.040 35.840 55.400 36.205 ;
        RECT 55.480 35.840 55.840 36.205 ;
        RECT 90.160 46.720 90.520 47.085 ;
        RECT 90.600 46.720 90.960 47.085 ;
        RECT 91.040 46.720 91.400 47.085 ;
        RECT 91.480 46.720 91.840 47.085 ;
        RECT 126.160 46.720 126.520 47.085 ;
        RECT 126.600 46.720 126.960 47.085 ;
        RECT 127.040 46.720 127.400 47.085 ;
        RECT 127.480 46.720 127.840 47.085 ;
        RECT 126.160 35.840 126.520 36.205 ;
        RECT 126.600 35.840 126.960 36.205 ;
        RECT 127.040 35.840 127.400 36.205 ;
        RECT 127.480 35.840 127.840 36.205 ;
        RECT 162.160 46.720 162.520 47.085 ;
        RECT 162.600 46.720 162.960 47.085 ;
        RECT 163.040 46.720 163.400 47.085 ;
        RECT 163.480 46.720 163.840 47.085 ;
        RECT 162.160 35.840 162.520 36.205 ;
        RECT 162.600 35.840 162.960 36.205 ;
        RECT 163.040 35.840 163.400 36.205 ;
        RECT 163.480 35.840 163.840 36.205 ;
        RECT 36.160 31.070 36.520 31.435 ;
        RECT 36.600 31.070 36.960 31.435 ;
        RECT 37.040 31.070 37.400 31.435 ;
        RECT 37.480 31.070 37.840 31.435 ;
        RECT 72.160 31.070 72.520 31.435 ;
        RECT 72.600 31.070 72.960 31.435 ;
        RECT 73.040 31.070 73.400 31.435 ;
        RECT 73.480 31.070 73.840 31.435 ;
        RECT 108.160 31.070 108.520 31.435 ;
        RECT 108.600 31.070 108.960 31.435 ;
        RECT 109.040 31.070 109.400 31.435 ;
        RECT 109.480 31.070 109.840 31.435 ;
        RECT 144.160 31.070 144.520 31.435 ;
        RECT 144.600 31.070 144.960 31.435 ;
        RECT 145.040 31.070 145.400 31.435 ;
        RECT 145.480 31.070 145.840 31.435 ;
        RECT 0.200 5.400 0.600 5.800 ;
        RECT 0.800 5.400 1.200 5.800 ;
        RECT 1.400 5.400 1.800 5.800 ;
        RECT 36.200 5.400 36.600 5.800 ;
        RECT 36.800 5.400 37.200 5.800 ;
        RECT 37.400 5.400 37.800 5.800 ;
        RECT 72.200 5.400 72.600 5.800 ;
        RECT 72.800 5.400 73.200 5.800 ;
        RECT 73.400 5.400 73.800 5.800 ;
        RECT 108.200 5.400 108.600 5.800 ;
        RECT 108.800 5.400 109.200 5.800 ;
        RECT 109.400 5.400 109.800 5.800 ;
        RECT 144.200 5.400 144.600 5.800 ;
        RECT 144.800 5.400 145.200 5.800 ;
        RECT 145.400 5.400 145.800 5.800 ;
        RECT 180.200 5.400 180.600 5.800 ;
        RECT 180.800 5.400 181.200 5.800 ;
        RECT 181.400 5.400 181.800 5.800 ;
        RECT 0.200 4.800 0.600 5.200 ;
        RECT 0.800 4.800 1.200 5.200 ;
        RECT 1.400 4.800 1.800 5.200 ;
        RECT 36.200 4.800 36.600 5.200 ;
        RECT 36.800 4.800 37.200 5.200 ;
        RECT 37.400 4.800 37.800 5.200 ;
        RECT 72.200 4.800 72.600 5.200 ;
        RECT 72.800 4.800 73.200 5.200 ;
        RECT 73.400 4.800 73.800 5.200 ;
        RECT 108.200 4.800 108.600 5.200 ;
        RECT 108.800 4.800 109.200 5.200 ;
        RECT 109.400 4.800 109.800 5.200 ;
        RECT 144.200 4.800 144.600 5.200 ;
        RECT 144.800 4.800 145.200 5.200 ;
        RECT 145.400 4.800 145.800 5.200 ;
        RECT 180.200 4.800 180.600 5.200 ;
        RECT 180.800 4.800 181.200 5.200 ;
        RECT 181.400 4.800 181.800 5.200 ;
        RECT 0.200 4.200 0.600 4.600 ;
        RECT 0.800 4.200 1.200 4.600 ;
        RECT 1.400 4.200 1.800 4.600 ;
        RECT 36.200 4.200 36.600 4.600 ;
        RECT 36.800 4.200 37.200 4.600 ;
        RECT 37.400 4.200 37.800 4.600 ;
        RECT 72.200 4.200 72.600 4.600 ;
        RECT 72.800 4.200 73.200 4.600 ;
        RECT 73.400 4.200 73.800 4.600 ;
        RECT 108.200 4.200 108.600 4.600 ;
        RECT 108.800 4.200 109.200 4.600 ;
        RECT 109.400 4.200 109.800 4.600 ;
        RECT 144.200 4.200 144.600 4.600 ;
        RECT 144.800 4.200 145.200 4.600 ;
        RECT 145.400 4.200 145.800 4.600 ;
        RECT 180.200 4.200 180.600 4.600 ;
        RECT 180.800 4.200 181.200 4.600 ;
        RECT 181.400 4.200 181.800 4.600 ;
        RECT 5.200 1.400 5.600 1.800 ;
        RECT 5.800 1.400 6.200 1.800 ;
        RECT 6.400 1.400 6.800 1.800 ;
        RECT 18.200 1.400 18.600 1.800 ;
        RECT 18.800 1.400 19.200 1.800 ;
        RECT 19.400 1.400 19.800 1.800 ;
        RECT 54.200 1.400 54.600 1.800 ;
        RECT 54.800 1.400 55.200 1.800 ;
        RECT 55.400 1.400 55.800 1.800 ;
        RECT 90.200 1.400 90.600 1.800 ;
        RECT 90.800 1.400 91.200 1.800 ;
        RECT 91.400 1.400 91.800 1.800 ;
        RECT 126.200 1.400 126.600 1.800 ;
        RECT 126.800 1.400 127.200 1.800 ;
        RECT 127.400 1.400 127.800 1.800 ;
        RECT 162.200 1.400 162.600 1.800 ;
        RECT 162.800 1.400 163.200 1.800 ;
        RECT 163.400 1.400 163.800 1.800 ;
        RECT 175.200 1.400 175.600 1.800 ;
        RECT 175.800 1.400 176.200 1.800 ;
        RECT 176.400 1.400 176.800 1.800 ;
        RECT 5.200 0.800 5.600 1.200 ;
        RECT 5.800 0.800 6.200 1.200 ;
        RECT 6.400 0.800 6.800 1.200 ;
        RECT 18.200 0.800 18.600 1.200 ;
        RECT 18.800 0.800 19.200 1.200 ;
        RECT 19.400 0.800 19.800 1.200 ;
        RECT 54.200 0.800 54.600 1.200 ;
        RECT 54.800 0.800 55.200 1.200 ;
        RECT 55.400 0.800 55.800 1.200 ;
        RECT 90.200 0.800 90.600 1.200 ;
        RECT 90.800 0.800 91.200 1.200 ;
        RECT 91.400 0.800 91.800 1.200 ;
        RECT 126.200 0.800 126.600 1.200 ;
        RECT 126.800 0.800 127.200 1.200 ;
        RECT 127.400 0.800 127.800 1.200 ;
        RECT 162.200 0.800 162.600 1.200 ;
        RECT 162.800 0.800 163.200 1.200 ;
        RECT 163.400 0.800 163.800 1.200 ;
        RECT 175.200 0.800 175.600 1.200 ;
        RECT 175.800 0.800 176.200 1.200 ;
        RECT 176.400 0.800 176.800 1.200 ;
        RECT 5.200 0.200 5.600 0.600 ;
        RECT 5.800 0.200 6.200 0.600 ;
        RECT 6.400 0.200 6.800 0.600 ;
        RECT 18.200 0.200 18.600 0.600 ;
        RECT 18.800 0.200 19.200 0.600 ;
        RECT 19.400 0.200 19.800 0.600 ;
        RECT 54.200 0.200 54.600 0.600 ;
        RECT 54.800 0.200 55.200 0.600 ;
        RECT 55.400 0.200 55.800 0.600 ;
        RECT 90.200 0.200 90.600 0.600 ;
        RECT 90.800 0.200 91.200 0.600 ;
        RECT 91.400 0.200 91.800 0.600 ;
        RECT 126.200 0.200 126.600 0.600 ;
        RECT 126.800 0.200 127.200 0.600 ;
        RECT 127.400 0.200 127.800 0.600 ;
        RECT 162.200 0.200 162.600 0.600 ;
        RECT 162.800 0.200 163.200 0.600 ;
        RECT 163.400 0.200 163.800 0.600 ;
        RECT 175.200 0.200 175.600 0.600 ;
        RECT 175.800 0.200 176.200 0.600 ;
        RECT 176.400 0.200 176.800 0.600 ;
  END
END vco_r100
END LIBRARY

