magic
tech sky130A
magscale 1 2
timestamp 1624928531
<< obsli1 >>
rect 1104 1377 179003 117521
<< obsm1 >>
rect 750 1368 179294 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5170 119200 5226 120000
rect 6734 119200 6790 120000
rect 8206 119200 8262 120000
rect 9678 119200 9734 120000
rect 11242 119200 11298 120000
rect 12714 119200 12770 120000
rect 14186 119200 14242 120000
rect 15750 119200 15806 120000
rect 17222 119200 17278 120000
rect 18694 119200 18750 120000
rect 20258 119200 20314 120000
rect 21730 119200 21786 120000
rect 23202 119200 23258 120000
rect 24674 119200 24730 120000
rect 26238 119200 26294 120000
rect 27710 119200 27766 120000
rect 29182 119200 29238 120000
rect 30746 119200 30802 120000
rect 32218 119200 32274 120000
rect 33690 119200 33746 120000
rect 35254 119200 35310 120000
rect 36726 119200 36782 120000
rect 38198 119200 38254 120000
rect 39762 119200 39818 120000
rect 41234 119200 41290 120000
rect 42706 119200 42762 120000
rect 44178 119200 44234 120000
rect 45742 119200 45798 120000
rect 47214 119200 47270 120000
rect 48686 119200 48742 120000
rect 50250 119200 50306 120000
rect 51722 119200 51778 120000
rect 53194 119200 53250 120000
rect 54758 119200 54814 120000
rect 56230 119200 56286 120000
rect 57702 119200 57758 120000
rect 59266 119200 59322 120000
rect 60738 119200 60794 120000
rect 62210 119200 62266 120000
rect 63682 119200 63738 120000
rect 65246 119200 65302 120000
rect 66718 119200 66774 120000
rect 68190 119200 68246 120000
rect 69754 119200 69810 120000
rect 71226 119200 71282 120000
rect 72698 119200 72754 120000
rect 74262 119200 74318 120000
rect 75734 119200 75790 120000
rect 77206 119200 77262 120000
rect 78770 119200 78826 120000
rect 80242 119200 80298 120000
rect 81714 119200 81770 120000
rect 83186 119200 83242 120000
rect 84750 119200 84806 120000
rect 86222 119200 86278 120000
rect 87694 119200 87750 120000
rect 89258 119200 89314 120000
rect 90730 119200 90786 120000
rect 92202 119200 92258 120000
rect 93766 119200 93822 120000
rect 95238 119200 95294 120000
rect 96710 119200 96766 120000
rect 98274 119200 98330 120000
rect 99746 119200 99802 120000
rect 101218 119200 101274 120000
rect 102690 119200 102746 120000
rect 104254 119200 104310 120000
rect 105726 119200 105782 120000
rect 107198 119200 107254 120000
rect 108762 119200 108818 120000
rect 110234 119200 110290 120000
rect 111706 119200 111762 120000
rect 113270 119200 113326 120000
rect 114742 119200 114798 120000
rect 116214 119200 116270 120000
rect 117778 119200 117834 120000
rect 119250 119200 119306 120000
rect 120722 119200 120778 120000
rect 122194 119200 122250 120000
rect 123758 119200 123814 120000
rect 125230 119200 125286 120000
rect 126702 119200 126758 120000
rect 128266 119200 128322 120000
rect 129738 119200 129794 120000
rect 131210 119200 131266 120000
rect 132774 119200 132830 120000
rect 134246 119200 134302 120000
rect 135718 119200 135774 120000
rect 137282 119200 137338 120000
rect 138754 119200 138810 120000
rect 140226 119200 140282 120000
rect 141698 119200 141754 120000
rect 143262 119200 143318 120000
rect 144734 119200 144790 120000
rect 146206 119200 146262 120000
rect 147770 119200 147826 120000
rect 149242 119200 149298 120000
rect 150714 119200 150770 120000
rect 152278 119200 152334 120000
rect 153750 119200 153806 120000
rect 155222 119200 155278 120000
rect 156786 119200 156842 120000
rect 158258 119200 158314 120000
rect 159730 119200 159786 120000
rect 161202 119200 161258 120000
rect 162766 119200 162822 120000
rect 164238 119200 164294 120000
rect 165710 119200 165766 120000
rect 167274 119200 167330 120000
rect 168746 119200 168802 120000
rect 170218 119200 170274 120000
rect 171782 119200 171838 120000
rect 173254 119200 173310 120000
rect 174726 119200 174782 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5814 0 5870 800
rect 7562 0 7618 800
rect 9218 0 9274 800
rect 10874 0 10930 800
rect 12622 0 12678 800
rect 14278 0 14334 800
rect 15934 0 15990 800
rect 17590 0 17646 800
rect 19338 0 19394 800
rect 20994 0 21050 800
rect 22650 0 22706 800
rect 24398 0 24454 800
rect 26054 0 26110 800
rect 27710 0 27766 800
rect 29366 0 29422 800
rect 31114 0 31170 800
rect 32770 0 32826 800
rect 34426 0 34482 800
rect 36174 0 36230 800
rect 37830 0 37886 800
rect 39486 0 39542 800
rect 41142 0 41198 800
rect 42890 0 42946 800
rect 44546 0 44602 800
rect 46202 0 46258 800
rect 47950 0 48006 800
rect 49606 0 49662 800
rect 51262 0 51318 800
rect 52918 0 52974 800
rect 54666 0 54722 800
rect 56322 0 56378 800
rect 57978 0 58034 800
rect 59726 0 59782 800
rect 61382 0 61438 800
rect 63038 0 63094 800
rect 64786 0 64842 800
rect 66442 0 66498 800
rect 68098 0 68154 800
rect 69754 0 69810 800
rect 71502 0 71558 800
rect 73158 0 73214 800
rect 74814 0 74870 800
rect 76562 0 76618 800
rect 78218 0 78274 800
rect 79874 0 79930 800
rect 81530 0 81586 800
rect 83278 0 83334 800
rect 84934 0 84990 800
rect 86590 0 86646 800
rect 88338 0 88394 800
rect 89994 0 90050 800
rect 91650 0 91706 800
rect 93306 0 93362 800
rect 95054 0 95110 800
rect 96710 0 96766 800
rect 98366 0 98422 800
rect 100114 0 100170 800
rect 101770 0 101826 800
rect 103426 0 103482 800
rect 105082 0 105138 800
rect 106830 0 106886 800
rect 108486 0 108542 800
rect 110142 0 110198 800
rect 111890 0 111946 800
rect 113546 0 113602 800
rect 115202 0 115258 800
rect 116858 0 116914 800
rect 118606 0 118662 800
rect 120262 0 120318 800
rect 121918 0 121974 800
rect 123666 0 123722 800
rect 125322 0 125378 800
rect 126978 0 127034 800
rect 128726 0 128782 800
rect 130382 0 130438 800
rect 132038 0 132094 800
rect 133694 0 133750 800
rect 135442 0 135498 800
rect 137098 0 137154 800
rect 138754 0 138810 800
rect 140502 0 140558 800
rect 142158 0 142214 800
rect 143814 0 143870 800
rect 145470 0 145526 800
rect 147218 0 147274 800
rect 148874 0 148930 800
rect 150530 0 150586 800
rect 152278 0 152334 800
rect 153934 0 153990 800
rect 155590 0 155646 800
rect 157246 0 157302 800
rect 158994 0 159050 800
rect 160650 0 160706 800
rect 162306 0 162362 800
rect 164054 0 164110 800
rect 165710 0 165766 800
rect 167366 0 167422 800
rect 169022 0 169078 800
rect 170770 0 170826 800
rect 172426 0 172482 800
rect 174082 0 174138 800
rect 175830 0 175886 800
rect 177486 0 177542 800
rect 179142 0 179198 800
<< obsm2 >>
rect 866 119144 2170 119377
rect 2338 119144 3642 119377
rect 3810 119144 5114 119377
rect 5282 119144 6678 119377
rect 6846 119144 8150 119377
rect 8318 119144 9622 119377
rect 9790 119144 11186 119377
rect 11354 119144 12658 119377
rect 12826 119144 14130 119377
rect 14298 119144 15694 119377
rect 15862 119144 17166 119377
rect 17334 119144 18638 119377
rect 18806 119144 20202 119377
rect 20370 119144 21674 119377
rect 21842 119144 23146 119377
rect 23314 119144 24618 119377
rect 24786 119144 26182 119377
rect 26350 119144 27654 119377
rect 27822 119144 29126 119377
rect 29294 119144 30690 119377
rect 30858 119144 32162 119377
rect 32330 119144 33634 119377
rect 33802 119144 35198 119377
rect 35366 119144 36670 119377
rect 36838 119144 38142 119377
rect 38310 119144 39706 119377
rect 39874 119144 41178 119377
rect 41346 119144 42650 119377
rect 42818 119144 44122 119377
rect 44290 119144 45686 119377
rect 45854 119144 47158 119377
rect 47326 119144 48630 119377
rect 48798 119144 50194 119377
rect 50362 119144 51666 119377
rect 51834 119144 53138 119377
rect 53306 119144 54702 119377
rect 54870 119144 56174 119377
rect 56342 119144 57646 119377
rect 57814 119144 59210 119377
rect 59378 119144 60682 119377
rect 60850 119144 62154 119377
rect 62322 119144 63626 119377
rect 63794 119144 65190 119377
rect 65358 119144 66662 119377
rect 66830 119144 68134 119377
rect 68302 119144 69698 119377
rect 69866 119144 71170 119377
rect 71338 119144 72642 119377
rect 72810 119144 74206 119377
rect 74374 119144 75678 119377
rect 75846 119144 77150 119377
rect 77318 119144 78714 119377
rect 78882 119144 80186 119377
rect 80354 119144 81658 119377
rect 81826 119144 83130 119377
rect 83298 119144 84694 119377
rect 84862 119144 86166 119377
rect 86334 119144 87638 119377
rect 87806 119144 89202 119377
rect 89370 119144 90674 119377
rect 90842 119144 92146 119377
rect 92314 119144 93710 119377
rect 93878 119144 95182 119377
rect 95350 119144 96654 119377
rect 96822 119144 98218 119377
rect 98386 119144 99690 119377
rect 99858 119144 101162 119377
rect 101330 119144 102634 119377
rect 102802 119144 104198 119377
rect 104366 119144 105670 119377
rect 105838 119144 107142 119377
rect 107310 119144 108706 119377
rect 108874 119144 110178 119377
rect 110346 119144 111650 119377
rect 111818 119144 113214 119377
rect 113382 119144 114686 119377
rect 114854 119144 116158 119377
rect 116326 119144 117722 119377
rect 117890 119144 119194 119377
rect 119362 119144 120666 119377
rect 120834 119144 122138 119377
rect 122306 119144 123702 119377
rect 123870 119144 125174 119377
rect 125342 119144 126646 119377
rect 126814 119144 128210 119377
rect 128378 119144 129682 119377
rect 129850 119144 131154 119377
rect 131322 119144 132718 119377
rect 132886 119144 134190 119377
rect 134358 119144 135662 119377
rect 135830 119144 137226 119377
rect 137394 119144 138698 119377
rect 138866 119144 140170 119377
rect 140338 119144 141642 119377
rect 141810 119144 143206 119377
rect 143374 119144 144678 119377
rect 144846 119144 146150 119377
rect 146318 119144 147714 119377
rect 147882 119144 149186 119377
rect 149354 119144 150658 119377
rect 150826 119144 152222 119377
rect 152390 119144 153694 119377
rect 153862 119144 155166 119377
rect 155334 119144 156730 119377
rect 156898 119144 158202 119377
rect 158370 119144 159674 119377
rect 159842 119144 161146 119377
rect 161314 119144 162710 119377
rect 162878 119144 164182 119377
rect 164350 119144 165654 119377
rect 165822 119144 167218 119377
rect 167386 119144 168690 119377
rect 168858 119144 170162 119377
rect 170330 119144 171726 119377
rect 171894 119144 173198 119377
rect 173366 119144 174670 119377
rect 174838 119144 176234 119377
rect 176402 119144 177706 119377
rect 177874 119144 179178 119377
rect 756 856 179288 119144
rect 756 439 790 856
rect 958 439 2446 856
rect 2614 439 4102 856
rect 4270 439 5758 856
rect 5926 439 7506 856
rect 7674 439 9162 856
rect 9330 439 10818 856
rect 10986 439 12566 856
rect 12734 439 14222 856
rect 14390 439 15878 856
rect 16046 439 17534 856
rect 17702 439 19282 856
rect 19450 439 20938 856
rect 21106 439 22594 856
rect 22762 439 24342 856
rect 24510 439 25998 856
rect 26166 439 27654 856
rect 27822 439 29310 856
rect 29478 439 31058 856
rect 31226 439 32714 856
rect 32882 439 34370 856
rect 34538 439 36118 856
rect 36286 439 37774 856
rect 37942 439 39430 856
rect 39598 439 41086 856
rect 41254 439 42834 856
rect 43002 439 44490 856
rect 44658 439 46146 856
rect 46314 439 47894 856
rect 48062 439 49550 856
rect 49718 439 51206 856
rect 51374 439 52862 856
rect 53030 439 54610 856
rect 54778 439 56266 856
rect 56434 439 57922 856
rect 58090 439 59670 856
rect 59838 439 61326 856
rect 61494 439 62982 856
rect 63150 439 64730 856
rect 64898 439 66386 856
rect 66554 439 68042 856
rect 68210 439 69698 856
rect 69866 439 71446 856
rect 71614 439 73102 856
rect 73270 439 74758 856
rect 74926 439 76506 856
rect 76674 439 78162 856
rect 78330 439 79818 856
rect 79986 439 81474 856
rect 81642 439 83222 856
rect 83390 439 84878 856
rect 85046 439 86534 856
rect 86702 439 88282 856
rect 88450 439 89938 856
rect 90106 439 91594 856
rect 91762 439 93250 856
rect 93418 439 94998 856
rect 95166 439 96654 856
rect 96822 439 98310 856
rect 98478 439 100058 856
rect 100226 439 101714 856
rect 101882 439 103370 856
rect 103538 439 105026 856
rect 105194 439 106774 856
rect 106942 439 108430 856
rect 108598 439 110086 856
rect 110254 439 111834 856
rect 112002 439 113490 856
rect 113658 439 115146 856
rect 115314 439 116802 856
rect 116970 439 118550 856
rect 118718 439 120206 856
rect 120374 439 121862 856
rect 122030 439 123610 856
rect 123778 439 125266 856
rect 125434 439 126922 856
rect 127090 439 128670 856
rect 128838 439 130326 856
rect 130494 439 131982 856
rect 132150 439 133638 856
rect 133806 439 135386 856
rect 135554 439 137042 856
rect 137210 439 138698 856
rect 138866 439 140446 856
rect 140614 439 142102 856
rect 142270 439 143758 856
rect 143926 439 145414 856
rect 145582 439 147162 856
rect 147330 439 148818 856
rect 148986 439 150474 856
rect 150642 439 152222 856
rect 152390 439 153878 856
rect 154046 439 155534 856
rect 155702 439 157190 856
rect 157358 439 158938 856
rect 159106 439 160594 856
rect 160762 439 162250 856
rect 162418 439 163998 856
rect 164166 439 165654 856
rect 165822 439 167310 856
rect 167478 439 168966 856
rect 169134 439 170714 856
rect 170882 439 172370 856
rect 172538 439 174026 856
rect 174194 439 175774 856
rect 175942 439 177430 856
rect 177598 439 179086 856
rect 179254 439 179288 856
<< metal3 >>
rect 0 119280 800 119400
rect 179200 119280 180000 119400
rect 0 118328 800 118448
rect 179200 118192 180000 118312
rect 0 117376 800 117496
rect 179200 117104 180000 117224
rect 0 116424 800 116544
rect 179200 116016 180000 116136
rect 0 115336 800 115456
rect 179200 114928 180000 115048
rect 0 114384 800 114504
rect 179200 113840 180000 113960
rect 0 113432 800 113552
rect 179200 112752 180000 112872
rect 0 112480 800 112600
rect 179200 111664 180000 111784
rect 0 111392 800 111512
rect 0 110440 800 110560
rect 179200 110576 180000 110696
rect 0 109488 800 109608
rect 179200 109488 180000 109608
rect 0 108536 800 108656
rect 179200 108400 180000 108520
rect 0 107584 800 107704
rect 179200 107312 180000 107432
rect 0 106496 800 106616
rect 179200 106224 180000 106344
rect 0 105544 800 105664
rect 179200 105136 180000 105256
rect 0 104592 800 104712
rect 179200 104048 180000 104168
rect 0 103640 800 103760
rect 179200 102960 180000 103080
rect 0 102552 800 102672
rect 179200 101872 180000 101992
rect 0 101600 800 101720
rect 0 100648 800 100768
rect 179200 100784 180000 100904
rect 0 99696 800 99816
rect 179200 99832 180000 99952
rect 0 98608 800 98728
rect 179200 98744 180000 98864
rect 0 97656 800 97776
rect 179200 97656 180000 97776
rect 0 96704 800 96824
rect 179200 96568 180000 96688
rect 0 95752 800 95872
rect 179200 95480 180000 95600
rect 0 94800 800 94920
rect 179200 94392 180000 94512
rect 0 93712 800 93832
rect 179200 93304 180000 93424
rect 0 92760 800 92880
rect 179200 92216 180000 92336
rect 0 91808 800 91928
rect 179200 91128 180000 91248
rect 0 90856 800 90976
rect 179200 90040 180000 90160
rect 0 89768 800 89888
rect 0 88816 800 88936
rect 179200 88952 180000 89072
rect 0 87864 800 87984
rect 179200 87864 180000 87984
rect 0 86912 800 87032
rect 179200 86776 180000 86896
rect 0 85824 800 85944
rect 179200 85688 180000 85808
rect 0 84872 800 84992
rect 179200 84600 180000 84720
rect 0 83920 800 84040
rect 179200 83512 180000 83632
rect 0 82968 800 83088
rect 179200 82424 180000 82544
rect 0 82016 800 82136
rect 179200 81336 180000 81456
rect 0 80928 800 81048
rect 179200 80384 180000 80504
rect 0 79976 800 80096
rect 179200 79296 180000 79416
rect 0 79024 800 79144
rect 0 78072 800 78192
rect 179200 78208 180000 78328
rect 0 76984 800 77104
rect 179200 77120 180000 77240
rect 0 76032 800 76152
rect 179200 76032 180000 76152
rect 0 75080 800 75200
rect 179200 74944 180000 75064
rect 0 74128 800 74248
rect 179200 73856 180000 73976
rect 0 73040 800 73160
rect 179200 72768 180000 72888
rect 0 72088 800 72208
rect 179200 71680 180000 71800
rect 0 71136 800 71256
rect 179200 70592 180000 70712
rect 0 70184 800 70304
rect 179200 69504 180000 69624
rect 0 69232 800 69352
rect 179200 68416 180000 68536
rect 0 68144 800 68264
rect 0 67192 800 67312
rect 179200 67328 180000 67448
rect 0 66240 800 66360
rect 179200 66240 180000 66360
rect 0 65288 800 65408
rect 179200 65152 180000 65272
rect 0 64200 800 64320
rect 179200 64064 180000 64184
rect 0 63248 800 63368
rect 179200 62976 180000 63096
rect 0 62296 800 62416
rect 179200 61888 180000 62008
rect 0 61344 800 61464
rect 179200 60800 180000 60920
rect 0 60392 800 60512
rect 179200 59848 180000 59968
rect 0 59304 800 59424
rect 179200 58760 180000 58880
rect 0 58352 800 58472
rect 179200 57672 180000 57792
rect 0 57400 800 57520
rect 0 56448 800 56568
rect 179200 56584 180000 56704
rect 0 55360 800 55480
rect 179200 55496 180000 55616
rect 0 54408 800 54528
rect 179200 54408 180000 54528
rect 0 53456 800 53576
rect 179200 53320 180000 53440
rect 0 52504 800 52624
rect 179200 52232 180000 52352
rect 0 51416 800 51536
rect 179200 51144 180000 51264
rect 0 50464 800 50584
rect 179200 50056 180000 50176
rect 0 49512 800 49632
rect 179200 48968 180000 49088
rect 0 48560 800 48680
rect 179200 47880 180000 48000
rect 0 47608 800 47728
rect 179200 46792 180000 46912
rect 0 46520 800 46640
rect 0 45568 800 45688
rect 179200 45704 180000 45824
rect 0 44616 800 44736
rect 179200 44616 180000 44736
rect 0 43664 800 43784
rect 179200 43528 180000 43648
rect 0 42576 800 42696
rect 179200 42440 180000 42560
rect 0 41624 800 41744
rect 179200 41352 180000 41472
rect 0 40672 800 40792
rect 179200 40400 180000 40520
rect 0 39720 800 39840
rect 179200 39312 180000 39432
rect 0 38632 800 38752
rect 179200 38224 180000 38344
rect 0 37680 800 37800
rect 179200 37136 180000 37256
rect 0 36728 800 36848
rect 179200 36048 180000 36168
rect 0 35776 800 35896
rect 0 34824 800 34944
rect 179200 34960 180000 35080
rect 0 33736 800 33856
rect 179200 33872 180000 33992
rect 0 32784 800 32904
rect 179200 32784 180000 32904
rect 0 31832 800 31952
rect 179200 31696 180000 31816
rect 0 30880 800 31000
rect 179200 30608 180000 30728
rect 0 29792 800 29912
rect 179200 29520 180000 29640
rect 0 28840 800 28960
rect 179200 28432 180000 28552
rect 0 27888 800 28008
rect 179200 27344 180000 27464
rect 0 26936 800 27056
rect 179200 26256 180000 26376
rect 0 25848 800 25968
rect 179200 25168 180000 25288
rect 0 24896 800 25016
rect 0 23944 800 24064
rect 179200 24080 180000 24200
rect 0 22992 800 23112
rect 179200 22992 180000 23112
rect 0 22040 800 22160
rect 179200 21904 180000 22024
rect 0 20952 800 21072
rect 179200 20816 180000 20936
rect 0 20000 800 20120
rect 179200 19864 180000 19984
rect 0 19048 800 19168
rect 179200 18776 180000 18896
rect 0 18096 800 18216
rect 179200 17688 180000 17808
rect 0 17008 800 17128
rect 179200 16600 180000 16720
rect 0 16056 800 16176
rect 179200 15512 180000 15632
rect 0 15104 800 15224
rect 179200 14424 180000 14544
rect 0 14152 800 14272
rect 179200 13336 180000 13456
rect 0 13064 800 13184
rect 0 12112 800 12232
rect 179200 12248 180000 12368
rect 0 11160 800 11280
rect 179200 11160 180000 11280
rect 0 10208 800 10328
rect 179200 10072 180000 10192
rect 0 9256 800 9376
rect 179200 8984 180000 9104
rect 0 8168 800 8288
rect 179200 7896 180000 8016
rect 0 7216 800 7336
rect 179200 6808 180000 6928
rect 0 6264 800 6384
rect 179200 5720 180000 5840
rect 0 5312 800 5432
rect 179200 4632 180000 4752
rect 0 4224 800 4344
rect 179200 3544 180000 3664
rect 0 3272 800 3392
rect 0 2320 800 2440
rect 179200 2456 180000 2576
rect 0 1368 800 1488
rect 179200 1368 180000 1488
rect 0 416 800 536
rect 179200 416 180000 536
<< obsm3 >>
rect 880 119200 179120 119373
rect 800 118528 179200 119200
rect 880 118392 179200 118528
rect 880 118248 179120 118392
rect 800 118112 179120 118248
rect 800 117576 179200 118112
rect 880 117304 179200 117576
rect 880 117296 179120 117304
rect 800 117024 179120 117296
rect 800 116624 179200 117024
rect 880 116344 179200 116624
rect 800 116216 179200 116344
rect 800 115936 179120 116216
rect 800 115536 179200 115936
rect 880 115256 179200 115536
rect 800 115128 179200 115256
rect 800 114848 179120 115128
rect 800 114584 179200 114848
rect 880 114304 179200 114584
rect 800 114040 179200 114304
rect 800 113760 179120 114040
rect 800 113632 179200 113760
rect 880 113352 179200 113632
rect 800 112952 179200 113352
rect 800 112680 179120 112952
rect 880 112672 179120 112680
rect 880 112400 179200 112672
rect 800 111864 179200 112400
rect 800 111592 179120 111864
rect 880 111584 179120 111592
rect 880 111312 179200 111584
rect 800 110776 179200 111312
rect 800 110640 179120 110776
rect 880 110496 179120 110640
rect 880 110360 179200 110496
rect 800 109688 179200 110360
rect 880 109408 179120 109688
rect 800 108736 179200 109408
rect 880 108600 179200 108736
rect 880 108456 179120 108600
rect 800 108320 179120 108456
rect 800 107784 179200 108320
rect 880 107512 179200 107784
rect 880 107504 179120 107512
rect 800 107232 179120 107504
rect 800 106696 179200 107232
rect 880 106424 179200 106696
rect 880 106416 179120 106424
rect 800 106144 179120 106416
rect 800 105744 179200 106144
rect 880 105464 179200 105744
rect 800 105336 179200 105464
rect 800 105056 179120 105336
rect 800 104792 179200 105056
rect 880 104512 179200 104792
rect 800 104248 179200 104512
rect 800 103968 179120 104248
rect 800 103840 179200 103968
rect 880 103560 179200 103840
rect 800 103160 179200 103560
rect 800 102880 179120 103160
rect 800 102752 179200 102880
rect 880 102472 179200 102752
rect 800 102072 179200 102472
rect 800 101800 179120 102072
rect 880 101792 179120 101800
rect 880 101520 179200 101792
rect 800 100984 179200 101520
rect 800 100848 179120 100984
rect 880 100704 179120 100848
rect 880 100568 179200 100704
rect 800 100032 179200 100568
rect 800 99896 179120 100032
rect 880 99752 179120 99896
rect 880 99616 179200 99752
rect 800 98944 179200 99616
rect 800 98808 179120 98944
rect 880 98664 179120 98808
rect 880 98528 179200 98664
rect 800 97856 179200 98528
rect 880 97576 179120 97856
rect 800 96904 179200 97576
rect 880 96768 179200 96904
rect 880 96624 179120 96768
rect 800 96488 179120 96624
rect 800 95952 179200 96488
rect 880 95680 179200 95952
rect 880 95672 179120 95680
rect 800 95400 179120 95672
rect 800 95000 179200 95400
rect 880 94720 179200 95000
rect 800 94592 179200 94720
rect 800 94312 179120 94592
rect 800 93912 179200 94312
rect 880 93632 179200 93912
rect 800 93504 179200 93632
rect 800 93224 179120 93504
rect 800 92960 179200 93224
rect 880 92680 179200 92960
rect 800 92416 179200 92680
rect 800 92136 179120 92416
rect 800 92008 179200 92136
rect 880 91728 179200 92008
rect 800 91328 179200 91728
rect 800 91056 179120 91328
rect 880 91048 179120 91056
rect 880 90776 179200 91048
rect 800 90240 179200 90776
rect 800 89968 179120 90240
rect 880 89960 179120 89968
rect 880 89688 179200 89960
rect 800 89152 179200 89688
rect 800 89016 179120 89152
rect 880 88872 179120 89016
rect 880 88736 179200 88872
rect 800 88064 179200 88736
rect 880 87784 179120 88064
rect 800 87112 179200 87784
rect 880 86976 179200 87112
rect 880 86832 179120 86976
rect 800 86696 179120 86832
rect 800 86024 179200 86696
rect 880 85888 179200 86024
rect 880 85744 179120 85888
rect 800 85608 179120 85744
rect 800 85072 179200 85608
rect 880 84800 179200 85072
rect 880 84792 179120 84800
rect 800 84520 179120 84792
rect 800 84120 179200 84520
rect 880 83840 179200 84120
rect 800 83712 179200 83840
rect 800 83432 179120 83712
rect 800 83168 179200 83432
rect 880 82888 179200 83168
rect 800 82624 179200 82888
rect 800 82344 179120 82624
rect 800 82216 179200 82344
rect 880 81936 179200 82216
rect 800 81536 179200 81936
rect 800 81256 179120 81536
rect 800 81128 179200 81256
rect 880 80848 179200 81128
rect 800 80584 179200 80848
rect 800 80304 179120 80584
rect 800 80176 179200 80304
rect 880 79896 179200 80176
rect 800 79496 179200 79896
rect 800 79224 179120 79496
rect 880 79216 179120 79224
rect 880 78944 179200 79216
rect 800 78408 179200 78944
rect 800 78272 179120 78408
rect 880 78128 179120 78272
rect 880 77992 179200 78128
rect 800 77320 179200 77992
rect 800 77184 179120 77320
rect 880 77040 179120 77184
rect 880 76904 179200 77040
rect 800 76232 179200 76904
rect 880 75952 179120 76232
rect 800 75280 179200 75952
rect 880 75144 179200 75280
rect 880 75000 179120 75144
rect 800 74864 179120 75000
rect 800 74328 179200 74864
rect 880 74056 179200 74328
rect 880 74048 179120 74056
rect 800 73776 179120 74048
rect 800 73240 179200 73776
rect 880 72968 179200 73240
rect 880 72960 179120 72968
rect 800 72688 179120 72960
rect 800 72288 179200 72688
rect 880 72008 179200 72288
rect 800 71880 179200 72008
rect 800 71600 179120 71880
rect 800 71336 179200 71600
rect 880 71056 179200 71336
rect 800 70792 179200 71056
rect 800 70512 179120 70792
rect 800 70384 179200 70512
rect 880 70104 179200 70384
rect 800 69704 179200 70104
rect 800 69432 179120 69704
rect 880 69424 179120 69432
rect 880 69152 179200 69424
rect 800 68616 179200 69152
rect 800 68344 179120 68616
rect 880 68336 179120 68344
rect 880 68064 179200 68336
rect 800 67528 179200 68064
rect 800 67392 179120 67528
rect 880 67248 179120 67392
rect 880 67112 179200 67248
rect 800 66440 179200 67112
rect 880 66160 179120 66440
rect 800 65488 179200 66160
rect 880 65352 179200 65488
rect 880 65208 179120 65352
rect 800 65072 179120 65208
rect 800 64400 179200 65072
rect 880 64264 179200 64400
rect 880 64120 179120 64264
rect 800 63984 179120 64120
rect 800 63448 179200 63984
rect 880 63176 179200 63448
rect 880 63168 179120 63176
rect 800 62896 179120 63168
rect 800 62496 179200 62896
rect 880 62216 179200 62496
rect 800 62088 179200 62216
rect 800 61808 179120 62088
rect 800 61544 179200 61808
rect 880 61264 179200 61544
rect 800 61000 179200 61264
rect 800 60720 179120 61000
rect 800 60592 179200 60720
rect 880 60312 179200 60592
rect 800 60048 179200 60312
rect 800 59768 179120 60048
rect 800 59504 179200 59768
rect 880 59224 179200 59504
rect 800 58960 179200 59224
rect 800 58680 179120 58960
rect 800 58552 179200 58680
rect 880 58272 179200 58552
rect 800 57872 179200 58272
rect 800 57600 179120 57872
rect 880 57592 179120 57600
rect 880 57320 179200 57592
rect 800 56784 179200 57320
rect 800 56648 179120 56784
rect 880 56504 179120 56648
rect 880 56368 179200 56504
rect 800 55696 179200 56368
rect 800 55560 179120 55696
rect 880 55416 179120 55560
rect 880 55280 179200 55416
rect 800 54608 179200 55280
rect 880 54328 179120 54608
rect 800 53656 179200 54328
rect 880 53520 179200 53656
rect 880 53376 179120 53520
rect 800 53240 179120 53376
rect 800 52704 179200 53240
rect 880 52432 179200 52704
rect 880 52424 179120 52432
rect 800 52152 179120 52424
rect 800 51616 179200 52152
rect 880 51344 179200 51616
rect 880 51336 179120 51344
rect 800 51064 179120 51336
rect 800 50664 179200 51064
rect 880 50384 179200 50664
rect 800 50256 179200 50384
rect 800 49976 179120 50256
rect 800 49712 179200 49976
rect 880 49432 179200 49712
rect 800 49168 179200 49432
rect 800 48888 179120 49168
rect 800 48760 179200 48888
rect 880 48480 179200 48760
rect 800 48080 179200 48480
rect 800 47808 179120 48080
rect 880 47800 179120 47808
rect 880 47528 179200 47800
rect 800 46992 179200 47528
rect 800 46720 179120 46992
rect 880 46712 179120 46720
rect 880 46440 179200 46712
rect 800 45904 179200 46440
rect 800 45768 179120 45904
rect 880 45624 179120 45768
rect 880 45488 179200 45624
rect 800 44816 179200 45488
rect 880 44536 179120 44816
rect 800 43864 179200 44536
rect 880 43728 179200 43864
rect 880 43584 179120 43728
rect 800 43448 179120 43584
rect 800 42776 179200 43448
rect 880 42640 179200 42776
rect 880 42496 179120 42640
rect 800 42360 179120 42496
rect 800 41824 179200 42360
rect 880 41552 179200 41824
rect 880 41544 179120 41552
rect 800 41272 179120 41544
rect 800 40872 179200 41272
rect 880 40600 179200 40872
rect 880 40592 179120 40600
rect 800 40320 179120 40592
rect 800 39920 179200 40320
rect 880 39640 179200 39920
rect 800 39512 179200 39640
rect 800 39232 179120 39512
rect 800 38832 179200 39232
rect 880 38552 179200 38832
rect 800 38424 179200 38552
rect 800 38144 179120 38424
rect 800 37880 179200 38144
rect 880 37600 179200 37880
rect 800 37336 179200 37600
rect 800 37056 179120 37336
rect 800 36928 179200 37056
rect 880 36648 179200 36928
rect 800 36248 179200 36648
rect 800 35976 179120 36248
rect 880 35968 179120 35976
rect 880 35696 179200 35968
rect 800 35160 179200 35696
rect 800 35024 179120 35160
rect 880 34880 179120 35024
rect 880 34744 179200 34880
rect 800 34072 179200 34744
rect 800 33936 179120 34072
rect 880 33792 179120 33936
rect 880 33656 179200 33792
rect 800 32984 179200 33656
rect 880 32704 179120 32984
rect 800 32032 179200 32704
rect 880 31896 179200 32032
rect 880 31752 179120 31896
rect 800 31616 179120 31752
rect 800 31080 179200 31616
rect 880 30808 179200 31080
rect 880 30800 179120 30808
rect 800 30528 179120 30800
rect 800 29992 179200 30528
rect 880 29720 179200 29992
rect 880 29712 179120 29720
rect 800 29440 179120 29712
rect 800 29040 179200 29440
rect 880 28760 179200 29040
rect 800 28632 179200 28760
rect 800 28352 179120 28632
rect 800 28088 179200 28352
rect 880 27808 179200 28088
rect 800 27544 179200 27808
rect 800 27264 179120 27544
rect 800 27136 179200 27264
rect 880 26856 179200 27136
rect 800 26456 179200 26856
rect 800 26176 179120 26456
rect 800 26048 179200 26176
rect 880 25768 179200 26048
rect 800 25368 179200 25768
rect 800 25096 179120 25368
rect 880 25088 179120 25096
rect 880 24816 179200 25088
rect 800 24280 179200 24816
rect 800 24144 179120 24280
rect 880 24000 179120 24144
rect 880 23864 179200 24000
rect 800 23192 179200 23864
rect 880 22912 179120 23192
rect 800 22240 179200 22912
rect 880 22104 179200 22240
rect 880 21960 179120 22104
rect 800 21824 179120 21960
rect 800 21152 179200 21824
rect 880 21016 179200 21152
rect 880 20872 179120 21016
rect 800 20736 179120 20872
rect 800 20200 179200 20736
rect 880 20064 179200 20200
rect 880 19920 179120 20064
rect 800 19784 179120 19920
rect 800 19248 179200 19784
rect 880 18976 179200 19248
rect 880 18968 179120 18976
rect 800 18696 179120 18968
rect 800 18296 179200 18696
rect 880 18016 179200 18296
rect 800 17888 179200 18016
rect 800 17608 179120 17888
rect 800 17208 179200 17608
rect 880 16928 179200 17208
rect 800 16800 179200 16928
rect 800 16520 179120 16800
rect 800 16256 179200 16520
rect 880 15976 179200 16256
rect 800 15712 179200 15976
rect 800 15432 179120 15712
rect 800 15304 179200 15432
rect 880 15024 179200 15304
rect 800 14624 179200 15024
rect 800 14352 179120 14624
rect 880 14344 179120 14352
rect 880 14072 179200 14344
rect 800 13536 179200 14072
rect 800 13264 179120 13536
rect 880 13256 179120 13264
rect 880 12984 179200 13256
rect 800 12448 179200 12984
rect 800 12312 179120 12448
rect 880 12168 179120 12312
rect 880 12032 179200 12168
rect 800 11360 179200 12032
rect 880 11080 179120 11360
rect 800 10408 179200 11080
rect 880 10272 179200 10408
rect 880 10128 179120 10272
rect 800 9992 179120 10128
rect 800 9456 179200 9992
rect 880 9184 179200 9456
rect 880 9176 179120 9184
rect 800 8904 179120 9176
rect 800 8368 179200 8904
rect 880 8096 179200 8368
rect 880 8088 179120 8096
rect 800 7816 179120 8088
rect 800 7416 179200 7816
rect 880 7136 179200 7416
rect 800 7008 179200 7136
rect 800 6728 179120 7008
rect 800 6464 179200 6728
rect 880 6184 179200 6464
rect 800 5920 179200 6184
rect 800 5640 179120 5920
rect 800 5512 179200 5640
rect 880 5232 179200 5512
rect 800 4832 179200 5232
rect 800 4552 179120 4832
rect 800 4424 179200 4552
rect 880 4144 179200 4424
rect 800 3744 179200 4144
rect 800 3472 179120 3744
rect 880 3464 179120 3472
rect 880 3192 179200 3464
rect 800 2656 179200 3192
rect 800 2520 179120 2656
rect 880 2376 179120 2520
rect 880 2240 179200 2376
rect 800 1568 179200 2240
rect 880 1288 179120 1568
rect 800 616 179200 1288
rect 880 443 179120 616
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< labels >>
rlabel metal3 s 179200 11160 180000 11280 6 adc0_dat_i[0]
port 1 nsew signal input
rlabel metal3 s 179200 46792 180000 46912 6 adc0_dat_i[10]
port 2 nsew signal input
rlabel metal3 s 179200 50056 180000 50176 6 adc0_dat_i[11]
port 3 nsew signal input
rlabel metal3 s 179200 53320 180000 53440 6 adc0_dat_i[12]
port 4 nsew signal input
rlabel metal3 s 179200 56584 180000 56704 6 adc0_dat_i[13]
port 5 nsew signal input
rlabel metal3 s 179200 59848 180000 59968 6 adc0_dat_i[14]
port 6 nsew signal input
rlabel metal3 s 179200 62976 180000 63096 6 adc0_dat_i[15]
port 7 nsew signal input
rlabel metal3 s 179200 66240 180000 66360 6 adc0_dat_i[16]
port 8 nsew signal input
rlabel metal3 s 179200 69504 180000 69624 6 adc0_dat_i[17]
port 9 nsew signal input
rlabel metal3 s 179200 72768 180000 72888 6 adc0_dat_i[18]
port 10 nsew signal input
rlabel metal3 s 179200 76032 180000 76152 6 adc0_dat_i[19]
port 11 nsew signal input
rlabel metal3 s 179200 15512 180000 15632 6 adc0_dat_i[1]
port 12 nsew signal input
rlabel metal3 s 179200 79296 180000 79416 6 adc0_dat_i[20]
port 13 nsew signal input
rlabel metal3 s 179200 82424 180000 82544 6 adc0_dat_i[21]
port 14 nsew signal input
rlabel metal3 s 179200 85688 180000 85808 6 adc0_dat_i[22]
port 15 nsew signal input
rlabel metal3 s 179200 88952 180000 89072 6 adc0_dat_i[23]
port 16 nsew signal input
rlabel metal3 s 179200 92216 180000 92336 6 adc0_dat_i[24]
port 17 nsew signal input
rlabel metal3 s 179200 95480 180000 95600 6 adc0_dat_i[25]
port 18 nsew signal input
rlabel metal3 s 179200 98744 180000 98864 6 adc0_dat_i[26]
port 19 nsew signal input
rlabel metal3 s 179200 101872 180000 101992 6 adc0_dat_i[27]
port 20 nsew signal input
rlabel metal3 s 179200 105136 180000 105256 6 adc0_dat_i[28]
port 21 nsew signal input
rlabel metal3 s 179200 108400 180000 108520 6 adc0_dat_i[29]
port 22 nsew signal input
rlabel metal3 s 179200 19864 180000 19984 6 adc0_dat_i[2]
port 23 nsew signal input
rlabel metal3 s 179200 111664 180000 111784 6 adc0_dat_i[30]
port 24 nsew signal input
rlabel metal3 s 179200 114928 180000 115048 6 adc0_dat_i[31]
port 25 nsew signal input
rlabel metal3 s 179200 24080 180000 24200 6 adc0_dat_i[3]
port 26 nsew signal input
rlabel metal3 s 179200 27344 180000 27464 6 adc0_dat_i[4]
port 27 nsew signal input
rlabel metal3 s 179200 30608 180000 30728 6 adc0_dat_i[5]
port 28 nsew signal input
rlabel metal3 s 179200 33872 180000 33992 6 adc0_dat_i[6]
port 29 nsew signal input
rlabel metal3 s 179200 37136 180000 37256 6 adc0_dat_i[7]
port 30 nsew signal input
rlabel metal3 s 179200 40400 180000 40520 6 adc0_dat_i[8]
port 31 nsew signal input
rlabel metal3 s 179200 43528 180000 43648 6 adc0_dat_i[9]
port 32 nsew signal input
rlabel metal3 s 179200 12248 180000 12368 6 adc1_dat_i[0]
port 33 nsew signal input
rlabel metal3 s 179200 47880 180000 48000 6 adc1_dat_i[10]
port 34 nsew signal input
rlabel metal3 s 179200 51144 180000 51264 6 adc1_dat_i[11]
port 35 nsew signal input
rlabel metal3 s 179200 54408 180000 54528 6 adc1_dat_i[12]
port 36 nsew signal input
rlabel metal3 s 179200 57672 180000 57792 6 adc1_dat_i[13]
port 37 nsew signal input
rlabel metal3 s 179200 60800 180000 60920 6 adc1_dat_i[14]
port 38 nsew signal input
rlabel metal3 s 179200 64064 180000 64184 6 adc1_dat_i[15]
port 39 nsew signal input
rlabel metal3 s 179200 67328 180000 67448 6 adc1_dat_i[16]
port 40 nsew signal input
rlabel metal3 s 179200 70592 180000 70712 6 adc1_dat_i[17]
port 41 nsew signal input
rlabel metal3 s 179200 73856 180000 73976 6 adc1_dat_i[18]
port 42 nsew signal input
rlabel metal3 s 179200 77120 180000 77240 6 adc1_dat_i[19]
port 43 nsew signal input
rlabel metal3 s 179200 16600 180000 16720 6 adc1_dat_i[1]
port 44 nsew signal input
rlabel metal3 s 179200 80384 180000 80504 6 adc1_dat_i[20]
port 45 nsew signal input
rlabel metal3 s 179200 83512 180000 83632 6 adc1_dat_i[21]
port 46 nsew signal input
rlabel metal3 s 179200 86776 180000 86896 6 adc1_dat_i[22]
port 47 nsew signal input
rlabel metal3 s 179200 90040 180000 90160 6 adc1_dat_i[23]
port 48 nsew signal input
rlabel metal3 s 179200 93304 180000 93424 6 adc1_dat_i[24]
port 49 nsew signal input
rlabel metal3 s 179200 96568 180000 96688 6 adc1_dat_i[25]
port 50 nsew signal input
rlabel metal3 s 179200 99832 180000 99952 6 adc1_dat_i[26]
port 51 nsew signal input
rlabel metal3 s 179200 102960 180000 103080 6 adc1_dat_i[27]
port 52 nsew signal input
rlabel metal3 s 179200 106224 180000 106344 6 adc1_dat_i[28]
port 53 nsew signal input
rlabel metal3 s 179200 109488 180000 109608 6 adc1_dat_i[29]
port 54 nsew signal input
rlabel metal3 s 179200 20816 180000 20936 6 adc1_dat_i[2]
port 55 nsew signal input
rlabel metal3 s 179200 112752 180000 112872 6 adc1_dat_i[30]
port 56 nsew signal input
rlabel metal3 s 179200 116016 180000 116136 6 adc1_dat_i[31]
port 57 nsew signal input
rlabel metal3 s 179200 25168 180000 25288 6 adc1_dat_i[3]
port 58 nsew signal input
rlabel metal3 s 179200 28432 180000 28552 6 adc1_dat_i[4]
port 59 nsew signal input
rlabel metal3 s 179200 31696 180000 31816 6 adc1_dat_i[5]
port 60 nsew signal input
rlabel metal3 s 179200 34960 180000 35080 6 adc1_dat_i[6]
port 61 nsew signal input
rlabel metal3 s 179200 38224 180000 38344 6 adc1_dat_i[7]
port 62 nsew signal input
rlabel metal3 s 179200 41352 180000 41472 6 adc1_dat_i[8]
port 63 nsew signal input
rlabel metal3 s 179200 44616 180000 44736 6 adc1_dat_i[9]
port 64 nsew signal input
rlabel metal3 s 179200 13336 180000 13456 6 adc2_dat_i[0]
port 65 nsew signal input
rlabel metal3 s 179200 48968 180000 49088 6 adc2_dat_i[10]
port 66 nsew signal input
rlabel metal3 s 179200 52232 180000 52352 6 adc2_dat_i[11]
port 67 nsew signal input
rlabel metal3 s 179200 55496 180000 55616 6 adc2_dat_i[12]
port 68 nsew signal input
rlabel metal3 s 179200 58760 180000 58880 6 adc2_dat_i[13]
port 69 nsew signal input
rlabel metal3 s 179200 61888 180000 62008 6 adc2_dat_i[14]
port 70 nsew signal input
rlabel metal3 s 179200 65152 180000 65272 6 adc2_dat_i[15]
port 71 nsew signal input
rlabel metal3 s 179200 68416 180000 68536 6 adc2_dat_i[16]
port 72 nsew signal input
rlabel metal3 s 179200 71680 180000 71800 6 adc2_dat_i[17]
port 73 nsew signal input
rlabel metal3 s 179200 74944 180000 75064 6 adc2_dat_i[18]
port 74 nsew signal input
rlabel metal3 s 179200 78208 180000 78328 6 adc2_dat_i[19]
port 75 nsew signal input
rlabel metal3 s 179200 17688 180000 17808 6 adc2_dat_i[1]
port 76 nsew signal input
rlabel metal3 s 179200 81336 180000 81456 6 adc2_dat_i[20]
port 77 nsew signal input
rlabel metal3 s 179200 84600 180000 84720 6 adc2_dat_i[21]
port 78 nsew signal input
rlabel metal3 s 179200 87864 180000 87984 6 adc2_dat_i[22]
port 79 nsew signal input
rlabel metal3 s 179200 91128 180000 91248 6 adc2_dat_i[23]
port 80 nsew signal input
rlabel metal3 s 179200 94392 180000 94512 6 adc2_dat_i[24]
port 81 nsew signal input
rlabel metal3 s 179200 97656 180000 97776 6 adc2_dat_i[25]
port 82 nsew signal input
rlabel metal3 s 179200 100784 180000 100904 6 adc2_dat_i[26]
port 83 nsew signal input
rlabel metal3 s 179200 104048 180000 104168 6 adc2_dat_i[27]
port 84 nsew signal input
rlabel metal3 s 179200 107312 180000 107432 6 adc2_dat_i[28]
port 85 nsew signal input
rlabel metal3 s 179200 110576 180000 110696 6 adc2_dat_i[29]
port 86 nsew signal input
rlabel metal3 s 179200 21904 180000 22024 6 adc2_dat_i[2]
port 87 nsew signal input
rlabel metal3 s 179200 113840 180000 113960 6 adc2_dat_i[30]
port 88 nsew signal input
rlabel metal3 s 179200 117104 180000 117224 6 adc2_dat_i[31]
port 89 nsew signal input
rlabel metal3 s 179200 26256 180000 26376 6 adc2_dat_i[3]
port 90 nsew signal input
rlabel metal3 s 179200 29520 180000 29640 6 adc2_dat_i[4]
port 91 nsew signal input
rlabel metal3 s 179200 32784 180000 32904 6 adc2_dat_i[5]
port 92 nsew signal input
rlabel metal3 s 179200 36048 180000 36168 6 adc2_dat_i[6]
port 93 nsew signal input
rlabel metal3 s 179200 39312 180000 39432 6 adc2_dat_i[7]
port 94 nsew signal input
rlabel metal3 s 179200 42440 180000 42560 6 adc2_dat_i[8]
port 95 nsew signal input
rlabel metal3 s 179200 45704 180000 45824 6 adc2_dat_i[9]
port 96 nsew signal input
rlabel metal3 s 179200 14424 180000 14544 6 adc_dvalid_i[0]
port 97 nsew signal input
rlabel metal3 s 179200 18776 180000 18896 6 adc_dvalid_i[1]
port 98 nsew signal input
rlabel metal3 s 179200 22992 180000 23112 6 adc_dvalid_i[2]
port 99 nsew signal input
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 100 nsew signal input
rlabel metal2 s 45742 119200 45798 120000 6 io_in[10]
port 101 nsew signal input
rlabel metal2 s 50250 119200 50306 120000 6 io_in[11]
port 102 nsew signal input
rlabel metal2 s 54758 119200 54814 120000 6 io_in[12]
port 103 nsew signal input
rlabel metal2 s 59266 119200 59322 120000 6 io_in[13]
port 104 nsew signal input
rlabel metal2 s 63682 119200 63738 120000 6 io_in[14]
port 105 nsew signal input
rlabel metal2 s 68190 119200 68246 120000 6 io_in[15]
port 106 nsew signal input
rlabel metal2 s 72698 119200 72754 120000 6 io_in[16]
port 107 nsew signal input
rlabel metal2 s 77206 119200 77262 120000 6 io_in[17]
port 108 nsew signal input
rlabel metal2 s 81714 119200 81770 120000 6 io_in[18]
port 109 nsew signal input
rlabel metal2 s 86222 119200 86278 120000 6 io_in[19]
port 110 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[1]
port 111 nsew signal input
rlabel metal2 s 90730 119200 90786 120000 6 io_in[20]
port 112 nsew signal input
rlabel metal2 s 95238 119200 95294 120000 6 io_in[21]
port 113 nsew signal input
rlabel metal2 s 99746 119200 99802 120000 6 io_in[22]
port 114 nsew signal input
rlabel metal2 s 104254 119200 104310 120000 6 io_in[23]
port 115 nsew signal input
rlabel metal2 s 108762 119200 108818 120000 6 io_in[24]
port 116 nsew signal input
rlabel metal2 s 113270 119200 113326 120000 6 io_in[25]
port 117 nsew signal input
rlabel metal2 s 117778 119200 117834 120000 6 io_in[26]
port 118 nsew signal input
rlabel metal2 s 122194 119200 122250 120000 6 io_in[27]
port 119 nsew signal input
rlabel metal2 s 126702 119200 126758 120000 6 io_in[28]
port 120 nsew signal input
rlabel metal2 s 131210 119200 131266 120000 6 io_in[29]
port 121 nsew signal input
rlabel metal2 s 9678 119200 9734 120000 6 io_in[2]
port 122 nsew signal input
rlabel metal2 s 135718 119200 135774 120000 6 io_in[30]
port 123 nsew signal input
rlabel metal2 s 140226 119200 140282 120000 6 io_in[31]
port 124 nsew signal input
rlabel metal2 s 144734 119200 144790 120000 6 io_in[32]
port 125 nsew signal input
rlabel metal2 s 149242 119200 149298 120000 6 io_in[33]
port 126 nsew signal input
rlabel metal2 s 153750 119200 153806 120000 6 io_in[34]
port 127 nsew signal input
rlabel metal2 s 158258 119200 158314 120000 6 io_in[35]
port 128 nsew signal input
rlabel metal2 s 162766 119200 162822 120000 6 io_in[36]
port 129 nsew signal input
rlabel metal2 s 167274 119200 167330 120000 6 io_in[37]
port 130 nsew signal input
rlabel metal2 s 14186 119200 14242 120000 6 io_in[3]
port 131 nsew signal input
rlabel metal2 s 18694 119200 18750 120000 6 io_in[4]
port 132 nsew signal input
rlabel metal2 s 23202 119200 23258 120000 6 io_in[5]
port 133 nsew signal input
rlabel metal2 s 27710 119200 27766 120000 6 io_in[6]
port 134 nsew signal input
rlabel metal2 s 32218 119200 32274 120000 6 io_in[7]
port 135 nsew signal input
rlabel metal2 s 36726 119200 36782 120000 6 io_in[8]
port 136 nsew signal input
rlabel metal2 s 41234 119200 41290 120000 6 io_in[9]
port 137 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 138 nsew signal output
rlabel metal2 s 47214 119200 47270 120000 6 io_oeb[10]
port 139 nsew signal output
rlabel metal2 s 51722 119200 51778 120000 6 io_oeb[11]
port 140 nsew signal output
rlabel metal2 s 56230 119200 56286 120000 6 io_oeb[12]
port 141 nsew signal output
rlabel metal2 s 60738 119200 60794 120000 6 io_oeb[13]
port 142 nsew signal output
rlabel metal2 s 65246 119200 65302 120000 6 io_oeb[14]
port 143 nsew signal output
rlabel metal2 s 69754 119200 69810 120000 6 io_oeb[15]
port 144 nsew signal output
rlabel metal2 s 74262 119200 74318 120000 6 io_oeb[16]
port 145 nsew signal output
rlabel metal2 s 78770 119200 78826 120000 6 io_oeb[17]
port 146 nsew signal output
rlabel metal2 s 83186 119200 83242 120000 6 io_oeb[18]
port 147 nsew signal output
rlabel metal2 s 87694 119200 87750 120000 6 io_oeb[19]
port 148 nsew signal output
rlabel metal2 s 6734 119200 6790 120000 6 io_oeb[1]
port 149 nsew signal output
rlabel metal2 s 92202 119200 92258 120000 6 io_oeb[20]
port 150 nsew signal output
rlabel metal2 s 96710 119200 96766 120000 6 io_oeb[21]
port 151 nsew signal output
rlabel metal2 s 101218 119200 101274 120000 6 io_oeb[22]
port 152 nsew signal output
rlabel metal2 s 105726 119200 105782 120000 6 io_oeb[23]
port 153 nsew signal output
rlabel metal2 s 110234 119200 110290 120000 6 io_oeb[24]
port 154 nsew signal output
rlabel metal2 s 114742 119200 114798 120000 6 io_oeb[25]
port 155 nsew signal output
rlabel metal2 s 119250 119200 119306 120000 6 io_oeb[26]
port 156 nsew signal output
rlabel metal2 s 123758 119200 123814 120000 6 io_oeb[27]
port 157 nsew signal output
rlabel metal2 s 128266 119200 128322 120000 6 io_oeb[28]
port 158 nsew signal output
rlabel metal2 s 132774 119200 132830 120000 6 io_oeb[29]
port 159 nsew signal output
rlabel metal2 s 11242 119200 11298 120000 6 io_oeb[2]
port 160 nsew signal output
rlabel metal2 s 137282 119200 137338 120000 6 io_oeb[30]
port 161 nsew signal output
rlabel metal2 s 141698 119200 141754 120000 6 io_oeb[31]
port 162 nsew signal output
rlabel metal2 s 146206 119200 146262 120000 6 io_oeb[32]
port 163 nsew signal output
rlabel metal2 s 150714 119200 150770 120000 6 io_oeb[33]
port 164 nsew signal output
rlabel metal2 s 155222 119200 155278 120000 6 io_oeb[34]
port 165 nsew signal output
rlabel metal2 s 159730 119200 159786 120000 6 io_oeb[35]
port 166 nsew signal output
rlabel metal2 s 164238 119200 164294 120000 6 io_oeb[36]
port 167 nsew signal output
rlabel metal2 s 168746 119200 168802 120000 6 io_oeb[37]
port 168 nsew signal output
rlabel metal2 s 15750 119200 15806 120000 6 io_oeb[3]
port 169 nsew signal output
rlabel metal2 s 20258 119200 20314 120000 6 io_oeb[4]
port 170 nsew signal output
rlabel metal2 s 24674 119200 24730 120000 6 io_oeb[5]
port 171 nsew signal output
rlabel metal2 s 29182 119200 29238 120000 6 io_oeb[6]
port 172 nsew signal output
rlabel metal2 s 33690 119200 33746 120000 6 io_oeb[7]
port 173 nsew signal output
rlabel metal2 s 38198 119200 38254 120000 6 io_oeb[8]
port 174 nsew signal output
rlabel metal2 s 42706 119200 42762 120000 6 io_oeb[9]
port 175 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 176 nsew signal output
rlabel metal2 s 48686 119200 48742 120000 6 io_out[10]
port 177 nsew signal output
rlabel metal2 s 53194 119200 53250 120000 6 io_out[11]
port 178 nsew signal output
rlabel metal2 s 57702 119200 57758 120000 6 io_out[12]
port 179 nsew signal output
rlabel metal2 s 62210 119200 62266 120000 6 io_out[13]
port 180 nsew signal output
rlabel metal2 s 66718 119200 66774 120000 6 io_out[14]
port 181 nsew signal output
rlabel metal2 s 71226 119200 71282 120000 6 io_out[15]
port 182 nsew signal output
rlabel metal2 s 75734 119200 75790 120000 6 io_out[16]
port 183 nsew signal output
rlabel metal2 s 80242 119200 80298 120000 6 io_out[17]
port 184 nsew signal output
rlabel metal2 s 84750 119200 84806 120000 6 io_out[18]
port 185 nsew signal output
rlabel metal2 s 89258 119200 89314 120000 6 io_out[19]
port 186 nsew signal output
rlabel metal2 s 8206 119200 8262 120000 6 io_out[1]
port 187 nsew signal output
rlabel metal2 s 93766 119200 93822 120000 6 io_out[20]
port 188 nsew signal output
rlabel metal2 s 98274 119200 98330 120000 6 io_out[21]
port 189 nsew signal output
rlabel metal2 s 102690 119200 102746 120000 6 io_out[22]
port 190 nsew signal output
rlabel metal2 s 107198 119200 107254 120000 6 io_out[23]
port 191 nsew signal output
rlabel metal2 s 111706 119200 111762 120000 6 io_out[24]
port 192 nsew signal output
rlabel metal2 s 116214 119200 116270 120000 6 io_out[25]
port 193 nsew signal output
rlabel metal2 s 120722 119200 120778 120000 6 io_out[26]
port 194 nsew signal output
rlabel metal2 s 125230 119200 125286 120000 6 io_out[27]
port 195 nsew signal output
rlabel metal2 s 129738 119200 129794 120000 6 io_out[28]
port 196 nsew signal output
rlabel metal2 s 134246 119200 134302 120000 6 io_out[29]
port 197 nsew signal output
rlabel metal2 s 12714 119200 12770 120000 6 io_out[2]
port 198 nsew signal output
rlabel metal2 s 138754 119200 138810 120000 6 io_out[30]
port 199 nsew signal output
rlabel metal2 s 143262 119200 143318 120000 6 io_out[31]
port 200 nsew signal output
rlabel metal2 s 147770 119200 147826 120000 6 io_out[32]
port 201 nsew signal output
rlabel metal2 s 152278 119200 152334 120000 6 io_out[33]
port 202 nsew signal output
rlabel metal2 s 156786 119200 156842 120000 6 io_out[34]
port 203 nsew signal output
rlabel metal2 s 161202 119200 161258 120000 6 io_out[35]
port 204 nsew signal output
rlabel metal2 s 165710 119200 165766 120000 6 io_out[36]
port 205 nsew signal output
rlabel metal2 s 170218 119200 170274 120000 6 io_out[37]
port 206 nsew signal output
rlabel metal2 s 17222 119200 17278 120000 6 io_out[3]
port 207 nsew signal output
rlabel metal2 s 21730 119200 21786 120000 6 io_out[4]
port 208 nsew signal output
rlabel metal2 s 26238 119200 26294 120000 6 io_out[5]
port 209 nsew signal output
rlabel metal2 s 30746 119200 30802 120000 6 io_out[6]
port 210 nsew signal output
rlabel metal2 s 35254 119200 35310 120000 6 io_out[7]
port 211 nsew signal output
rlabel metal2 s 39762 119200 39818 120000 6 io_out[8]
port 212 nsew signal output
rlabel metal2 s 44178 119200 44234 120000 6 io_out[9]
port 213 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 irq[0]
port 214 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 irq[1]
port 215 nsew signal output
rlabel metal3 s 179200 119280 180000 119400 6 irq[2]
port 216 nsew signal output
rlabel metal3 s 0 416 800 536 6 mem1_data_i[0]
port 217 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 mem1_data_i[10]
port 218 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 mem1_data_i[11]
port 219 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 mem1_data_i[12]
port 220 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 mem1_data_i[13]
port 221 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 mem1_data_i[14]
port 222 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 mem1_data_i[15]
port 223 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 mem1_data_i[16]
port 224 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 mem1_data_i[17]
port 225 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 mem1_data_i[18]
port 226 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 mem1_data_i[19]
port 227 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 mem1_data_i[1]
port 228 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 mem1_data_i[20]
port 229 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 mem1_data_i[21]
port 230 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 mem1_data_i[22]
port 231 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 mem1_data_i[23]
port 232 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 mem1_data_i[24]
port 233 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 mem1_data_i[25]
port 234 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 mem1_data_i[26]
port 235 nsew signal input
rlabel metal3 s 0 101600 800 101720 6 mem1_data_i[27]
port 236 nsew signal input
rlabel metal3 s 0 104592 800 104712 6 mem1_data_i[28]
port 237 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 mem1_data_i[29]
port 238 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 mem1_data_i[2]
port 239 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 mem1_data_i[30]
port 240 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 mem1_data_i[31]
port 241 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 mem1_data_i[3]
port 242 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 mem1_data_i[4]
port 243 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 mem1_data_i[5]
port 244 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 mem1_data_i[6]
port 245 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 mem1_data_i[7]
port 246 nsew signal input
rlabel metal3 s 0 43664 800 43784 6 mem1_data_i[8]
port 247 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 mem1_data_i[9]
port 248 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 mem_data_i[0]
port 249 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 mem_data_i[10]
port 250 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 mem_data_i[11]
port 251 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 mem_data_i[12]
port 252 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 mem_data_i[13]
port 253 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 mem_data_i[14]
port 254 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 mem_data_i[15]
port 255 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 mem_data_i[16]
port 256 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 mem_data_i[17]
port 257 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 mem_data_i[18]
port 258 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 mem_data_i[19]
port 259 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 mem_data_i[1]
port 260 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 mem_data_i[20]
port 261 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 mem_data_i[21]
port 262 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 mem_data_i[22]
port 263 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 mem_data_i[23]
port 264 nsew signal input
rlabel metal3 s 0 93712 800 93832 6 mem_data_i[24]
port 265 nsew signal input
rlabel metal3 s 0 96704 800 96824 6 mem_data_i[25]
port 266 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 mem_data_i[26]
port 267 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 mem_data_i[27]
port 268 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 mem_data_i[28]
port 269 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 mem_data_i[29]
port 270 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 mem_data_i[2]
port 271 nsew signal input
rlabel metal3 s 0 111392 800 111512 6 mem_data_i[30]
port 272 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 mem_data_i[31]
port 273 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 mem_data_i[3]
port 274 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 mem_data_i[4]
port 275 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 mem_data_i[5]
port 276 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 mem_data_i[6]
port 277 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 mem_data_i[7]
port 278 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 mem_data_i[8]
port 279 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 mem_data_i[9]
port 280 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 mem_data_o[0]
port 281 nsew signal output
rlabel metal3 s 0 53456 800 53576 6 mem_data_o[10]
port 282 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 mem_data_o[11]
port 283 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 mem_data_o[12]
port 284 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 mem_data_o[13]
port 285 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 mem_data_o[14]
port 286 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 mem_data_o[15]
port 287 nsew signal output
rlabel metal3 s 0 71136 800 71256 6 mem_data_o[16]
port 288 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 mem_data_o[17]
port 289 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 mem_data_o[18]
port 290 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 mem_data_o[19]
port 291 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 mem_data_o[1]
port 292 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 mem_data_o[20]
port 293 nsew signal output
rlabel metal3 s 0 85824 800 85944 6 mem_data_o[21]
port 294 nsew signal output
rlabel metal3 s 0 88816 800 88936 6 mem_data_o[22]
port 295 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 mem_data_o[23]
port 296 nsew signal output
rlabel metal3 s 0 94800 800 94920 6 mem_data_o[24]
port 297 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 mem_data_o[25]
port 298 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 mem_data_o[26]
port 299 nsew signal output
rlabel metal3 s 0 103640 800 103760 6 mem_data_o[27]
port 300 nsew signal output
rlabel metal3 s 0 106496 800 106616 6 mem_data_o[28]
port 301 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 mem_data_o[29]
port 302 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 mem_data_o[2]
port 303 nsew signal output
rlabel metal3 s 0 112480 800 112600 6 mem_data_o[30]
port 304 nsew signal output
rlabel metal3 s 0 115336 800 115456 6 mem_data_o[31]
port 305 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 mem_data_o[3]
port 306 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 mem_data_o[4]
port 307 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 mem_data_o[5]
port 308 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 mem_data_o[6]
port 309 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 mem_data_o[7]
port 310 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 mem_data_o[8]
port 311 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 mem_data_o[9]
port 312 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 mem_raddr_o[0]
port 313 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 mem_raddr_o[1]
port 314 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 mem_raddr_o[2]
port 315 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 mem_raddr_o[3]
port 316 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 mem_raddr_o[4]
port 317 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 mem_raddr_o[5]
port 318 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 mem_raddr_o[6]
port 319 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 mem_raddr_o[7]
port 320 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 mem_raddr_o[8]
port 321 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 mem_renb_o[0]
port 322 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 mem_renb_o[1]
port 323 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 mem_waddr_o[0]
port 324 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 mem_waddr_o[1]
port 325 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 mem_waddr_o[2]
port 326 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 mem_waddr_o[3]
port 327 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 mem_waddr_o[4]
port 328 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 mem_waddr_o[5]
port 329 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 mem_waddr_o[6]
port 330 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 mem_waddr_o[7]
port 331 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 mem_waddr_o[8]
port 332 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 mem_wenb_o[0]
port 333 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 mem_wenb_o[1]
port 334 nsew signal output
rlabel metal3 s 179200 416 180000 536 6 oversample_o[0]
port 335 nsew signal output
rlabel metal3 s 179200 1368 180000 1488 6 oversample_o[1]
port 336 nsew signal output
rlabel metal3 s 179200 2456 180000 2576 6 oversample_o[2]
port 337 nsew signal output
rlabel metal3 s 179200 3544 180000 3664 6 oversample_o[3]
port 338 nsew signal output
rlabel metal3 s 179200 4632 180000 4752 6 oversample_o[4]
port 339 nsew signal output
rlabel metal3 s 179200 5720 180000 5840 6 oversample_o[5]
port 340 nsew signal output
rlabel metal3 s 179200 6808 180000 6928 6 oversample_o[6]
port 341 nsew signal output
rlabel metal3 s 179200 7896 180000 8016 6 oversample_o[7]
port 342 nsew signal output
rlabel metal3 s 179200 8984 180000 9104 6 oversample_o[8]
port 343 nsew signal output
rlabel metal3 s 179200 10072 180000 10192 6 oversample_o[9]
port 344 nsew signal output
rlabel metal2 s 176290 119200 176346 120000 6 sinc3_en_o[0]
port 345 nsew signal output
rlabel metal2 s 177762 119200 177818 120000 6 sinc3_en_o[1]
port 346 nsew signal output
rlabel metal2 s 179234 119200 179290 120000 6 sinc3_en_o[2]
port 347 nsew signal output
rlabel metal2 s 171782 119200 171838 120000 6 vco_enb_o[0]
port 348 nsew signal output
rlabel metal2 s 173254 119200 173310 120000 6 vco_enb_o[1]
port 349 nsew signal output
rlabel metal2 s 174726 119200 174782 120000 6 vco_enb_o[2]
port 350 nsew signal output
rlabel metal2 s 846 0 902 800 6 wb_clk_i
port 351 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wb_rst_i
port 352 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_ack_o
port 353 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_adr_i[0]
port 354 nsew signal input
rlabel metal2 s 68098 0 68154 800 6 wbs_adr_i[10]
port 355 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 wbs_adr_i[11]
port 356 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 wbs_adr_i[12]
port 357 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 wbs_adr_i[13]
port 358 nsew signal input
rlabel metal2 s 88338 0 88394 800 6 wbs_adr_i[14]
port 359 nsew signal input
rlabel metal2 s 93306 0 93362 800 6 wbs_adr_i[15]
port 360 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 wbs_adr_i[16]
port 361 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 wbs_adr_i[17]
port 362 nsew signal input
rlabel metal2 s 108486 0 108542 800 6 wbs_adr_i[18]
port 363 nsew signal input
rlabel metal2 s 113546 0 113602 800 6 wbs_adr_i[19]
port 364 nsew signal input
rlabel metal2 s 17590 0 17646 800 6 wbs_adr_i[1]
port 365 nsew signal input
rlabel metal2 s 118606 0 118662 800 6 wbs_adr_i[20]
port 366 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 wbs_adr_i[21]
port 367 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 wbs_adr_i[22]
port 368 nsew signal input
rlabel metal2 s 133694 0 133750 800 6 wbs_adr_i[23]
port 369 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 wbs_adr_i[24]
port 370 nsew signal input
rlabel metal2 s 143814 0 143870 800 6 wbs_adr_i[25]
port 371 nsew signal input
rlabel metal2 s 148874 0 148930 800 6 wbs_adr_i[26]
port 372 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 wbs_adr_i[27]
port 373 nsew signal input
rlabel metal2 s 158994 0 159050 800 6 wbs_adr_i[28]
port 374 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 wbs_adr_i[29]
port 375 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[2]
port 376 nsew signal input
rlabel metal2 s 169022 0 169078 800 6 wbs_adr_i[30]
port 377 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 wbs_adr_i[31]
port 378 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 wbs_adr_i[3]
port 379 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 wbs_adr_i[4]
port 380 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[5]
port 381 nsew signal input
rlabel metal2 s 47950 0 48006 800 6 wbs_adr_i[6]
port 382 nsew signal input
rlabel metal2 s 52918 0 52974 800 6 wbs_adr_i[7]
port 383 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 wbs_adr_i[8]
port 384 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_adr_i[9]
port 385 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_cyc_i
port 386 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_i[0]
port 387 nsew signal input
rlabel metal2 s 69754 0 69810 800 6 wbs_dat_i[10]
port 388 nsew signal input
rlabel metal2 s 74814 0 74870 800 6 wbs_dat_i[11]
port 389 nsew signal input
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_i[12]
port 390 nsew signal input
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_i[13]
port 391 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_i[14]
port 392 nsew signal input
rlabel metal2 s 95054 0 95110 800 6 wbs_dat_i[15]
port 393 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 wbs_dat_i[16]
port 394 nsew signal input
rlabel metal2 s 105082 0 105138 800 6 wbs_dat_i[17]
port 395 nsew signal input
rlabel metal2 s 110142 0 110198 800 6 wbs_dat_i[18]
port 396 nsew signal input
rlabel metal2 s 115202 0 115258 800 6 wbs_dat_i[19]
port 397 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 wbs_dat_i[1]
port 398 nsew signal input
rlabel metal2 s 120262 0 120318 800 6 wbs_dat_i[20]
port 399 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 wbs_dat_i[21]
port 400 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 wbs_dat_i[22]
port 401 nsew signal input
rlabel metal2 s 135442 0 135498 800 6 wbs_dat_i[23]
port 402 nsew signal input
rlabel metal2 s 140502 0 140558 800 6 wbs_dat_i[24]
port 403 nsew signal input
rlabel metal2 s 145470 0 145526 800 6 wbs_dat_i[25]
port 404 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 wbs_dat_i[26]
port 405 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 wbs_dat_i[27]
port 406 nsew signal input
rlabel metal2 s 160650 0 160706 800 6 wbs_dat_i[28]
port 407 nsew signal input
rlabel metal2 s 165710 0 165766 800 6 wbs_dat_i[29]
port 408 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 wbs_dat_i[2]
port 409 nsew signal input
rlabel metal2 s 170770 0 170826 800 6 wbs_dat_i[30]
port 410 nsew signal input
rlabel metal2 s 175830 0 175886 800 6 wbs_dat_i[31]
port 411 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 wbs_dat_i[3]
port 412 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 wbs_dat_i[4]
port 413 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 wbs_dat_i[5]
port 414 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[6]
port 415 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 wbs_dat_i[7]
port 416 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_i[8]
port 417 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 wbs_dat_i[9]
port 418 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_o[0]
port 419 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 wbs_dat_o[10]
port 420 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 wbs_dat_o[11]
port 421 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 wbs_dat_o[12]
port 422 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_o[13]
port 423 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 wbs_dat_o[14]
port 424 nsew signal output
rlabel metal2 s 96710 0 96766 800 6 wbs_dat_o[15]
port 425 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 wbs_dat_o[16]
port 426 nsew signal output
rlabel metal2 s 106830 0 106886 800 6 wbs_dat_o[17]
port 427 nsew signal output
rlabel metal2 s 111890 0 111946 800 6 wbs_dat_o[18]
port 428 nsew signal output
rlabel metal2 s 116858 0 116914 800 6 wbs_dat_o[19]
port 429 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 wbs_dat_o[1]
port 430 nsew signal output
rlabel metal2 s 121918 0 121974 800 6 wbs_dat_o[20]
port 431 nsew signal output
rlabel metal2 s 126978 0 127034 800 6 wbs_dat_o[21]
port 432 nsew signal output
rlabel metal2 s 132038 0 132094 800 6 wbs_dat_o[22]
port 433 nsew signal output
rlabel metal2 s 137098 0 137154 800 6 wbs_dat_o[23]
port 434 nsew signal output
rlabel metal2 s 142158 0 142214 800 6 wbs_dat_o[24]
port 435 nsew signal output
rlabel metal2 s 147218 0 147274 800 6 wbs_dat_o[25]
port 436 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 wbs_dat_o[26]
port 437 nsew signal output
rlabel metal2 s 157246 0 157302 800 6 wbs_dat_o[27]
port 438 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 wbs_dat_o[28]
port 439 nsew signal output
rlabel metal2 s 167366 0 167422 800 6 wbs_dat_o[29]
port 440 nsew signal output
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_o[2]
port 441 nsew signal output
rlabel metal2 s 172426 0 172482 800 6 wbs_dat_o[30]
port 442 nsew signal output
rlabel metal2 s 177486 0 177542 800 6 wbs_dat_o[31]
port 443 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 wbs_dat_o[3]
port 444 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 wbs_dat_o[4]
port 445 nsew signal output
rlabel metal2 s 46202 0 46258 800 6 wbs_dat_o[5]
port 446 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[6]
port 447 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 wbs_dat_o[7]
port 448 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 wbs_dat_o[8]
port 449 nsew signal output
rlabel metal2 s 66442 0 66498 800 6 wbs_dat_o[9]
port 450 nsew signal output
rlabel metal2 s 15934 0 15990 800 6 wbs_sel_i[0]
port 451 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 wbs_sel_i[1]
port 452 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wbs_sel_i[2]
port 453 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_sel_i[3]
port 454 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_stb_i
port 455 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_we_i
port 456 nsew signal input
rlabel metal3 s 0 117376 800 117496 6 wmask_o[0]
port 457 nsew signal output
rlabel metal3 s 179200 118192 180000 118312 6 wmask_o[1]
port 458 nsew signal output
rlabel metal3 s 0 119280 800 119400 6 wmask_o[2]
port 459 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 wmask_o[3]
port 460 nsew signal output
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 461 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 462 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 463 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 464 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 465 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 466 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 467 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 468 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 469 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 470 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 471 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 472 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 473 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 474 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 475 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 476 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 477 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 478 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 479 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 480 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 481 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 482 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 483 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 484 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 485 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 486 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 487 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 488 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 489 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 490 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 491 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 492 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 493 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 494 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 495 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 496 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 497 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 498 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 499 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 500 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 501 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 502 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 503 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 504 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 505 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 506 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 507 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 508 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 9222838
string GDS_START 666706
<< end >>

