module user_project_wrapper (user_clock2,
    wb_clk_i,
    wb_rst_i,
    wbs_ack_o,
    wbs_cyc_i,
    wbs_stb_i,
    wbs_we_i,
    vccd1,
    vssd1,
    vccd2,
    vssd2,
    vdda1,
    vssa1,
    vdda2,
    vssa2,
    analog_io,
    io_in,
    io_oeb,
    io_out,
    la_data_in,
    la_data_out,
    la_oenb,
    user_irq,
    wbs_adr_i,
    wbs_dat_i,
    wbs_dat_o,
    wbs_sel_i);
 input user_clock2;
 input wb_clk_i;
 input wb_rst_i;
 output wbs_ack_o;
 input wbs_cyc_i;
 input wbs_stb_i;
 input wbs_we_i;
 input vccd1;
 input vssd1;
 input vccd2;
 input vssd2;
 input vdda1;
 input vssa1;
 input vdda2;
 input vssa2;
 inout [28:0] analog_io;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;
 input [127:0] la_data_in;
 output [127:0] la_data_out;
 input [127:0] la_oenb;
 output [2:0] user_irq;
 input [31:0] wbs_adr_i;
 input [31:0] wbs_dat_i;
 output [31:0] wbs_dat_o;
 input [3:0] wbs_sel_i;

 sky130_sram_2kbyte_1rw1r_32x512_8 mem_0 (.csb0(\wenb[0] ),
    .csb1(\renb[0] ),
    .web0(\wenb[0] ),
    .clk0(wb_clk_i),
    .clk1(wb_clk_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\waddr[8] ,
    \waddr[7] ,
    \waddr[6] ,
    \waddr[5] ,
    \waddr[4] ,
    \waddr[3] ,
    \waddr[2] ,
    \waddr[1] ,
    \waddr[0] }),
    .addr1({\raddr[8] ,
    \raddr[7] ,
    \raddr[6] ,
    \raddr[5] ,
    \raddr[4] ,
    \raddr[3] ,
    \raddr[2] ,
    \raddr[1] ,
    \raddr[0] }),
    .din0({\w2m_data[31] ,
    \w2m_data[30] ,
    \w2m_data[29] ,
    \w2m_data[28] ,
    \w2m_data[27] ,
    \w2m_data[26] ,
    \w2m_data[25] ,
    \w2m_data[24] ,
    \w2m_data[23] ,
    \w2m_data[22] ,
    \w2m_data[21] ,
    \w2m_data[20] ,
    \w2m_data[19] ,
    \w2m_data[18] ,
    \w2m_data[17] ,
    \w2m_data[16] ,
    \w2m_data[15] ,
    \w2m_data[14] ,
    \w2m_data[13] ,
    \w2m_data[12] ,
    \w2m_data[11] ,
    \w2m_data[10] ,
    \w2m_data[9] ,
    \w2m_data[8] ,
    \w2m_data[7] ,
    \w2m_data[6] ,
    \w2m_data[5] ,
    \w2m_data[4] ,
    \w2m_data[3] ,
    \w2m_data[2] ,
    \w2m_data[1] ,
    \w2m_data[0] }),
    .dout0({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .dout1({\m2w_data0[31] ,
    \m2w_data0[30] ,
    \m2w_data0[29] ,
    \m2w_data0[28] ,
    \m2w_data0[27] ,
    \m2w_data0[26] ,
    \m2w_data0[25] ,
    \m2w_data0[24] ,
    \m2w_data0[23] ,
    \m2w_data0[22] ,
    \m2w_data0[21] ,
    \m2w_data0[20] ,
    \m2w_data0[19] ,
    \m2w_data0[18] ,
    \m2w_data0[17] ,
    \m2w_data0[16] ,
    \m2w_data0[15] ,
    \m2w_data0[14] ,
    \m2w_data0[13] ,
    \m2w_data0[12] ,
    \m2w_data0[11] ,
    \m2w_data0[10] ,
    \m2w_data0[9] ,
    \m2w_data0[8] ,
    \m2w_data0[7] ,
    \m2w_data0[6] ,
    \m2w_data0[5] ,
    \m2w_data0[4] ,
    \m2w_data0[3] ,
    \m2w_data0[2] ,
    \m2w_data0[1] ,
    \m2w_data0[0] }),
    .wmask0({\wmask[3] ,
    \wmask[2] ,
    \wmask[1] ,
    \wmask[0] }));
 sky130_sram_2kbyte_1rw1r_32x512_8 mem_1 (.csb0(\wenb[1] ),
    .csb1(\renb[1] ),
    .web0(\wenb[1] ),
    .clk0(wb_clk_i),
    .clk1(wb_clk_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .addr0({\waddr[8] ,
    \waddr[7] ,
    \waddr[6] ,
    \waddr[5] ,
    \waddr[4] ,
    \waddr[3] ,
    \waddr[2] ,
    \waddr[1] ,
    \waddr[0] }),
    .addr1({\raddr[8] ,
    \raddr[7] ,
    \raddr[6] ,
    \raddr[5] ,
    \raddr[4] ,
    \raddr[3] ,
    \raddr[2] ,
    \raddr[1] ,
    \raddr[0] }),
    .din0({\w2m_data[31] ,
    \w2m_data[30] ,
    \w2m_data[29] ,
    \w2m_data[28] ,
    \w2m_data[27] ,
    \w2m_data[26] ,
    \w2m_data[25] ,
    \w2m_data[24] ,
    \w2m_data[23] ,
    \w2m_data[22] ,
    \w2m_data[21] ,
    \w2m_data[20] ,
    \w2m_data[19] ,
    \w2m_data[18] ,
    \w2m_data[17] ,
    \w2m_data[16] ,
    \w2m_data[15] ,
    \w2m_data[14] ,
    \w2m_data[13] ,
    \w2m_data[12] ,
    \w2m_data[11] ,
    \w2m_data[10] ,
    \w2m_data[9] ,
    \w2m_data[8] ,
    \w2m_data[7] ,
    \w2m_data[6] ,
    \w2m_data[5] ,
    \w2m_data[4] ,
    \w2m_data[3] ,
    \w2m_data[2] ,
    \w2m_data[1] ,
    \w2m_data[0] }),
    .dout0({_NC33,
    _NC34,
    _NC35,
    _NC36,
    _NC37,
    _NC38,
    _NC39,
    _NC40,
    _NC41,
    _NC42,
    _NC43,
    _NC44,
    _NC45,
    _NC46,
    _NC47,
    _NC48,
    _NC49,
    _NC50,
    _NC51,
    _NC52,
    _NC53,
    _NC54,
    _NC55,
    _NC56,
    _NC57,
    _NC58,
    _NC59,
    _NC60,
    _NC61,
    _NC62,
    _NC63,
    _NC64}),
    .dout1({\m2w_data1[31] ,
    \m2w_data1[30] ,
    \m2w_data1[29] ,
    \m2w_data1[28] ,
    \m2w_data1[27] ,
    \m2w_data1[26] ,
    \m2w_data1[25] ,
    \m2w_data1[24] ,
    \m2w_data1[23] ,
    \m2w_data1[22] ,
    \m2w_data1[21] ,
    \m2w_data1[20] ,
    \m2w_data1[19] ,
    \m2w_data1[18] ,
    \m2w_data1[17] ,
    \m2w_data1[16] ,
    \m2w_data1[15] ,
    \m2w_data1[14] ,
    \m2w_data1[13] ,
    \m2w_data1[12] ,
    \m2w_data1[11] ,
    \m2w_data1[10] ,
    \m2w_data1[9] ,
    \m2w_data1[8] ,
    \m2w_data1[7] ,
    \m2w_data1[6] ,
    \m2w_data1[5] ,
    \m2w_data1[4] ,
    \m2w_data1[3] ,
    \m2w_data1[2] ,
    \m2w_data1[1] ,
    \m2w_data1[0] }),
    .wmask0({\wmask[3] ,
    \wmask[2] ,
    \wmask[1] ,
    \wmask[0] }));
 vco_r100 vco_0 (.input_analog(analog_io[9]),
    .vccd2(vccd2),
    .vssd2(vssd2),
    .enb(\vco_enb[0] ),
    .p({\phase0[10] ,
    \phase0[9] ,
    \phase0[8] ,
    \phase0[7] ,
    analog_io[10],
    \phase0[5] ,
    \phase0[4] ,
    \phase0[3] ,
    \phase0[2] ,
    \phase0[1] ,
    \phase0[0] }));
 vco vco_1 (.input_analog(analog_io[12]),
    .vccd2(vccd2),
    .vssd2(vssd2),
    .enb(\vco_enb[1] ),
    .p({\phase1[10] ,
    \phase1[9] ,
    \phase1[8] ,
    \phase1[7] ,
    analog_io[13],
    \phase1[5] ,
    \phase1[4] ,
    \phase1[3] ,
    \phase1[2] ,
    \phase1[1] ,
    \phase1[0] }));
 vco_r100 vco_2 (.input_analog(analog_io[15]),
    .vccd2(vccd2),
    .vssd2(vssd2),
    .enb(\vco_enb[2] ),
    .p({\phase2[10] ,
    \phase2[9] ,
    \phase2[8] ,
    \phase2[7] ,
    analog_io[16],
    \phase2[5] ,
    \phase2[4] ,
    \phase2[3] ,
    \phase2[2] ,
    \phase2[1] ,
    \phase2[0] }));
 vco_adc vco_adc_0 (.clk(wb_clk_i),
    .data_valid_out(\sinc3_dvalid[0] ),
    .enable_in(\en[0] ),
    .rst(wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .data_out({\adc_out_0[31] ,
    \adc_out_0[30] ,
    \adc_out_0[29] ,
    \adc_out_0[28] ,
    \adc_out_0[27] ,
    \adc_out_0[26] ,
    \adc_out_0[25] ,
    \adc_out_0[24] ,
    \adc_out_0[23] ,
    \adc_out_0[22] ,
    \adc_out_0[21] ,
    \adc_out_0[20] ,
    \adc_out_0[19] ,
    \adc_out_0[18] ,
    \adc_out_0[17] ,
    \adc_out_0[16] ,
    \adc_out_0[15] ,
    \adc_out_0[14] ,
    \adc_out_0[13] ,
    \adc_out_0[12] ,
    \adc_out_0[11] ,
    \adc_out_0[10] ,
    \adc_out_0[9] ,
    \adc_out_0[8] ,
    \adc_out_0[7] ,
    \adc_out_0[6] ,
    \adc_out_0[5] ,
    \adc_out_0[4] ,
    \adc_out_0[3] ,
    \adc_out_0[2] ,
    \adc_out_0[1] ,
    \adc_out_0[0] }),
    .oversample_in({\oversample[9] ,
    \oversample[8] ,
    \oversample[7] ,
    \oversample[6] ,
    \oversample[5] ,
    \oversample[4] ,
    \oversample[3] ,
    \oversample[2] ,
    \oversample[1] ,
    \oversample[0] }),
    .phase_in({\phase0[10] ,
    \phase0[9] ,
    \phase0[8] ,
    \phase0[7] ,
    analog_io[10],
    \phase0[5] ,
    \phase0[4] ,
    \phase0[3] ,
    \phase0[2] ,
    \phase0[1] ,
    \phase0[0] }));
 vco_adc vco_adc_1 (.clk(wb_clk_i),
    .data_valid_out(\sinc3_dvalid[1] ),
    .enable_in(\en[1] ),
    .rst(wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .data_out({\adc_out_1[31] ,
    \adc_out_1[30] ,
    \adc_out_1[29] ,
    \adc_out_1[28] ,
    \adc_out_1[27] ,
    \adc_out_1[26] ,
    \adc_out_1[25] ,
    \adc_out_1[24] ,
    \adc_out_1[23] ,
    \adc_out_1[22] ,
    \adc_out_1[21] ,
    \adc_out_1[20] ,
    \adc_out_1[19] ,
    \adc_out_1[18] ,
    \adc_out_1[17] ,
    \adc_out_1[16] ,
    \adc_out_1[15] ,
    \adc_out_1[14] ,
    \adc_out_1[13] ,
    \adc_out_1[12] ,
    \adc_out_1[11] ,
    \adc_out_1[10] ,
    \adc_out_1[9] ,
    \adc_out_1[8] ,
    \adc_out_1[7] ,
    \adc_out_1[6] ,
    \adc_out_1[5] ,
    \adc_out_1[4] ,
    \adc_out_1[3] ,
    \adc_out_1[2] ,
    \adc_out_1[1] ,
    \adc_out_1[0] }),
    .oversample_in({\oversample[9] ,
    \oversample[8] ,
    \oversample[7] ,
    \oversample[6] ,
    \oversample[5] ,
    \oversample[4] ,
    \oversample[3] ,
    \oversample[2] ,
    \oversample[1] ,
    \oversample[0] }),
    .phase_in({\phase1[10] ,
    \phase1[9] ,
    \phase1[8] ,
    \phase1[7] ,
    analog_io[13],
    \phase1[5] ,
    \phase1[4] ,
    \phase1[3] ,
    \phase1[2] ,
    \phase1[1] ,
    \phase1[0] }));
 vco_adc vco_adc_2 (.clk(wb_clk_i),
    .data_valid_out(\sinc3_dvalid[2] ),
    .enable_in(\en[2] ),
    .rst(wb_rst_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .data_out({\adc_out_2[31] ,
    \adc_out_2[30] ,
    \adc_out_2[29] ,
    \adc_out_2[28] ,
    \adc_out_2[27] ,
    \adc_out_2[26] ,
    \adc_out_2[25] ,
    \adc_out_2[24] ,
    \adc_out_2[23] ,
    \adc_out_2[22] ,
    \adc_out_2[21] ,
    \adc_out_2[20] ,
    \adc_out_2[19] ,
    \adc_out_2[18] ,
    \adc_out_2[17] ,
    \adc_out_2[16] ,
    \adc_out_2[15] ,
    \adc_out_2[14] ,
    \adc_out_2[13] ,
    \adc_out_2[12] ,
    \adc_out_2[11] ,
    \adc_out_2[10] ,
    \adc_out_2[9] ,
    \adc_out_2[8] ,
    \adc_out_2[7] ,
    \adc_out_2[6] ,
    \adc_out_2[5] ,
    \adc_out_2[4] ,
    \adc_out_2[3] ,
    \adc_out_2[2] ,
    \adc_out_2[1] ,
    \adc_out_2[0] }),
    .oversample_in({\oversample[9] ,
    \oversample[8] ,
    \oversample[7] ,
    \oversample[6] ,
    \oversample[5] ,
    \oversample[4] ,
    \oversample[3] ,
    \oversample[2] ,
    \oversample[1] ,
    \oversample[0] }),
    .phase_in({\phase2[10] ,
    \phase2[9] ,
    \phase2[8] ,
    \phase2[7] ,
    analog_io[16],
    \phase2[5] ,
    \phase2[4] ,
    \phase2[3] ,
    \phase2[2] ,
    \phase2[1] ,
    \phase2[0] }));
 vco_adc_wrapper vco_adc_wrapper_1 (.wb_clk_i(wb_clk_i),
    .wb_rst_i(wb_rst_i),
    .wbs_ack_o(wbs_ack_o),
    .wbs_cyc_i(wbs_cyc_i),
    .wbs_stb_i(wbs_stb_i),
    .wbs_we_i(wbs_we_i),
    .vccd1(vccd1),
    .vssd1(vssd1),
    .vccd2(vccd2),
    .vssd2(vssd2),
    .vdda1(vdda1),
    .vssa1(vssa1),
    .vdda2(vdda2),
    .vssa2(vssa2),
    .adc0_dat_i({\adc_out_0[31] ,
    \adc_out_0[30] ,
    \adc_out_0[29] ,
    \adc_out_0[28] ,
    \adc_out_0[27] ,
    \adc_out_0[26] ,
    \adc_out_0[25] ,
    \adc_out_0[24] ,
    \adc_out_0[23] ,
    \adc_out_0[22] ,
    \adc_out_0[21] ,
    \adc_out_0[20] ,
    \adc_out_0[19] ,
    \adc_out_0[18] ,
    \adc_out_0[17] ,
    \adc_out_0[16] ,
    \adc_out_0[15] ,
    \adc_out_0[14] ,
    \adc_out_0[13] ,
    \adc_out_0[12] ,
    \adc_out_0[11] ,
    \adc_out_0[10] ,
    \adc_out_0[9] ,
    \adc_out_0[8] ,
    \adc_out_0[7] ,
    \adc_out_0[6] ,
    \adc_out_0[5] ,
    \adc_out_0[4] ,
    \adc_out_0[3] ,
    \adc_out_0[2] ,
    \adc_out_0[1] ,
    \adc_out_0[0] }),
    .adc1_dat_i({\adc_out_1[31] ,
    \adc_out_1[30] ,
    \adc_out_1[29] ,
    \adc_out_1[28] ,
    \adc_out_1[27] ,
    \adc_out_1[26] ,
    \adc_out_1[25] ,
    \adc_out_1[24] ,
    \adc_out_1[23] ,
    \adc_out_1[22] ,
    \adc_out_1[21] ,
    \adc_out_1[20] ,
    \adc_out_1[19] ,
    \adc_out_1[18] ,
    \adc_out_1[17] ,
    \adc_out_1[16] ,
    \adc_out_1[15] ,
    \adc_out_1[14] ,
    \adc_out_1[13] ,
    \adc_out_1[12] ,
    \adc_out_1[11] ,
    \adc_out_1[10] ,
    \adc_out_1[9] ,
    \adc_out_1[8] ,
    \adc_out_1[7] ,
    \adc_out_1[6] ,
    \adc_out_1[5] ,
    \adc_out_1[4] ,
    \adc_out_1[3] ,
    \adc_out_1[2] ,
    \adc_out_1[1] ,
    \adc_out_1[0] }),
    .adc2_dat_i({\adc_out_2[31] ,
    \adc_out_2[30] ,
    \adc_out_2[29] ,
    \adc_out_2[28] ,
    \adc_out_2[27] ,
    \adc_out_2[26] ,
    \adc_out_2[25] ,
    \adc_out_2[24] ,
    \adc_out_2[23] ,
    \adc_out_2[22] ,
    \adc_out_2[21] ,
    \adc_out_2[20] ,
    \adc_out_2[19] ,
    \adc_out_2[18] ,
    \adc_out_2[17] ,
    \adc_out_2[16] ,
    \adc_out_2[15] ,
    \adc_out_2[14] ,
    \adc_out_2[13] ,
    \adc_out_2[12] ,
    \adc_out_2[11] ,
    \adc_out_2[10] ,
    \adc_out_2[9] ,
    \adc_out_2[8] ,
    \adc_out_2[7] ,
    \adc_out_2[6] ,
    \adc_out_2[5] ,
    \adc_out_2[4] ,
    \adc_out_2[3] ,
    \adc_out_2[2] ,
    \adc_out_2[1] ,
    \adc_out_2[0] }),
    .adc_dvalid_i({\sinc3_dvalid[2] ,
    \sinc3_dvalid[1] ,
    \sinc3_dvalid[0] }),
    .io_in({io_in[37],
    io_in[36],
    io_in[35],
    io_in[34],
    io_in[33],
    io_in[32],
    io_in[31],
    io_in[30],
    io_in[29],
    io_in[28],
    io_in[27],
    io_in[26],
    io_in[25],
    io_in[24],
    io_in[23],
    io_in[22],
    io_in[21],
    io_in[20],
    io_in[19],
    io_in[18],
    io_in[17],
    io_in[16],
    io_in[15],
    io_in[14],
    io_in[13],
    io_in[12],
    io_in[11],
    io_in[10],
    io_in[9],
    io_in[8],
    io_in[7],
    io_in[6],
    io_in[5],
    io_in[4],
    io_in[3],
    io_in[2],
    io_in[1],
    io_in[0]}),
    .io_oeb({io_oeb[37],
    io_oeb[36],
    io_oeb[35],
    io_oeb[34],
    io_oeb[33],
    io_oeb[32],
    io_oeb[31],
    io_oeb[30],
    io_oeb[29],
    io_oeb[28],
    io_oeb[27],
    io_oeb[26],
    io_oeb[25],
    io_oeb[24],
    io_oeb[23],
    io_oeb[22],
    io_oeb[21],
    io_oeb[20],
    io_oeb[19],
    io_oeb[18],
    io_oeb[17],
    io_oeb[16],
    io_oeb[15],
    io_oeb[14],
    io_oeb[13],
    io_oeb[12],
    io_oeb[11],
    io_oeb[10],
    io_oeb[9],
    io_oeb[8],
    io_oeb[7],
    io_oeb[6],
    io_oeb[5],
    io_oeb[4],
    io_oeb[3],
    io_oeb[2],
    io_oeb[1],
    io_oeb[0]}),
    .io_out({io_out[37],
    io_out[36],
    io_out[35],
    io_out[34],
    io_out[33],
    io_out[32],
    io_out[31],
    io_out[30],
    io_out[29],
    io_out[28],
    io_out[27],
    io_out[26],
    io_out[25],
    io_out[24],
    io_out[23],
    io_out[22],
    io_out[21],
    io_out[20],
    io_out[19],
    io_out[18],
    io_out[17],
    io_out[16],
    io_out[15],
    io_out[14],
    io_out[13],
    io_out[12],
    io_out[11],
    io_out[10],
    io_out[9],
    io_out[8],
    io_out[7],
    io_out[6],
    io_out[5],
    io_out[4],
    io_out[3],
    io_out[2],
    io_out[1],
    io_out[0]}),
    .irq({user_irq[2],
    user_irq[1],
    user_irq[0]}),
    .mem1_data_i({\m2w_data1[31] ,
    \m2w_data1[30] ,
    \m2w_data1[29] ,
    \m2w_data1[28] ,
    \m2w_data1[27] ,
    \m2w_data1[26] ,
    \m2w_data1[25] ,
    \m2w_data1[24] ,
    \m2w_data1[23] ,
    \m2w_data1[22] ,
    \m2w_data1[21] ,
    \m2w_data1[20] ,
    \m2w_data1[19] ,
    \m2w_data1[18] ,
    \m2w_data1[17] ,
    \m2w_data1[16] ,
    \m2w_data1[15] ,
    \m2w_data1[14] ,
    \m2w_data1[13] ,
    \m2w_data1[12] ,
    \m2w_data1[11] ,
    \m2w_data1[10] ,
    \m2w_data1[9] ,
    \m2w_data1[8] ,
    \m2w_data1[7] ,
    \m2w_data1[6] ,
    \m2w_data1[5] ,
    \m2w_data1[4] ,
    \m2w_data1[3] ,
    \m2w_data1[2] ,
    \m2w_data1[1] ,
    \m2w_data1[0] }),
    .mem_data_i({\m2w_data0[31] ,
    \m2w_data0[30] ,
    \m2w_data0[29] ,
    \m2w_data0[28] ,
    \m2w_data0[27] ,
    \m2w_data0[26] ,
    \m2w_data0[25] ,
    \m2w_data0[24] ,
    \m2w_data0[23] ,
    \m2w_data0[22] ,
    \m2w_data0[21] ,
    \m2w_data0[20] ,
    \m2w_data0[19] ,
    \m2w_data0[18] ,
    \m2w_data0[17] ,
    \m2w_data0[16] ,
    \m2w_data0[15] ,
    \m2w_data0[14] ,
    \m2w_data0[13] ,
    \m2w_data0[12] ,
    \m2w_data0[11] ,
    \m2w_data0[10] ,
    \m2w_data0[9] ,
    \m2w_data0[8] ,
    \m2w_data0[7] ,
    \m2w_data0[6] ,
    \m2w_data0[5] ,
    \m2w_data0[4] ,
    \m2w_data0[3] ,
    \m2w_data0[2] ,
    \m2w_data0[1] ,
    \m2w_data0[0] }),
    .mem_data_o({\w2m_data[31] ,
    \w2m_data[30] ,
    \w2m_data[29] ,
    \w2m_data[28] ,
    \w2m_data[27] ,
    \w2m_data[26] ,
    \w2m_data[25] ,
    \w2m_data[24] ,
    \w2m_data[23] ,
    \w2m_data[22] ,
    \w2m_data[21] ,
    \w2m_data[20] ,
    \w2m_data[19] ,
    \w2m_data[18] ,
    \w2m_data[17] ,
    \w2m_data[16] ,
    \w2m_data[15] ,
    \w2m_data[14] ,
    \w2m_data[13] ,
    \w2m_data[12] ,
    \w2m_data[11] ,
    \w2m_data[10] ,
    \w2m_data[9] ,
    \w2m_data[8] ,
    \w2m_data[7] ,
    \w2m_data[6] ,
    \w2m_data[5] ,
    \w2m_data[4] ,
    \w2m_data[3] ,
    \w2m_data[2] ,
    \w2m_data[1] ,
    \w2m_data[0] }),
    .mem_raddr_o({\raddr[8] ,
    \raddr[7] ,
    \raddr[6] ,
    \raddr[5] ,
    \raddr[4] ,
    \raddr[3] ,
    \raddr[2] ,
    \raddr[1] ,
    \raddr[0] }),
    .mem_renb_o({\renb[1] ,
    \renb[0] }),
    .mem_waddr_o({\waddr[8] ,
    \waddr[7] ,
    \waddr[6] ,
    \waddr[5] ,
    \waddr[4] ,
    \waddr[3] ,
    \waddr[2] ,
    \waddr[1] ,
    \waddr[0] }),
    .mem_wenb_o({\wenb[1] ,
    \wenb[0] }),
    .oversample_o({\oversample[9] ,
    \oversample[8] ,
    \oversample[7] ,
    \oversample[6] ,
    \oversample[5] ,
    \oversample[4] ,
    \oversample[3] ,
    \oversample[2] ,
    \oversample[1] ,
    \oversample[0] }),
    .sinc3_en_o({\en[2] ,
    \en[1] ,
    \en[0] }),
    .vco_enb_o({\vco_enb[2] ,
    \vco_enb[1] ,
    \vco_enb[0] }),
    .wbs_adr_i({wbs_adr_i[31],
    wbs_adr_i[30],
    wbs_adr_i[29],
    wbs_adr_i[28],
    wbs_adr_i[27],
    wbs_adr_i[26],
    wbs_adr_i[25],
    wbs_adr_i[24],
    wbs_adr_i[23],
    wbs_adr_i[22],
    wbs_adr_i[21],
    wbs_adr_i[20],
    wbs_adr_i[19],
    wbs_adr_i[18],
    wbs_adr_i[17],
    wbs_adr_i[16],
    wbs_adr_i[15],
    wbs_adr_i[14],
    wbs_adr_i[13],
    wbs_adr_i[12],
    wbs_adr_i[11],
    wbs_adr_i[10],
    wbs_adr_i[9],
    wbs_adr_i[8],
    wbs_adr_i[7],
    wbs_adr_i[6],
    wbs_adr_i[5],
    wbs_adr_i[4],
    wbs_adr_i[3],
    wbs_adr_i[2],
    wbs_adr_i[1],
    wbs_adr_i[0]}),
    .wbs_dat_i({wbs_dat_i[31],
    wbs_dat_i[30],
    wbs_dat_i[29],
    wbs_dat_i[28],
    wbs_dat_i[27],
    wbs_dat_i[26],
    wbs_dat_i[25],
    wbs_dat_i[24],
    wbs_dat_i[23],
    wbs_dat_i[22],
    wbs_dat_i[21],
    wbs_dat_i[20],
    wbs_dat_i[19],
    wbs_dat_i[18],
    wbs_dat_i[17],
    wbs_dat_i[16],
    wbs_dat_i[15],
    wbs_dat_i[14],
    wbs_dat_i[13],
    wbs_dat_i[12],
    wbs_dat_i[11],
    wbs_dat_i[10],
    wbs_dat_i[9],
    wbs_dat_i[8],
    wbs_dat_i[7],
    wbs_dat_i[6],
    wbs_dat_i[5],
    wbs_dat_i[4],
    wbs_dat_i[3],
    wbs_dat_i[2],
    wbs_dat_i[1],
    wbs_dat_i[0]}),
    .wbs_dat_o({wbs_dat_o[31],
    wbs_dat_o[30],
    wbs_dat_o[29],
    wbs_dat_o[28],
    wbs_dat_o[27],
    wbs_dat_o[26],
    wbs_dat_o[25],
    wbs_dat_o[24],
    wbs_dat_o[23],
    wbs_dat_o[22],
    wbs_dat_o[21],
    wbs_dat_o[20],
    wbs_dat_o[19],
    wbs_dat_o[18],
    wbs_dat_o[17],
    wbs_dat_o[16],
    wbs_dat_o[15],
    wbs_dat_o[14],
    wbs_dat_o[13],
    wbs_dat_o[12],
    wbs_dat_o[11],
    wbs_dat_o[10],
    wbs_dat_o[9],
    wbs_dat_o[8],
    wbs_dat_o[7],
    wbs_dat_o[6],
    wbs_dat_o[5],
    wbs_dat_o[4],
    wbs_dat_o[3],
    wbs_dat_o[2],
    wbs_dat_o[1],
    wbs_dat_o[0]}),
    .wbs_sel_i({wbs_sel_i[3],
    wbs_sel_i[2],
    wbs_sel_i[1],
    wbs_sel_i[0]}),
    .wmask_o({\wmask[3] ,
    \wmask[2] ,
    \wmask[1] ,
    \wmask[0] }));
endmodule
