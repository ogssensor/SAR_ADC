* NGSPICE file created from vco_adc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s50_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s50_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

.subckt vco_adc clk data_out[0] data_out[10] data_out[11] data_out[12] data_out[13]
+ data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[1]
+ data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26]
+ data_out[27] data_out[28] data_out[29] data_out[2] data_out[30] data_out[31] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] data_valid_out
+ enable_in oversample_in[0] oversample_in[1] oversample_in[2] oversample_in[3] oversample_in[4]
+ oversample_in[5] oversample_in[6] oversample_in[7] oversample_in[8] oversample_in[9]
+ phase_in[0] phase_in[10] phase_in[1] phase_in[2] phase_in[3] phase_in[4] phase_in[5]
+ phase_in[6] phase_in[7] phase_in[8] phase_in[9] rst vccd1 vssd1
XFILLER_67_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3155_ _5161_/Q _3672_/B vssd1 vssd1 vccd1 vccd1 _3158_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3086_ _3086_/A _3086_/B vssd1 vssd1 vccd1 vccd1 _3087_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3988_ _4019_/B vssd1 vssd1 vccd1 vccd1 _4012_/B sky130_fd_sc_hd__inv_2
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2939_ _5234_/Q vssd1 vssd1 vccd1 vccd1 _3733_/B sky130_fd_sc_hd__inv_2
X_4609_ _4609_/A _4769_/B vssd1 vssd1 vccd1 vccd1 _4610_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4960_ _4964_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 _4960_/Q sky130_fd_sc_hd__dfxtp_1
X_3911_ _5081_/Q vssd1 vssd1 vccd1 vccd1 _4339_/A sky130_fd_sc_hd__inv_2
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4891_ _4891_/A _4891_/B vssd1 vssd1 vccd1 vccd1 _4894_/B sky130_fd_sc_hd__nor2_1
XFILLER_44_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3842_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4501_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3773_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3784_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2724_ _2854_/B _2724_/B vssd1 vssd1 vccd1 vccd1 _2869_/C sky130_fd_sc_hd__nand2_1
X_2655_ _5262_/Q _4574_/A vssd1 vssd1 vccd1 vccd1 _2957_/B sky130_fd_sc_hd__or2_1
X_4325_ _4427_/A _4427_/B _4324_/Y vssd1 vssd1 vccd1 vccd1 _4406_/B sky130_fd_sc_hd__a21oi_2
X_2586_ _4996_/Q vssd1 vssd1 vccd1 vccd1 _2667_/A sky130_fd_sc_hd__inv_2
XFILLER_59_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _4517_/A _4520_/B _4524_/B vssd1 vssd1 vccd1 vccd1 _4507_/A sky130_fd_sc_hd__nand3_1
XFILLER_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4187_ _4185_/Y _4178_/B _4535_/A vssd1 vssd1 vccd1 vccd1 _4187_/Y sky130_fd_sc_hd__a21oi_1
X_3207_ _3208_/A _3208_/B _3208_/C vssd1 vssd1 vccd1 vccd1 _3207_/X sky130_fd_sc_hd__a21o_1
XFILLER_67_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3138_ _3138_/A vssd1 vssd1 vccd1 vccd1 _3138_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3069_ _5137_/Q _3736_/B vssd1 vssd1 vccd1 vccd1 _3071_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4110_ _4110_/A _4110_/B vssd1 vssd1 vccd1 vccd1 _4115_/A sky130_fd_sc_hd__nand2_1
X_5090_ _5090_/CLK _5090_/D vssd1 vssd1 vccd1 vccd1 _5090_/Q sky130_fd_sc_hd__dfxtp_1
X_4041_ _4142_/B _5066_/Q _5063_/Q vssd1 vssd1 vccd1 vccd1 _4126_/A sky130_fd_sc_hd__and3_1
XFILLER_68_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4943_ _4934_/X _4933_/A _4951_/S vssd1 vssd1 vccd1 vccd1 _4943_/X sky130_fd_sc_hd__mux2_1
XFILLER_32_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4874_ _5094_/Q _3887_/Y _5089_/Q _3891_/Y vssd1 vssd1 vccd1 vccd1 _4874_/X sky130_fd_sc_hd__o22a_1
X_3825_ _5104_/Q _3819_/X _3816_/X _3824_/Y vssd1 vssd1 vccd1 vccd1 _5104_/D sky130_fd_sc_hd__o211a_1
X_3756_ _3758_/A _3756_/B vssd1 vssd1 vccd1 vccd1 _3756_/Y sky130_fd_sc_hd__nand2_1
X_2707_ _5272_/Q vssd1 vssd1 vccd1 vccd1 _2708_/A sky130_fd_sc_hd__inv_2
X_3687_ _5156_/Q _3685_/X _3682_/X _3686_/Y vssd1 vssd1 vccd1 vccd1 _5156_/D sky130_fd_sc_hd__o211a_1
X_2638_ _5275_/Q _4628_/A vssd1 vssd1 vccd1 vccd1 _2716_/A sky130_fd_sc_hd__nor2_1
X_2569_ _5000_/Q vssd1 vssd1 vccd1 vccd1 _4598_/A sky130_fd_sc_hd__inv_2
XFILLER_87_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5288_ _5288_/CLK _5288_/D vssd1 vssd1 vccd1 vccd1 _5288_/Q sky130_fd_sc_hd__dfxtp_1
X_4308_ _5040_/Q vssd1 vssd1 vccd1 vccd1 _4628_/B sky130_fd_sc_hd__inv_2
X_4239_ _5030_/Q vssd1 vssd1 vccd1 vccd1 _4569_/B sky130_fd_sc_hd__inv_2
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3610_ _5173_/Q _3580_/X _3608_/Y _3609_/X _3587_/X vssd1 vssd1 vccd1 vccd1 _5173_/D
+ sky130_fd_sc_hd__o221a_1
X_4590_ _4590_/A _4800_/C vssd1 vssd1 vccd1 vccd1 _4796_/A sky130_fd_sc_hd__and2_1
X_3541_ _3541_/A _3541_/B vssd1 vssd1 vccd1 vccd1 _3576_/A sky130_fd_sc_hd__and2_1
X_3472_ _3476_/A _3472_/B vssd1 vssd1 vccd1 vccd1 _3472_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5211_ _5215_/CLK _5211_/D vssd1 vssd1 vccd1 vccd1 _5211_/Q sky130_fd_sc_hd__dfxtp_1
X_5142_ _5254_/CLK _5142_/D vssd1 vssd1 vccd1 vccd1 _5142_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5073_ _5074_/CLK _5073_/D vssd1 vssd1 vccd1 vccd1 _5073_/Q sky130_fd_sc_hd__dfxtp_1
X_4024_ _4021_/Y _4016_/A _5056_/Q _4023_/Y vssd1 vssd1 vccd1 vccd1 _4185_/B sky130_fd_sc_hd__o211ai_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4926_ _4931_/B _4928_/C vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__and2_1
X_4857_ _4873_/A input8/X vssd1 vssd1 vccd1 vccd1 _4858_/A sky130_fd_sc_hd__or2_1
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3808_ _3810_/A _3808_/B vssd1 vssd1 vccd1 vccd1 _3808_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4788_ _4788_/A _4788_/B vssd1 vssd1 vccd1 vccd1 _4793_/B sky130_fd_sc_hd__or2_1
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3739_ _3792_/A vssd1 vssd1 vccd1 vccd1 _3739_/X sky130_fd_sc_hd__buf_2
XFILLER_69_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2972_ _3230_/B vssd1 vssd1 vccd1 vccd1 _2972_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_34_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4711_ _4711_/A vssd1 vssd1 vccd1 vccd1 _4711_/X sky130_fd_sc_hd__clkbuf_2
X_4642_ _4731_/A _4734_/A vssd1 vssd1 vccd1 vccd1 _4643_/B sky130_fd_sc_hd__nand2_1
X_4573_ _4573_/A _4573_/B vssd1 vssd1 vccd1 vccd1 _4810_/B sky130_fd_sc_hd__nor2_1
X_3524_ _3528_/A _3354_/Y _3355_/B _2850_/X vssd1 vssd1 vccd1 vccd1 _3524_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_89_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3455_ _5214_/Q vssd1 vssd1 vccd1 vccd1 _3787_/B sky130_fd_sc_hd__inv_2
X_3386_ _5198_/Q vssd1 vssd1 vccd1 vccd1 _3830_/B sky130_fd_sc_hd__inv_2
XFILLER_57_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5125_ _5195_/CLK _5125_/D vssd1 vssd1 vccd1 vccd1 _5125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5056_ _5058_/CLK _5056_/D vssd1 vssd1 vccd1 vccd1 _5056_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4007_ _4007_/A _4020_/B _4018_/A vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__nand3_1
XFILLER_72_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4909_ _4909_/A _4913_/B vssd1 vssd1 vccd1 vccd1 _4910_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _3240_/A _3240_/B vssd1 vssd1 vccd1 vccd1 _3248_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3171_ _3148_/Y _3151_/Y _3170_/Y vssd1 vssd1 vccd1 vccd1 _3171_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2955_ _2955_/A _2955_/B vssd1 vssd1 vccd1 vccd1 _2957_/C sky130_fd_sc_hd__nor2_1
X_2886_ _3505_/A _5244_/Q vssd1 vssd1 vccd1 vccd1 _2886_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4625_ _5009_/Q _5041_/Q vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__xor2_1
X_4556_ _4764_/A _4556_/B vssd1 vssd1 vccd1 vccd1 _4619_/B sky130_fd_sc_hd__nor2_1
X_3507_ _3507_/A _3507_/B vssd1 vssd1 vccd1 vccd1 _3508_/A sky130_fd_sc_hd__or2_1
X_4487_ _4487_/A _4487_/B vssd1 vssd1 vccd1 vccd1 _4487_/Y sky130_fd_sc_hd__nor2_1
X_3438_ _3594_/A _3594_/B _3437_/X vssd1 vssd1 vccd1 vccd1 _3581_/B sky130_fd_sc_hd__a21oi_1
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _3571_/A _3449_/A vssd1 vssd1 vccd1 vccd1 _3369_/Y sky130_fd_sc_hd__nor2_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5108_ _5209_/CLK _5108_/D vssd1 vssd1 vccd1 vccd1 _5108_/Q sky130_fd_sc_hd__dfxtp_1
X_5039_ _5051_/CLK _5039_/D vssd1 vssd1 vccd1 vccd1 _5039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput31 _5178_/Q vssd1 vssd1 vccd1 vccd1 data_out[16] sky130_fd_sc_hd__buf_2
Xoutput42 _5188_/Q vssd1 vssd1 vccd1 vccd1 data_out[26] sky130_fd_sc_hd__buf_2
Xoutput53 _5169_/Q vssd1 vssd1 vccd1 vccd1 data_out[7] sky130_fd_sc_hd__buf_2
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2740_ _2729_/A _2857_/B _2736_/Y _2739_/Y vssd1 vssd1 vccd1 vccd1 _2824_/B sky130_fd_sc_hd__o211a_1
X_2671_ _2770_/A _2671_/B vssd1 vssd1 vccd1 vccd1 _2768_/A sky130_fd_sc_hd__nand2_1
X_4410_ _4410_/A _4410_/B vssd1 vssd1 vccd1 vccd1 _4427_/C sky130_fd_sc_hd__nand2_1
X_4341_ _5082_/Q _5050_/Q vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__nor2_1
X_4272_ _4272_/A _4598_/B vssd1 vssd1 vccd1 vccd1 _4273_/B sky130_fd_sc_hd__nor2_1
X_3223_ _3229_/B _3229_/A vssd1 vssd1 vccd1 vccd1 _3230_/A sky130_fd_sc_hd__or2_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3154_ _5257_/Q vssd1 vssd1 vccd1 vccd1 _3672_/B sky130_fd_sc_hd__inv_2
XFILLER_82_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3085_ _3726_/B _5141_/Q vssd1 vssd1 vccd1 vccd1 _3086_/B sky130_fd_sc_hd__and2_1
XFILLER_82_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3987_ _3987_/A _3987_/B vssd1 vssd1 vccd1 vccd1 _4019_/B sky130_fd_sc_hd__or2_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2938_ _2938_/A _2938_/B vssd1 vssd1 vccd1 vccd1 _2938_/X sky130_fd_sc_hd__xor2_2
X_2869_ _2869_/A _2869_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__and3_1
X_4608_ _5003_/Q _5035_/Q vssd1 vssd1 vccd1 vccd1 _4769_/B sky130_fd_sc_hd__nand2_1
X_4539_ _5013_/Q _5045_/Q vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__nor2_1
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_41_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3910_ _5082_/Q vssd1 vssd1 vccd1 vccd1 _4343_/A sky130_fd_sc_hd__inv_2
X_4890_ _4890_/A _4890_/B vssd1 vssd1 vccd1 vccd1 _4891_/B sky130_fd_sc_hd__nor2_1
X_3841_ _4841_/A vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3772_ _5124_/Q _3766_/X _3763_/X _3771_/Y vssd1 vssd1 vccd1 vccd1 _5124_/D sky130_fd_sc_hd__o211a_1
X_2723_ _4735_/A _5278_/Q vssd1 vssd1 vccd1 vccd1 _2724_/B sky130_fd_sc_hd__nand2_1
X_2654_ _2922_/B vssd1 vssd1 vccd1 vccd1 _2654_/Y sky130_fd_sc_hd__inv_2
X_2585_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__clkbuf_2
X_4324_ _4324_/A _4324_/B vssd1 vssd1 vccd1 vccd1 _4324_/Y sky130_fd_sc_hd__nand2_1
X_4255_ _5057_/Q _5025_/Q vssd1 vssd1 vccd1 vccd1 _4524_/B sky130_fd_sc_hd__nand2_1
X_4186_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4535_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_67_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3206_ _3206_/A _3206_/B vssd1 vssd1 vccd1 vccd1 _3208_/C sky130_fd_sc_hd__nor2_1
X_3137_ _3118_/A _3136_/Y _3118_/B vssd1 vssd1 vccd1 vccd1 _3138_/A sky130_fd_sc_hd__o21ba_1
XFILLER_82_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3068_ _5233_/Q vssd1 vssd1 vccd1 vccd1 _3736_/B sky130_fd_sc_hd__inv_2
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4040_ _4278_/A _4272_/A vssd1 vssd1 vccd1 vccd1 _4142_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4942_ _4937_/X _4936_/A _4951_/S vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__mux2_1
X_4873_ _4873_/A _4873_/B vssd1 vssd1 vccd1 vccd1 _4975_/D sky130_fd_sc_hd__nor2_1
X_3824_ _3824_/A _3824_/B vssd1 vssd1 vccd1 vccd1 _3824_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3755_ _5131_/Q _3753_/X _3750_/X _3754_/Y vssd1 vssd1 vccd1 vccd1 _5131_/D sky130_fd_sc_hd__o211a_1
X_3686_ _3690_/A _3686_/B vssd1 vssd1 vccd1 vccd1 _3686_/Y sky130_fd_sc_hd__nand2_1
X_2706_ _2704_/Y _2706_/B vssd1 vssd1 vccd1 vccd1 _2901_/A sky130_fd_sc_hd__and2b_1
X_2637_ _2880_/B _2880_/C _2877_/B vssd1 vssd1 vccd1 vccd1 _2643_/A sky130_fd_sc_hd__and3_1
XFILLER_58_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2568_ _5268_/Q _2564_/X _2565_/X _2567_/Y vssd1 vssd1 vccd1 vccd1 _5268_/D sky130_fd_sc_hd__o211a_1
X_4307_ _5072_/Q _5040_/Q vssd1 vssd1 vccd1 vccd1 _4445_/A sky130_fd_sc_hd__nor2_1
X_2499_ _5018_/Q vssd1 vssd1 vccd1 vccd1 _4702_/A sky130_fd_sc_hd__clkinv_2
X_5287_ _5287_/CLK _5287_/D vssd1 vssd1 vccd1 vccd1 _5287_/Q sky130_fd_sc_hd__dfxtp_1
X_4238_ _5061_/Q _5029_/Q vssd1 vssd1 vccd1 vccd1 _4497_/C sky130_fd_sc_hd__nand2_1
XFILLER_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ _4169_/A _4169_/B _4179_/A _4169_/D vssd1 vssd1 vccd1 vccd1 _4169_/X sky130_fd_sc_hd__and4_1
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _5186_/Q _3537_/X _3303_/X _3539_/Y vssd1 vssd1 vccd1 vccd1 _5186_/D sky130_fd_sc_hd__o211a_1
XFILLER_6_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5210_ _5215_/CLK _5210_/D vssd1 vssd1 vccd1 vccd1 _5210_/Q sky130_fd_sc_hd__dfxtp_1
X_3471_ _3784_/B _5119_/Q vssd1 vssd1 vccd1 vccd1 _3472_/B sky130_fd_sc_hd__and2_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5141_ _5251_/CLK _5141_/D vssd1 vssd1 vccd1 vccd1 _5141_/Q sky130_fd_sc_hd__dfxtp_1
X_5072_ _5074_/CLK _5072_/D vssd1 vssd1 vccd1 vccd1 _5072_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4023_ _4023_/A _4192_/B vssd1 vssd1 vccd1 vccd1 _4023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_37_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4925_ _4925_/A _4925_/B vssd1 vssd1 vccd1 vccd1 _4928_/C sky130_fd_sc_hd__nand2_1
X_4856_ _4856_/A vssd1 vssd1 vccd1 vccd1 _4984_/D sky130_fd_sc_hd__clkbuf_1
X_3807_ _5111_/Q _3805_/X _3802_/X _3806_/Y vssd1 vssd1 vccd1 vccd1 _5111_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4787_ _5001_/Q _4987_/Q _4784_/X _4786_/X vssd1 vssd1 vccd1 vccd1 _5001_/D sky130_fd_sc_hd__o211a_1
X_3738_ _3738_/A vssd1 vssd1 vccd1 vccd1 _3792_/A sky130_fd_sc_hd__buf_2
XFILLER_69_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3669_ _5162_/Q _3634_/X _3667_/Y _3668_/Y _3642_/X vssd1 vssd1 vccd1 vccd1 _5162_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2971_ _5229_/Q _2907_/X _2969_/Y _2970_/X _2914_/X vssd1 vssd1 vccd1 vccd1 _5229_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_61_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4710_ _4710_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4710_/Y sky130_fd_sc_hd__nor2_1
X_4641_ _4641_/A _4641_/B vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__nor2_1
X_4572_ _4811_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4573_/B sky130_fd_sc_hd__nor2_1
X_3523_ _3528_/A _3355_/B _3354_/Y vssd1 vssd1 vccd1 vccd1 _3523_/X sky130_fd_sc_hd__a21o_1
XFILLER_6_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3454_ _3541_/A _3541_/B _3453_/X vssd1 vssd1 vccd1 vccd1 _3454_/Y sky130_fd_sc_hd__a21oi_1
X_3385_ _5199_/Q vssd1 vssd1 vccd1 vccd1 _3827_/B sky130_fd_sc_hd__inv_2
XFILLER_69_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5124_ _5193_/CLK _5124_/D vssd1 vssd1 vccd1 vccd1 _5124_/Q sky130_fd_sc_hd__dfxtp_1
X_5055_ _5058_/CLK _5055_/D vssd1 vssd1 vccd1 vccd1 _5055_/Q sky130_fd_sc_hd__dfxtp_2
X_4006_ _4009_/C _4005_/A _4004_/A _4004_/B vssd1 vssd1 vccd1 vccd1 _4018_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_72_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4908_ _4912_/B vssd1 vssd1 vccd1 vccd1 _4913_/B sky130_fd_sc_hd__inv_2
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4839_ _4839_/A _4990_/Q vssd1 vssd1 vccd1 vccd1 _4839_/X sky130_fd_sc_hd__and2_1
XFILLER_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold20 hold20/A vssd1 vssd1 vccd1 vccd1 hold20/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_48_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ _3170_/A _3170_/B vssd1 vssd1 vccd1 vccd1 _3170_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2954_ _5263_/Q _4811_/A vssd1 vssd1 vccd1 vccd1 _2955_/A sky130_fd_sc_hd__nor2_1
X_2885_ _2877_/Y _2876_/Y _2875_/X _2884_/Y vssd1 vssd1 vccd1 vccd1 _2885_/X sky130_fd_sc_hd__a31o_1
X_4624_ _4637_/C _4624_/B vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__nor2_1
X_4555_ _5006_/Q _5038_/Q vssd1 vssd1 vccd1 vccd1 _4617_/A sky130_fd_sc_hd__nor2_1
X_3506_ _3504_/Y _3505_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5192_/D sky130_fd_sc_hd__a21oi_1
X_4486_ _4486_/A _4486_/B vssd1 vssd1 vccd1 vccd1 _4487_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3437_ _3593_/A _3593_/B _3602_/B vssd1 vssd1 vccd1 vccd1 _3437_/X sky130_fd_sc_hd__or3_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _5114_/Q _3797_/B vssd1 vssd1 vccd1 vccd1 _3449_/A sky130_fd_sc_hd__nor2_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5107_ _5206_/CLK _5107_/D vssd1 vssd1 vccd1 vccd1 _5107_/Q sky130_fd_sc_hd__dfxtp_1
X_3299_ _3299_/A _3299_/B vssd1 vssd1 vccd1 vccd1 _3300_/A sky130_fd_sc_hd__nand2_1
X_5038_ _5272_/CLK _5038_/D vssd1 vssd1 vccd1 vccd1 _5038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput32 _5179_/Q vssd1 vssd1 vccd1 vccd1 data_out[17] sky130_fd_sc_hd__buf_2
Xoutput43 _5189_/Q vssd1 vssd1 vccd1 vccd1 data_out[27] sky130_fd_sc_hd__buf_2
Xoutput54 _5170_/Q vssd1 vssd1 vccd1 vccd1 data_out[8] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2670_ _4589_/A _5264_/Q vssd1 vssd1 vccd1 vccd1 _2671_/B sky130_fd_sc_hd__nand2_1
X_4340_ _4340_/A _4340_/B vssd1 vssd1 vccd1 vccd1 _4396_/B sky130_fd_sc_hd__nand2_1
X_4271_ _5032_/Q vssd1 vssd1 vccd1 vccd1 _4598_/B sky130_fd_sc_hd__inv_2
X_3222_ _3113_/C _3236_/B _3031_/X vssd1 vssd1 vccd1 vccd1 _3229_/A sky130_fd_sc_hd__o21ba_1
X_3153_ _3165_/B _3165_/A _3170_/A _3152_/Y vssd1 vssd1 vccd1 vccd1 _3167_/B sky130_fd_sc_hd__o22ai_2
XFILLER_82_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3084_ _5141_/Q _3726_/B vssd1 vssd1 vccd1 vccd1 _3086_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3986_ _3986_/A _3986_/B _3986_/C vssd1 vssd1 vccd1 vccd1 _4019_/A sky130_fd_sc_hd__nand3_1
X_2937_ _5235_/Q _2907_/X _2935_/Y _2936_/X _2914_/X vssd1 vssd1 vccd1 vccd1 _5235_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2868_ _5247_/Q _2814_/X _2865_/Y _2867_/X _2822_/X vssd1 vssd1 vccd1 vccd1 _5247_/D
+ sky130_fd_sc_hd__o221a_1
X_4607_ _4607_/A _4607_/B vssd1 vssd1 vccd1 vccd1 _4609_/A sky130_fd_sc_hd__nand2_1
X_2799_ _2809_/A vssd1 vssd1 vccd1 vccd1 _3505_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4538_ hold24/A _4538_/B vssd1 vssd1 vccd1 vccd1 _4690_/B sky130_fd_sc_hd__nor2_1
X_4469_ _4784_/A vssd1 vssd1 vccd1 vccd1 _4469_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_77_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3840_ _5098_/Q _3832_/X _3829_/X _3839_/Y vssd1 vssd1 vccd1 vccd1 _5098_/D sky130_fd_sc_hd__o211a_1
X_3771_ _3771_/A _3771_/B vssd1 vssd1 vccd1 vccd1 _3771_/Y sky130_fd_sc_hd__nand2_1
X_2722_ _2722_/A vssd1 vssd1 vccd1 vccd1 _2854_/B sky130_fd_sc_hd__inv_2
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2653_ _2683_/B _2681_/A _2652_/Y vssd1 vssd1 vccd1 vccd1 _2922_/B sky130_fd_sc_hd__o21a_1
X_2584_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2584_/X sky130_fd_sc_hd__clkbuf_2
X_4323_ _4423_/B _4410_/A _4410_/B vssd1 vssd1 vccd1 vccd1 _4324_/B sky130_fd_sc_hd__and3_1
X_4254_ _5058_/Q _5026_/Q vssd1 vssd1 vccd1 vccd1 _4520_/B sky130_fd_sc_hd__nand2_1
X_4185_ _4185_/A _4185_/B vssd1 vssd1 vccd1 vccd1 _4185_/Y sky130_fd_sc_hd__nand2_1
X_3205_ _3212_/B _3212_/A vssd1 vssd1 vccd1 vccd1 _3208_/A sky130_fd_sc_hd__or2_1
X_3136_ _5150_/Q _3701_/B vssd1 vssd1 vccd1 vccd1 _3136_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3067_ _3287_/B _3067_/B vssd1 vssd1 vccd1 vccd1 _3292_/B sky130_fd_sc_hd__nand2_1
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3969_ _3967_/A _3967_/B _3994_/A _3975_/A vssd1 vssd1 vccd1 vccd1 _3969_/X sky130_fd_sc_hd__o211a_1
XFILLER_88_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4941_ _5289_/Q _3832_/X _4784_/X _4940_/Y vssd1 vssd1 vccd1 vccd1 _5289_/D sky130_fd_sc_hd__o211a_1
X_4872_ _4872_/A _4987_/Q vssd1 vssd1 vccd1 vccd1 _4873_/B sky130_fd_sc_hd__nand2_1
X_3823_ _5105_/Q _3819_/X _3816_/X _3822_/Y vssd1 vssd1 vccd1 vccd1 _5105_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3754_ _3758_/A _3754_/B vssd1 vssd1 vccd1 vccd1 _3754_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3685_ _3725_/A vssd1 vssd1 vccd1 vccd1 _3685_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2705_ _4761_/A _5273_/Q vssd1 vssd1 vccd1 vccd1 _2706_/B sky130_fd_sc_hd__nand2_1
X_2636_ _4637_/A _5276_/Q vssd1 vssd1 vccd1 vccd1 _2877_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2567_ _2573_/A _4603_/A vssd1 vssd1 vccd1 vccd1 _2567_/Y sky130_fd_sc_hd__nand2_1
X_4306_ _4440_/A _4430_/A vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__nand2_1
X_5286_ _5287_/CLK _5286_/D vssd1 vssd1 vccd1 vccd1 _5286_/Q sky130_fd_sc_hd__dfxtp_1
X_2498_ _2557_/A vssd1 vssd1 vccd1 vccd1 _2516_/A sky130_fd_sc_hd__clkbuf_2
X_4237_ _5062_/Q _5030_/Q vssd1 vssd1 vccd1 vccd1 _4263_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4168_ _4168_/A vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__inv_2
XFILLER_67_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4099_ _4099_/A _4144_/B vssd1 vssd1 vccd1 vccd1 _4099_/Y sky130_fd_sc_hd__nand2_1
X_3119_ _3119_/A vssd1 vssd1 vccd1 vccd1 _3132_/A sky130_fd_sc_hd__inv_2
XFILLER_43_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3470_ _5119_/Q _3784_/B vssd1 vssd1 vccd1 vccd1 _3476_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5140_ _5207_/CLK _5140_/D vssd1 vssd1 vccd1 vccd1 _5140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5071_ _5074_/CLK _5071_/D vssd1 vssd1 vccd1 vccd1 _5071_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4022_ _4022_/A _4022_/B vssd1 vssd1 vccd1 vccd1 _4023_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4924_ _4930_/B vssd1 vssd1 vccd1 vccd1 _4931_/B sky130_fd_sc_hd__inv_2
X_4855_ _4873_/A input9/X vssd1 vssd1 vccd1 vccd1 _4856_/A sky130_fd_sc_hd__or2_1
XFILLER_20_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3806_ _3810_/A _3806_/B vssd1 vssd1 vccd1 vccd1 _3806_/Y sky130_fd_sc_hd__nand2_1
X_4786_ _4781_/A _4785_/Y _4501_/X vssd1 vssd1 vccd1 vccd1 _4786_/X sky130_fd_sc_hd__a21o_1
X_3737_ _5137_/Q _3725_/X _3735_/X _3736_/Y vssd1 vssd1 vccd1 vccd1 _5137_/D sky130_fd_sc_hd__o211a_1
X_3668_ _3668_/A _3668_/B vssd1 vssd1 vccd1 vccd1 _3668_/Y sky130_fd_sc_hd__nand2_1
X_3599_ _3597_/B _3597_/A _3598_/X vssd1 vssd1 vccd1 vccd1 _3599_/X sky130_fd_sc_hd__a21o_1
X_2619_ _4656_/A _5284_/Q vssd1 vssd1 vccd1 vccd1 _2620_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5269_ _5288_/CLK _5269_/D vssd1 vssd1 vccd1 vccd1 _5269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2970_ _2969_/B _2969_/A _2912_/X vssd1 vssd1 vccd1 vccd1 _2970_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4640_ _5011_/Q _5043_/Q vssd1 vssd1 vccd1 vccd1 _4641_/A sky130_fd_sc_hd__nor2_1
X_4571_ _4996_/Q _5028_/Q vssd1 vssd1 vccd1 vccd1 _4573_/A sky130_fd_sc_hd__nor2_1
X_3522_ _3527_/A _3345_/Y vssd1 vssd1 vccd1 vccd1 _3528_/A sky130_fd_sc_hd__or2b_1
X_3453_ _3453_/A _3566_/B _3453_/C vssd1 vssd1 vccd1 vccd1 _3453_/X sky130_fd_sc_hd__or3_1
X_5123_ _5195_/CLK _5123_/D vssd1 vssd1 vccd1 vccd1 _5123_/Q sky130_fd_sc_hd__dfxtp_1
X_3384_ _3384_/A _3419_/A vssd1 vssd1 vccd1 vccd1 _3605_/A sky130_fd_sc_hd__nand2_1
X_5054_ _5070_/CLK _5054_/D vssd1 vssd1 vccd1 vccd1 _5054_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4005_ _4005_/A _4009_/C _4005_/C vssd1 vssd1 vccd1 vccd1 _4020_/B sky130_fd_sc_hd__nand3_2
XFILLER_65_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4907_ _4907_/A _5092_/Q vssd1 vssd1 vccd1 vccd1 _4912_/B sky130_fd_sc_hd__nand2_1
XFILLER_40_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4838_ _4990_/Q _4839_/A vssd1 vssd1 vccd1 vccd1 _4838_/Y sky130_fd_sc_hd__nor2_1
X_4769_ _4769_/A _4769_/B vssd1 vssd1 vccd1 vccd1 _4770_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold10 hold10/A vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_28_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2953_ _2953_/A vssd1 vssd1 vccd1 vccd1 _2957_/A sky130_fd_sc_hd__inv_2
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2884_ _2884_/A _2978_/A vssd1 vssd1 vccd1 vccd1 _2884_/Y sky130_fd_sc_hd__nand2_1
X_4623_ _4623_/A _4623_/B vssd1 vssd1 vccd1 vccd1 _4624_/B sky130_fd_sc_hd__nor2_1
X_4554_ _4554_/A vssd1 vssd1 vccd1 vccd1 _4716_/A sky130_fd_sc_hd__inv_2
X_3505_ _3505_/A _5192_/Q vssd1 vssd1 vccd1 vccd1 _3505_/Y sky130_fd_sc_hd__nand2_1
X_4485_ _4490_/B _4490_/A vssd1 vssd1 vccd1 vccd1 _4486_/A sky130_fd_sc_hd__or2_1
X_3436_ _3436_/A _3436_/B vssd1 vssd1 vccd1 vccd1 _3602_/B sky130_fd_sc_hd__or2_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3367_ _5115_/Q _3795_/B vssd1 vssd1 vccd1 vccd1 _3571_/A sky130_fd_sc_hd__nor2_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5106_ _5206_/CLK _5106_/D vssd1 vssd1 vccd1 vccd1 _5106_/Q sky130_fd_sc_hd__dfxtp_1
X_5037_ _5272_/CLK _5037_/D vssd1 vssd1 vccd1 vccd1 _5037_/Q sky130_fd_sc_hd__dfxtp_1
X_3298_ _3299_/A _3299_/B _3301_/A _2898_/X vssd1 vssd1 vccd1 vccd1 _3298_/X sky130_fd_sc_hd__a31o_1
XFILLER_72_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput33 _5180_/Q vssd1 vssd1 vccd1 vccd1 data_out[18] sky130_fd_sc_hd__buf_2
Xoutput55 _5171_/Q vssd1 vssd1 vccd1 vccd1 data_out[9] sky130_fd_sc_hd__buf_2
Xoutput44 _5190_/Q vssd1 vssd1 vccd1 vccd1 data_out[28] sky130_fd_sc_hd__buf_2
XFILLER_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4270_ _5064_/Q _5032_/Q vssd1 vssd1 vccd1 vccd1 _4273_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3221_ _3221_/A _3221_/B vssd1 vssd1 vccd1 vccd1 _3236_/B sky130_fd_sc_hd__and2_1
X_3152_ _3676_/B _5159_/Q _3148_/Y _3151_/Y vssd1 vssd1 vccd1 vccd1 _3152_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_39_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3083_ _5237_/Q vssd1 vssd1 vccd1 vccd1 _3726_/B sky130_fd_sc_hd__inv_2
XFILLER_35_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3985_ _3986_/C _3986_/A _3981_/A _3981_/B vssd1 vssd1 vccd1 vccd1 _4020_/C sky130_fd_sc_hd__o2bb2ai_1
XFILLER_22_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2936_ _2935_/B _2935_/A _2912_/X vssd1 vssd1 vccd1 vccd1 _2936_/X sky130_fd_sc_hd__a21o_1
XFILLER_50_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2867_ _2870_/B _2733_/X _2854_/B _2866_/X vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__a31o_1
X_4606_ _4777_/A _4777_/B _4605_/X vssd1 vssd1 vccd1 vccd1 _4767_/B sky130_fd_sc_hd__a21oi_1
XFILLER_7_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2798_ _2798_/A _3504_/C _2798_/C vssd1 vssd1 vccd1 vccd1 _2798_/Y sky130_fd_sc_hd__nand3_1
X_4537_ _4537_/A _4537_/B vssd1 vssd1 vccd1 vccd1 _4674_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4468_ _4987_/Q _5036_/Q _4466_/Y _4467_/X _4438_/X vssd1 vssd1 vccd1 vccd1 _5036_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3419_ _3419_/A _3419_/B vssd1 vssd1 vccd1 vccd1 _3614_/A sky130_fd_sc_hd__nand2_1
X_4399_ _4746_/A _5049_/Q vssd1 vssd1 vccd1 vccd1 _4399_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3770_ _5125_/Q _3766_/X _3763_/X _3769_/Y vssd1 vssd1 vccd1 vccd1 _5125_/D sky130_fd_sc_hd__o211a_1
X_2721_ _5278_/Q _4735_/A vssd1 vssd1 vccd1 vccd1 _2722_/A sky130_fd_sc_hd__nor2_1
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2652_ _2683_/A vssd1 vssd1 vccd1 vccd1 _2652_/Y sky130_fd_sc_hd__inv_2
X_2583_ _5264_/Q _2564_/X _2565_/X _2582_/Y vssd1 vssd1 vccd1 vccd1 _5264_/D sky130_fd_sc_hd__o211a_1
X_4322_ _4322_/A _4548_/B vssd1 vssd1 vccd1 vccd1 _4410_/B sky130_fd_sc_hd__nand2_1
X_4253_ _4529_/B _4523_/B _4524_/A vssd1 vssd1 vccd1 vccd1 _4517_/A sky130_fd_sc_hd__o21ai_1
XFILLER_59_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3204_ _3132_/A _3203_/Y _3138_/Y vssd1 vssd1 vccd1 vccd1 _3212_/A sky130_fd_sc_hd__o21a_1
XFILLER_86_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4184_ _4987_/Q _5057_/Q _4180_/Y _4182_/X _4183_/X vssd1 vssd1 vccd1 vccd1 _5057_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_67_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3135_ _3135_/A _3206_/A vssd1 vssd1 vccd1 vccd1 _3135_/Y sky130_fd_sc_hd__nor2_1
XFILLER_67_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3066_ _3740_/B _5136_/Q vssd1 vssd1 vccd1 vccd1 _3067_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3968_ _3975_/A _3994_/A _3975_/C vssd1 vssd1 vccd1 vccd1 _3968_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2919_ _3826_/A vssd1 vssd1 vccd1 vccd1 _4940_/A sky130_fd_sc_hd__clkbuf_4
X_3899_ _4984_/Q vssd1 vssd1 vccd1 vccd1 _3899_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _4940_/A _4940_/B vssd1 vssd1 vccd1 vccd1 _4940_/Y sky130_fd_sc_hd__nand2_1
X_4871_ _4873_/A _4871_/B vssd1 vssd1 vccd1 vccd1 _4976_/D sky130_fd_sc_hd__nor2_1
X_3822_ _3824_/A _3822_/B vssd1 vssd1 vccd1 vccd1 _3822_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3753_ _3792_/A vssd1 vssd1 vccd1 vccd1 _3753_/X sky130_fd_sc_hd__clkbuf_2
X_3684_ _5157_/Q _3671_/X _3682_/X _3683_/Y vssd1 vssd1 vccd1 vccd1 _5157_/D sky130_fd_sc_hd__o211a_1
X_2704_ _5273_/Q _4761_/A vssd1 vssd1 vccd1 vccd1 _2704_/Y sky130_fd_sc_hd__nor2_1
X_2635_ _2644_/A _2635_/B vssd1 vssd1 vccd1 vccd1 _2880_/B sky130_fd_sc_hd__nor2_1
X_4305_ _4319_/B _4305_/B vssd1 vssd1 vccd1 vccd1 _4430_/A sky130_fd_sc_hd__nor2_1
X_2566_ _5001_/Q vssd1 vssd1 vccd1 vccd1 _4603_/A sky130_fd_sc_hd__inv_2
X_2497_ _5286_/Q _2481_/X _2485_/X _2496_/Y vssd1 vssd1 vccd1 vccd1 _5286_/D sky130_fd_sc_hd__o211a_1
X_5285_ _5287_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _5285_/Q sky130_fd_sc_hd__dfxtp_1
X_4236_ _4476_/A _4478_/C _4476_/B vssd1 vssd1 vccd1 vccd1 _4463_/A sky130_fd_sc_hd__o21bai_1
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4167_ _4167_/A vssd1 vssd1 vccd1 vccd1 _5059_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3118_ _3118_/A _3118_/B vssd1 vssd1 vccd1 vccd1 _3119_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4098_ _4110_/A _5077_/Q _4098_/C vssd1 vssd1 vccd1 vccd1 _4104_/B sky130_fd_sc_hd__nand3_1
XFILLER_55_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3049_ _5228_/Q vssd1 vssd1 vccd1 vccd1 _3751_/B sky130_fd_sc_hd__clkinv_2
XFILLER_43_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5070_ _5070_/CLK _5070_/D vssd1 vssd1 vccd1 vccd1 _5070_/Q sky130_fd_sc_hd__dfxtp_1
X_4021_ _4021_/A _4021_/B vssd1 vssd1 vccd1 vccd1 _4021_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4923_ _4925_/B _4925_/A vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4854_ _4854_/A vssd1 vssd1 vccd1 vccd1 _4985_/D sky130_fd_sc_hd__clkbuf_1
X_3805_ _3832_/A vssd1 vssd1 vccd1 vccd1 _3805_/X sky130_fd_sc_hd__clkbuf_2
X_4785_ _4785_/A _4785_/B vssd1 vssd1 vccd1 vccd1 _4785_/Y sky130_fd_sc_hd__nand2_1
X_3736_ _3744_/A _3736_/B vssd1 vssd1 vccd1 vccd1 _3736_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3667_ _5098_/Q _3839_/B vssd1 vssd1 vccd1 vccd1 _3667_/Y sky130_fd_sc_hd__nor2_1
X_3598_ _3598_/A vssd1 vssd1 vccd1 vccd1 _3598_/X sky130_fd_sc_hd__clkbuf_2
X_2618_ _2622_/B _2828_/C vssd1 vssd1 vccd1 vccd1 _2630_/B sky130_fd_sc_hd__nor2_1
X_2549_ _2555_/A _4761_/A vssd1 vssd1 vccd1 vccd1 _2549_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5268_ _5288_/CLK _5268_/D vssd1 vssd1 vccd1 vccd1 _5268_/Q sky130_fd_sc_hd__dfxtp_1
X_4219_ _4322_/A _4548_/B vssd1 vssd1 vccd1 vccd1 _4421_/A sky130_fd_sc_hd__nor2_1
XFILLER_87_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5199_ _5203_/CLK _5199_/D vssd1 vssd1 vccd1 vccd1 _5199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4570_ _4591_/A _4800_/C _4591_/B vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__o21bai_1
X_3521_ _3483_/B _3532_/B _3350_/X vssd1 vssd1 vccd1 vccd1 _3527_/A sky130_fd_sc_hd__o21ba_1
X_3452_ _3571_/B _3571_/A _3576_/B vssd1 vssd1 vccd1 vccd1 _3453_/C sky130_fd_sc_hd__or3_1
X_3383_ _5107_/Q _3817_/B vssd1 vssd1 vccd1 vccd1 _3419_/A sky130_fd_sc_hd__or2_1
XFILLER_69_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5122_ _5195_/CLK _5122_/D vssd1 vssd1 vccd1 vccd1 _5122_/Q sky130_fd_sc_hd__dfxtp_1
X_5053_ _5070_/CLK _5053_/D vssd1 vssd1 vccd1 vccd1 _5053_/Q sky130_fd_sc_hd__dfxtp_1
X_4004_ _4004_/A _4004_/B vssd1 vssd1 vccd1 vccd1 _4005_/C sky130_fd_sc_hd__nor2_1
XFILLER_80_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4906_ _5092_/Q _4907_/A vssd1 vssd1 vccd1 vccd1 _4909_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4837_ _4846_/A _4840_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4839_/A sky130_fd_sc_hd__or3_1
X_4768_ _4774_/B _4774_/A vssd1 vssd1 vccd1 vccd1 _4769_/A sky130_fd_sc_hd__nand2_1
X_3719_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3730_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4699_ _4704_/B _4704_/A vssd1 vssd1 vccd1 vccd1 _4705_/B sky130_fd_sc_hd__nor2_1
Xhold22 hold22/A vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2952_ _2603_/X _2949_/Y _2903_/X _2951_/Y vssd1 vssd1 vccd1 vccd1 _5232_/D sky130_fd_sc_hd__o211a_1
X_2883_ _2803_/X _2879_/Y _2880_/X _2808_/X _2882_/Y vssd1 vssd1 vccd1 vccd1 _5245_/D
+ sky130_fd_sc_hd__o311a_1
X_4622_ _5010_/Q _5042_/Q vssd1 vssd1 vccd1 vccd1 _4637_/C sky130_fd_sc_hd__nor2_1
X_4553_ _4546_/Y _4550_/X _4544_/B _4552_/Y vssd1 vssd1 vccd1 vccd1 _4554_/A sky130_fd_sc_hd__a211oi_1
X_4484_ _4484_/A _4484_/B vssd1 vssd1 vccd1 vccd1 _4490_/A sky130_fd_sc_hd__nor2_1
X_3504_ _3504_/A _3504_/B _3504_/C vssd1 vssd1 vccd1 vccd1 _3504_/Y sky130_fd_sc_hd__nand3_1
X_3435_ _3808_/B _5110_/Q vssd1 vssd1 vccd1 vccd1 _3436_/B sky130_fd_sc_hd__and2_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3366_ _3795_/B _5115_/Q vssd1 vssd1 vccd1 vccd1 _3571_/B sky130_fd_sc_hd__and2_1
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ _5203_/CLK _5105_/D vssd1 vssd1 vccd1 vccd1 _5105_/Q sky130_fd_sc_hd__dfxtp_1
X_3297_ _3297_/A _3297_/B vssd1 vssd1 vccd1 vccd1 _3301_/A sky130_fd_sc_hd__nor2_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _5068_/CLK _5036_/D vssd1 vssd1 vccd1 vccd1 _5036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput34 _5181_/Q vssd1 vssd1 vccd1 vccd1 data_out[19] sky130_fd_sc_hd__buf_2
Xoutput56 _4939_/X vssd1 vssd1 vccd1 vccd1 data_valid_out sky130_fd_sc_hd__buf_2
Xoutput45 _5191_/Q vssd1 vssd1 vccd1 vccd1 data_out[29] sky130_fd_sc_hd__buf_2
XFILLER_0_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3220_ _5214_/Q _2928_/X _2962_/X _3219_/X vssd1 vssd1 vccd1 vccd1 _5214_/D sky130_fd_sc_hd__o211a_1
X_3151_ _3175_/A vssd1 vssd1 vccd1 vccd1 _3151_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3082_ _3267_/B _3082_/B vssd1 vssd1 vccd1 vccd1 _3271_/B sky130_fd_sc_hd__nand2_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _4956_/Q _4956_/D vssd1 vssd1 vccd1 vccd1 _4027_/A sky130_fd_sc_hd__xnor2_4
XFILLER_62_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2935_ _2935_/A _2935_/B vssd1 vssd1 vccd1 vccd1 _2935_/Y sky130_fd_sc_hd__nor2_1
X_2866_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2866_/X sky130_fd_sc_hd__buf_4
X_4605_ _4779_/B _4779_/A _4785_/B vssd1 vssd1 vccd1 vccd1 _4605_/X sky130_fd_sc_hd__or3_1
X_2797_ _2755_/Y _2797_/B _2797_/C vssd1 vssd1 vccd1 vccd1 _2798_/C sky130_fd_sc_hd__nand3b_1
X_4536_ _4535_/B _4534_/Y _4535_/Y _5055_/Q _4873_/A vssd1 vssd1 vccd1 vccd1 _5023_/D
+ sky130_fd_sc_hd__a221oi_1
XFILLER_89_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4467_ _4466_/B _4466_/A _4436_/X vssd1 vssd1 vccd1 vccd1 _4467_/X sky130_fd_sc_hd__a21o_1
X_4398_ _4701_/A vssd1 vssd1 vccd1 vccd1 _4746_/A sky130_fd_sc_hd__buf_2
X_3418_ _5202_/Q _5106_/Q vssd1 vssd1 vccd1 vccd1 _3621_/B sky130_fd_sc_hd__xor2_1
XFILLER_58_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3349_ _3774_/B _5123_/Q vssd1 vssd1 vccd1 vccd1 _3531_/B sky130_fd_sc_hd__and2_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5019_ _5272_/CLK _5019_/D vssd1 vssd1 vccd1 vccd1 _5019_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2720_ _2713_/Y _2715_/Y _2719_/X vssd1 vssd1 vccd1 vccd1 _2720_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_12_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2651_ _5267_/Q _4598_/A vssd1 vssd1 vccd1 vccd1 _2683_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2582_ _2594_/A _4589_/A vssd1 vssd1 vccd1 vccd1 _2582_/Y sky130_fd_sc_hd__nand2_1
X_4321_ _4321_/A _4321_/B vssd1 vssd1 vccd1 vccd1 _4423_/B sky130_fd_sc_hd__nor2_1
X_4252_ _5057_/Q _5025_/Q vssd1 vssd1 vccd1 vccd1 _4524_/A sky130_fd_sc_hd__or2_1
X_3203_ _3218_/B _3218_/A vssd1 vssd1 vccd1 vccd1 _3203_/Y sky130_fd_sc_hd__nand2_1
X_4183_ _4183_/A vssd1 vssd1 vccd1 vccd1 _4183_/X sky130_fd_sc_hd__buf_4
XFILLER_67_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3134_ _3201_/A _3201_/B _3133_/Y vssd1 vssd1 vccd1 vccd1 _3196_/A sky130_fd_sc_hd__o21bai_2
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3065_ _5136_/Q _3740_/B vssd1 vssd1 vccd1 vccd1 _3287_/B sky130_fd_sc_hd__or2_1
XFILLER_23_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3967_ _3967_/A _3967_/B vssd1 vssd1 vccd1 vccd1 _3975_/C sky130_fd_sc_hd__or2_1
X_2918_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3826_/A sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_30_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5193_/CLK sky130_fd_sc_hd__clkbuf_16
X_3898_ _4982_/Q _3898_/B vssd1 vssd1 vccd1 vccd1 _3898_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2849_ _2849_/A vssd1 vssd1 vccd1 vccd1 _3598_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4519_ _4520_/B _4520_/C _4520_/A vssd1 vssd1 vccd1 vccd1 _4519_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4964_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4870_ _4870_/A vssd1 vssd1 vccd1 vccd1 _4977_/D sky130_fd_sc_hd__clkbuf_1
X_3821_ _5106_/Q _3819_/X _3816_/X _3820_/Y vssd1 vssd1 vccd1 vccd1 _5106_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5080_/CLK sky130_fd_sc_hd__clkbuf_16
X_3752_ _5132_/Q _3739_/X _3750_/X _3751_/Y vssd1 vssd1 vccd1 vccd1 _5132_/D sky130_fd_sc_hd__o211a_1
X_3683_ _3690_/A hold17/X vssd1 vssd1 vccd1 vccd1 _3683_/Y sky130_fd_sc_hd__nand2_1
X_2703_ _2908_/A _2908_/B _2702_/Y vssd1 vssd1 vccd1 vccd1 _2703_/Y sky130_fd_sc_hd__a21oi_1
X_2634_ _2635_/B _2880_/C vssd1 vssd1 vccd1 vccd1 _2644_/B sky130_fd_sc_hd__nor2_1
X_2565_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2565_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4304_ _4304_/A _4623_/B vssd1 vssd1 vccd1 vccd1 _4305_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5284_ _5287_/CLK hold13/X vssd1 vssd1 vccd1 vccd1 _5284_/Q sky130_fd_sc_hd__dfxtp_1
X_2496_ _2496_/A hold24/X vssd1 vssd1 vccd1 vccd1 _2496_/Y sky130_fd_sc_hd__nand2_1
X_4235_ _4235_/A _4563_/B vssd1 vssd1 vccd1 vccd1 _4476_/B sky130_fd_sc_hd__nor2_1
XFILLER_4_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4166_ _4166_/A _4760_/A _4166_/C vssd1 vssd1 vccd1 vccd1 _4167_/A sky130_fd_sc_hd__and3_1
XFILLER_28_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3117_ _3699_/B _5151_/Q vssd1 vssd1 vccd1 vccd1 _3118_/B sky130_fd_sc_hd__and2_1
XFILLER_82_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4097_ _4097_/A vssd1 vssd1 vccd1 vccd1 _4098_/C sky130_fd_sc_hd__inv_2
XFILLER_82_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3048_ _5133_/Q vssd1 vssd1 vccd1 vccd1 _3048_/Y sky130_fd_sc_hd__inv_2
XFILLER_90_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4999_ _5265_/CLK _4999_/D vssd1 vssd1 vccd1 vccd1 _4999_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4020_ _4020_/A _4020_/B _4020_/C vssd1 vssd1 vccd1 vccd1 _4021_/B sky130_fd_sc_hd__nand3_1
Xclkbuf_leaf_1_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5137_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_49_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4922_ _4922_/A vssd1 vssd1 vccd1 vccd1 _4922_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4853_ _4853_/A _4853_/B vssd1 vssd1 vccd1 vccd1 _4854_/A sky130_fd_sc_hd__and2_1
X_3804_ _5112_/Q _3792_/X _3802_/X _3803_/Y vssd1 vssd1 vccd1 vccd1 _5112_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4784_ _4784_/A vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__buf_2
X_3735_ _3735_/A vssd1 vssd1 vccd1 vccd1 _3735_/X sky130_fd_sc_hd__buf_2
X_3666_ _5163_/Q _3634_/X _3664_/Y _3665_/X _3642_/X vssd1 vssd1 vccd1 vccd1 _5163_/D
+ sky130_fd_sc_hd__o221a_1
X_3597_ _3597_/A _3597_/B vssd1 vssd1 vccd1 vccd1 _3597_/Y sky130_fd_sc_hd__nor2_1
X_2617_ _5284_/Q _4656_/A vssd1 vssd1 vccd1 vccd1 _2828_/C sky130_fd_sc_hd__or2_1
X_2548_ _5006_/Q vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__inv_2
X_5267_ _5288_/CLK _5267_/D vssd1 vssd1 vccd1 vccd1 _5267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2479_ _2600_/A vssd1 vssd1 vccd1 vccd1 _2836_/A sky130_fd_sc_hd__clkbuf_1
X_4218_ _5043_/Q vssd1 vssd1 vccd1 vccd1 _4548_/B sky130_fd_sc_hd__inv_2
X_5198_ _5209_/CLK _5198_/D vssd1 vssd1 vccd1 vccd1 _5198_/Q sky130_fd_sc_hd__dfxtp_1
X_4149_ _4151_/A _5064_/Q _4141_/C _4873_/A vssd1 vssd1 vccd1 vccd1 _4149_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_55_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3520_ _3538_/A _3538_/C vssd1 vssd1 vccd1 vccd1 _3532_/B sky130_fd_sc_hd__and2_1
X_3451_ _3573_/B _3451_/B vssd1 vssd1 vccd1 vccd1 _3576_/B sky130_fd_sc_hd__nand2_1
X_3382_ _3820_/B _5106_/Q _3419_/B vssd1 vssd1 vccd1 vccd1 _3384_/A sky130_fd_sc_hd__or3b_1
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5121_ _5195_/CLK _5121_/D vssd1 vssd1 vccd1 vccd1 _5121_/Q sky130_fd_sc_hd__dfxtp_1
X_5052_ _5086_/CLK _5052_/D vssd1 vssd1 vccd1 vccd1 _5052_/Q sky130_fd_sc_hd__dfxtp_2
X_4003_ _4003_/A _4003_/B vssd1 vssd1 vccd1 vccd1 _4004_/B sky130_fd_sc_hd__and2_1
XFILLER_77_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4905_ _4905_/A vssd1 vssd1 vccd1 vccd1 _4905_/X sky130_fd_sc_hd__clkbuf_1
X_4836_ _4988_/Q vssd1 vssd1 vccd1 vccd1 _4846_/B sky130_fd_sc_hd__inv_2
X_4767_ _4767_/A _4767_/B vssd1 vssd1 vccd1 vccd1 _4774_/B sky130_fd_sc_hd__or2_1
X_4698_ _4704_/B _4704_/A _4661_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4698_/X sky130_fd_sc_hd__o211a_1
X_3718_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3773_/A sky130_fd_sc_hd__buf_2
X_3649_ _3649_/A _3649_/B vssd1 vssd1 vccd1 vccd1 _3651_/A sky130_fd_sc_hd__nand2_1
XFILLER_88_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold12 hold12/A vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold23 hold23/A vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_29_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2951_ _3199_/A _3740_/B vssd1 vssd1 vccd1 vccd1 _2951_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2882_ _3238_/A _3703_/B vssd1 vssd1 vccd1 vccd1 _2882_/Y sky130_fd_sc_hd__nand2_1
X_4621_ _4756_/A _4756_/B _4620_/Y vssd1 vssd1 vccd1 vccd1 _4737_/B sky130_fd_sc_hd__a21oi_1
XFILLER_30_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4552_ _4552_/A _4722_/B vssd1 vssd1 vccd1 vccd1 _4552_/Y sky130_fd_sc_hd__nor2_1
X_4483_ _4987_/Q _5033_/Q _4469_/X _4482_/X vssd1 vssd1 vccd1 vccd1 _5033_/D sky130_fd_sc_hd__o211a_1
X_3503_ _3507_/A _3503_/B _3503_/C vssd1 vssd1 vccd1 vccd1 _3504_/A sky130_fd_sc_hd__nand3b_1
XFILLER_89_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3434_ _3434_/A vssd1 vssd1 vccd1 vccd1 _3593_/B sky130_fd_sc_hd__inv_2
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ _5211_/Q vssd1 vssd1 vccd1 vccd1 _3795_/B sky130_fd_sc_hd__inv_2
XFILLER_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5104_ _5203_/CLK _5104_/D vssd1 vssd1 vccd1 vccd1 _5104_/Q sky130_fd_sc_hd__dfxtp_1
X_3296_ _5135_/Q _3742_/B vssd1 vssd1 vccd1 vccd1 _3297_/B sky130_fd_sc_hd__nor2_1
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _5068_/CLK _5035_/D vssd1 vssd1 vccd1 vccd1 _5035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4819_ _4819_/A _4819_/B _4819_/C vssd1 vssd1 vccd1 vccd1 _4819_/X sky130_fd_sc_hd__and3_1
XFILLER_5_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput24 _5162_/Q vssd1 vssd1 vccd1 vccd1 data_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput46 _5164_/Q vssd1 vssd1 vccd1 vccd1 data_out[2] sky130_fd_sc_hd__buf_2
Xoutput35 _5163_/Q vssd1 vssd1 vccd1 vccd1 data_out[1] sky130_fd_sc_hd__buf_2
XFILLER_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3150_ _5158_/Q _3679_/B vssd1 vssd1 vccd1 vccd1 _3175_/A sky130_fd_sc_hd__nor2_1
XFILLER_79_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3081_ _3728_/B _5140_/Q vssd1 vssd1 vccd1 vccd1 _3082_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3983_ _3987_/B _3987_/A _3992_/A _3982_/X vssd1 vssd1 vccd1 vccd1 _4026_/A sky130_fd_sc_hd__o22ai_4
X_2934_ _2938_/A _2938_/B _2681_/A vssd1 vssd1 vccd1 vccd1 _2935_/B sky130_fd_sc_hd__o21a_1
XFILLER_30_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2865_ _2870_/B _2854_/B _2733_/X vssd1 vssd1 vccd1 vccd1 _2865_/Y sky130_fd_sc_hd__a21oi_1
X_4604_ _4604_/A _4781_/C vssd1 vssd1 vccd1 vccd1 _4785_/B sky130_fd_sc_hd__nand2_1
X_4535_ _4535_/A _4535_/B vssd1 vssd1 vccd1 vccd1 _4535_/Y sky130_fd_sc_hd__nor2_1
X_2796_ _2978_/A vssd1 vssd1 vccd1 vccd1 _3504_/C sky130_fd_sc_hd__buf_2
XFILLER_89_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4466_ _4466_/A _4466_/B vssd1 vssd1 vccd1 vccd1 _4466_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4397_ _4745_/A _4397_/B _4397_/C vssd1 vssd1 vccd1 vccd1 _4397_/X sky130_fd_sc_hd__or3_1
X_3417_ _3414_/B _3626_/B _3414_/A vssd1 vssd1 vccd1 vccd1 _3615_/B sky130_fd_sc_hd__o21ba_1
XFILLER_58_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3348_ _5122_/Q _3777_/B vssd1 vssd1 vccd1 vccd1 _3533_/A sky130_fd_sc_hd__nor2_1
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3279_ _3279_/A _3279_/B vssd1 vssd1 vccd1 vccd1 _3279_/Y sky130_fd_sc_hd__nor2_1
X_5018_ _5272_/CLK _5018_/D vssd1 vssd1 vccd1 vccd1 _5018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2650_ _5266_/Q _4794_/A vssd1 vssd1 vccd1 vccd1 _2681_/A sky130_fd_sc_hd__or2_1
X_2581_ _4997_/Q vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__inv_2
X_4320_ _4304_/A _4623_/B _4318_/Y _4316_/A _4319_/X vssd1 vssd1 vccd1 vccd1 _4427_/B
+ sky130_fd_sc_hd__o221a_1
X_4251_ _5056_/Q _5024_/Q _5055_/Q _5023_/Q vssd1 vssd1 vccd1 vccd1 _4523_/B sky130_fd_sc_hd__o211a_1
X_3202_ _3202_/A vssd1 vssd1 vccd1 vccd1 _3218_/A sky130_fd_sc_hd__inv_2
X_4182_ _4185_/A _4178_/Y _4179_/Y _4181_/X vssd1 vssd1 vccd1 vccd1 _4182_/X sky130_fd_sc_hd__a31o_1
X_3133_ _3133_/A vssd1 vssd1 vccd1 vccd1 _3133_/Y sky130_fd_sc_hd__clkinv_2
XFILLER_55_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3064_ _3297_/A vssd1 vssd1 vccd1 vccd1 _3064_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3966_ _4968_/Q _4968_/D vssd1 vssd1 vccd1 vccd1 _3967_/B sky130_fd_sc_hd__and2_1
X_2917_ _2917_/A _2917_/B vssd1 vssd1 vccd1 vccd1 _2917_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3897_ _3897_/A _3897_/B _3897_/C _3897_/D vssd1 vssd1 vccd1 vccd1 _3897_/X sky130_fd_sc_hd__and4_1
X_2848_ _2843_/B _2841_/C _2841_/A vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__a21o_1
X_2779_ _2874_/A _2874_/B _2719_/X vssd1 vssd1 vccd1 vccd1 _2869_/A sky130_fd_sc_hd__o21bai_1
X_4518_ _4518_/A vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__inv_2
XFILLER_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4449_ _4987_/Q _5040_/Q _4446_/X _4448_/Y _4438_/X vssd1 vssd1 vccd1 vccd1 _5040_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_77_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3820_ _3824_/A _3820_/B vssd1 vssd1 vccd1 vccd1 _3820_/Y sky130_fd_sc_hd__nand2_1
X_3751_ _3758_/A _3751_/B vssd1 vssd1 vccd1 vccd1 _3751_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2702_ _2911_/A _2916_/A vssd1 vssd1 vccd1 vccd1 _2702_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3682_ _3735_/A vssd1 vssd1 vccd1 vccd1 _3682_/X sky130_fd_sc_hd__clkbuf_2
X_2633_ _5276_/Q _4637_/A vssd1 vssd1 vccd1 vccd1 _2880_/C sky130_fd_sc_hd__or2_1
X_2564_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2564_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4303_ _5042_/Q vssd1 vssd1 vccd1 vccd1 _4623_/B sky130_fd_sc_hd__inv_2
X_2495_ _5019_/Q vssd1 vssd1 vccd1 vccd1 hold24/A sky130_fd_sc_hd__clkinv_2
XFILLER_59_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5283_ _5283_/CLK _5283_/D vssd1 vssd1 vccd1 vccd1 _5283_/Q sky130_fd_sc_hd__dfxtp_1
X_4234_ _5034_/Q vssd1 vssd1 vccd1 vccd1 _4563_/B sky130_fd_sc_hd__inv_2
X_4165_ _4701_/A _4162_/C _4247_/A vssd1 vssd1 vccd1 vccd1 _4166_/C sky130_fd_sc_hd__o21ai_1
XFILLER_67_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3116_ _5151_/Q _3699_/B vssd1 vssd1 vccd1 vccd1 _3118_/A sky130_fd_sc_hd__nor2_1
XFILLER_28_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4096_ _4110_/B _4096_/B vssd1 vssd1 vccd1 vccd1 _4097_/A sky130_fd_sc_hd__nand2_1
X_3047_ _3742_/B _5135_/Q _3299_/B vssd1 vssd1 vccd1 vccd1 _3047_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4998_ _5265_/CLK _4998_/D vssd1 vssd1 vccd1 vccd1 _4998_/Q sky130_fd_sc_hd__dfxtp_1
X_3949_ _3949_/A _4003_/B vssd1 vssd1 vccd1 vccd1 _3993_/B sky130_fd_sc_hd__and2_1
XFILLER_58_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4921_ _4936_/B _4925_/A _4921_/C vssd1 vssd1 vccd1 vccd1 _4922_/A sky130_fd_sc_hd__and3_1
XFILLER_33_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4852_ _4852_/A vssd1 vssd1 vccd1 vccd1 _4986_/D sky130_fd_sc_hd__clkbuf_1
X_3803_ _3810_/A _3803_/B vssd1 vssd1 vccd1 vccd1 _3803_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4783_ _4516_/X _4780_/Y _4781_/X _4760_/X _4782_/Y vssd1 vssd1 vccd1 vccd1 _5002_/D
+ sky130_fd_sc_hd__o311a_1
X_3734_ _5138_/Q _3725_/X _3722_/X _3733_/Y vssd1 vssd1 vccd1 vccd1 _5138_/D sky130_fd_sc_hd__o211a_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3665_ _3668_/B _3664_/B _2866_/X vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__a21o_1
X_2616_ _4702_/A _5285_/Q vssd1 vssd1 vccd1 vccd1 _2622_/B sky130_fd_sc_hd__and2_1
X_3596_ _3808_/B _5110_/Q _3595_/X vssd1 vssd1 vccd1 vccd1 _3597_/B sky130_fd_sc_hd__o21a_1
X_2547_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2547_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2478_ _4841_/A _4871_/B vssd1 vssd1 vccd1 vccd1 _2600_/A sky130_fd_sc_hd__nor2_2
X_5266_ _5288_/CLK _5266_/D vssd1 vssd1 vccd1 vccd1 _5266_/Q sky130_fd_sc_hd__dfxtp_1
X_4217_ _4321_/B vssd1 vssd1 vccd1 vccd1 _4217_/Y sky130_fd_sc_hd__inv_2
X_5197_ _5219_/CLK _5197_/D vssd1 vssd1 vccd1 vccd1 _5197_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_28_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _4146_/Y _4278_/A _4147_/X vssd1 vssd1 vccd1 vccd1 _5065_/D sky130_fd_sc_hd__a21oi_1
X_4079_ _4092_/B _5080_/Q _5079_/Q vssd1 vssd1 vccd1 vccd1 _4080_/A sky130_fd_sc_hd__and3_1
XFILLER_28_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_3_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3450_ _3797_/B _5114_/Q vssd1 vssd1 vccd1 vccd1 _3451_/B sky130_fd_sc_hd__nand2_1
X_3381_ _3817_/B _5107_/Q vssd1 vssd1 vccd1 vccd1 _3419_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5120_ _5219_/CLK _5120_/D vssd1 vssd1 vccd1 vccd1 _5120_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5051_ _5051_/CLK _5051_/D vssd1 vssd1 vccd1 vccd1 _5051_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4002_ _4002_/A vssd1 vssd1 vccd1 vccd1 _4004_/A sky130_fd_sc_hd__inv_2
XFILLER_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4904_ _4915_/A _4904_/B vssd1 vssd1 vccd1 vccd1 _4905_/A sky130_fd_sc_hd__and2_1
X_4835_ _4989_/Q vssd1 vssd1 vccd1 vccd1 _4840_/A sky130_fd_sc_hd__inv_2
X_4766_ _4766_/A vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__inv_2
X_3717_ _5144_/Q _3711_/X _3708_/X _3716_/Y vssd1 vssd1 vccd1 vccd1 _5144_/D sky130_fd_sc_hd__o211a_1
X_4697_ _4696_/X _4663_/A _4665_/X vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__a21oi_2
XFILLER_20_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3648_ _3833_/B _5101_/Q vssd1 vssd1 vccd1 vccd1 _3649_/B sky130_fd_sc_hd__nand2_1
XFILLER_88_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3579_ _5178_/Q _3537_/X _3303_/X _3578_/X vssd1 vssd1 vccd1 vccd1 _5178_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold13 hold13/A vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold24 hold24/A vssd1 vssd1 vccd1 vccd1 hold24/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_5249_ _5282_/CLK _5249_/D vssd1 vssd1 vccd1 vccd1 _5249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2950_ _5232_/Q vssd1 vssd1 vccd1 vccd1 _3740_/B sky130_fd_sc_hd__clkinv_2
X_2881_ _5245_/Q vssd1 vssd1 vccd1 vccd1 _3703_/B sky130_fd_sc_hd__inv_2
X_4620_ _4759_/B _4763_/A vssd1 vssd1 vccd1 vccd1 _4620_/Y sky130_fd_sc_hd__nand2_1
X_4551_ _4551_/A vssd1 vssd1 vccd1 vccd1 _4722_/B sky130_fd_sc_hd__inv_2
X_4482_ _4478_/A _4481_/Y _4407_/X vssd1 vssd1 vccd1 vccd1 _4482_/X sky130_fd_sc_hd__a21o_1
X_3502_ _3502_/A _3502_/B vssd1 vssd1 vccd1 vccd1 _3503_/C sky130_fd_sc_hd__nor2_1
X_3433_ _3429_/B _3607_/B _3429_/A vssd1 vssd1 vccd1 vccd1 _3594_/B sky130_fd_sc_hd__o21ba_1
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _5168_/CLK _5103_/D vssd1 vssd1 vccd1 vccd1 _5103_/Q sky130_fd_sc_hd__dfxtp_1
X_3364_ _3370_/B _3364_/B vssd1 vssd1 vccd1 vccd1 _3566_/B sky130_fd_sc_hd__nand2_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _3295_/A vssd1 vssd1 vccd1 vccd1 _3299_/A sky130_fd_sc_hd__inv_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _5068_/CLK _5034_/D vssd1 vssd1 vccd1 vccd1 _5034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4818_ _4819_/B _4819_/C _4819_/A vssd1 vssd1 vccd1 vccd1 _4818_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4749_ _4753_/A _4753_/B _4632_/A vssd1 vssd1 vccd1 vccd1 _4750_/B sky130_fd_sc_hd__o21a_1
Xoutput25 _5172_/Q vssd1 vssd1 vccd1 vccd1 data_out[10] sky130_fd_sc_hd__buf_2
Xoutput36 _5182_/Q vssd1 vssd1 vccd1 vccd1 data_out[20] sky130_fd_sc_hd__buf_2
Xoutput47 _5192_/Q vssd1 vssd1 vccd1 vccd1 data_out[30] sky130_fd_sc_hd__buf_2
XFILLER_63_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3080_ _5140_/Q _3728_/B vssd1 vssd1 vccd1 vccd1 _3267_/B sky130_fd_sc_hd__or2_1
XFILLER_39_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3982_ _3969_/X _3979_/Y _3986_/B _3986_/A vssd1 vssd1 vccd1 vccd1 _3982_/X sky130_fd_sc_hd__o211a_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2933_ _2933_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _2938_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2864_ _5248_/Q _2847_/X _2609_/X _2863_/X vssd1 vssd1 vccd1 vccd1 _5248_/D sky130_fd_sc_hd__o211a_1
X_2795_ _2764_/Y _2788_/Y _2794_/Y vssd1 vssd1 vccd1 vccd1 _5257_/D sky130_fd_sc_hd__a21oi_1
X_4603_ _4603_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _4604_/A sky130_fd_sc_hd__nand2_1
X_4534_ _4987_/Q _5055_/Q vssd1 vssd1 vccd1 vccd1 _4534_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4465_ _4471_/B _4471_/A _4285_/B vssd1 vssd1 vccd1 vccd1 _4466_/B sky130_fd_sc_hd__o21ai_1
X_4396_ _4396_/A _4396_/B _4396_/C vssd1 vssd1 vccd1 vccd1 _4397_/B sky130_fd_sc_hd__and3_1
X_3416_ _3388_/Y _3635_/A _3406_/Y _3415_/Y vssd1 vssd1 vccd1 vccd1 _3615_/A sky130_fd_sc_hd__o211ai_1
X_3347_ _5123_/Q _3774_/B vssd1 vssd1 vccd1 vccd1 _3531_/A sky130_fd_sc_hd__nor2_1
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _3733_/B _5138_/Q _3277_/X vssd1 vssd1 vccd1 vccd1 _3279_/B sky130_fd_sc_hd__o21a_1
X_5017_ _5272_/CLK _5017_/D vssd1 vssd1 vccd1 vccd1 _5017_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_73_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2580_ _5265_/Q _2564_/X _2565_/X _2579_/Y vssd1 vssd1 vccd1 vccd1 _5265_/D sky130_fd_sc_hd__o211a_1
X_4250_ _5056_/Q _5024_/Q vssd1 vssd1 vccd1 vccd1 _4529_/B sky130_fd_sc_hd__and2_1
XFILLER_4_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4181_ _4711_/A vssd1 vssd1 vccd1 vccd1 _4181_/X sky130_fd_sc_hd__clkbuf_4
X_3201_ _3201_/A _3201_/B vssd1 vssd1 vccd1 vccd1 _3218_/B sky130_fd_sc_hd__or2_1
X_3132_ _3132_/A _3202_/A _3132_/C vssd1 vssd1 vccd1 vccd1 _3133_/A sky130_fd_sc_hd__nor3_1
X_3063_ _5231_/Q _3063_/B vssd1 vssd1 vccd1 vccd1 _3297_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3965_ _4968_/Q _4968_/D vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3896_ _5090_/Q _3895_/Y _4890_/A _4979_/Q vssd1 vssd1 vccd1 vccd1 _3897_/D sky130_fd_sc_hd__o22a_1
X_2916_ _2916_/A _2916_/B vssd1 vssd1 vccd1 vccd1 _2916_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2847_ _3601_/A vssd1 vssd1 vccd1 vccd1 _2847_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_12_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2778_ _2896_/A _2896_/B _2712_/Y vssd1 vssd1 vccd1 vccd1 _2874_/B sky130_fd_sc_hd__a21oi_1
X_4517_ _4517_/A _4524_/B vssd1 vssd1 vccd1 vccd1 _4518_/A sky130_fd_sc_hd__nand2_1
X_4448_ _4448_/A _4448_/B vssd1 vssd1 vccd1 vccd1 _4448_/Y sky130_fd_sc_hd__nor2_1
X_4379_ _4379_/A _4987_/Q vssd1 vssd1 vccd1 vccd1 _4379_/Y sky130_fd_sc_hd__nand2_1
XFILLER_58_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _3802_/A vssd1 vssd1 vccd1 vccd1 _3750_/X sky130_fd_sc_hd__clkbuf_2
X_2701_ _2917_/A vssd1 vssd1 vccd1 vccd1 _2916_/A sky130_fd_sc_hd__inv_2
XFILLER_9_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3681_ _4089_/A vssd1 vssd1 vccd1 vccd1 _3735_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2632_ _4623_/A _5277_/Q vssd1 vssd1 vccd1 vccd1 _2635_/B sky130_fd_sc_hd__and2_1
X_2563_ _5269_/Q _2544_/X _2547_/X _2562_/Y vssd1 vssd1 vccd1 vccd1 _5269_/D sky130_fd_sc_hd__o211a_1
X_4302_ _5074_/Q _5042_/Q vssd1 vssd1 vccd1 vccd1 _4319_/B sky130_fd_sc_hd__nor2_1
X_5282_ _5282_/CLK _5282_/D vssd1 vssd1 vccd1 vccd1 _5282_/Q sky130_fd_sc_hd__dfxtp_1
X_4233_ _5065_/Q _5033_/Q vssd1 vssd1 vccd1 vccd1 _4478_/C sky130_fd_sc_hd__nand2_1
X_2494_ _5287_/Q _2481_/X _2485_/X _2493_/Y vssd1 vssd1 vccd1 vccd1 _5287_/D sky130_fd_sc_hd__o211a_1
X_4164_ _4244_/A _4166_/A _4163_/X vssd1 vssd1 vccd1 vccd1 _5060_/D sky130_fd_sc_hd__a21oi_1
X_4095_ _5078_/Q vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__inv_2
XFILLER_28_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3115_ _5247_/Q vssd1 vssd1 vccd1 vccd1 _3699_/B sky130_fd_sc_hd__inv_2
X_3046_ _5134_/Q _3744_/B vssd1 vssd1 vccd1 vccd1 _3299_/B sky130_fd_sc_hd__or2_1
XFILLER_55_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4997_ _5265_/CLK _4997_/D vssd1 vssd1 vccd1 vccd1 _4997_/Q sky130_fd_sc_hd__dfxtp_1
X_3948_ _4003_/B _3949_/A vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__nor2_1
X_3879_ _3879_/A _4890_/A vssd1 vssd1 vccd1 vccd1 _3879_/Y sky130_fd_sc_hd__nand2_1
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4920_ _4920_/A vssd1 vssd1 vccd1 vccd1 _4920_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _4853_/A _4851_/B vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__and2_1
XFILLER_60_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3802_ _3802_/A vssd1 vssd1 vccd1 vccd1 _3802_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4782_ _4782_/A _4794_/B vssd1 vssd1 vccd1 vccd1 _4782_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3733_ _3744_/A _3733_/B vssd1 vssd1 vccd1 vccd1 _3733_/Y sky130_fd_sc_hd__nand2_1
X_3664_ _3668_/B _3664_/B vssd1 vssd1 vccd1 vccd1 _3664_/Y sky130_fd_sc_hd__nor2_1
X_2615_ _5285_/Q _4702_/A vssd1 vssd1 vccd1 vccd1 _2630_/A sky130_fd_sc_hd__nor2_1
X_3595_ _3602_/B _3602_/A vssd1 vssd1 vccd1 vccd1 _3595_/X sky130_fd_sc_hd__or2_1
X_2546_ _4089_/A vssd1 vssd1 vccd1 vccd1 _2903_/A sky130_fd_sc_hd__buf_2
X_2477_ _5087_/Q vssd1 vssd1 vccd1 vccd1 _4871_/B sky130_fd_sc_hd__inv_2
X_5265_ _5265_/CLK _5265_/D vssd1 vssd1 vccd1 vccd1 _5265_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4216_ _4216_/A _4547_/B vssd1 vssd1 vccd1 vccd1 _4321_/B sky130_fd_sc_hd__nor2_1
X_5196_ _5219_/CLK _5196_/D vssd1 vssd1 vccd1 vccd1 _5196_/Q sky130_fd_sc_hd__dfxtp_2
X_4147_ _4163_/B _4142_/B _4141_/C _4873_/A vssd1 vssd1 vccd1 vccd1 _4147_/X sky130_fd_sc_hd__a31o_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4078_ _4873_/A _4078_/B _4078_/C vssd1 vssd1 vccd1 vccd1 _5083_/D sky130_fd_sc_hd__nor3_1
XFILLER_43_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3029_ _5146_/Q _3712_/B vssd1 vssd1 vccd1 vccd1 _3110_/A sky130_fd_sc_hd__nor2_1
XFILLER_51_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3380_ _5203_/Q vssd1 vssd1 vccd1 vccd1 _3817_/B sky130_fd_sc_hd__inv_2
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5050_ _5051_/CLK _5050_/D vssd1 vssd1 vccd1 vccd1 _5050_/Q sky130_fd_sc_hd__dfxtp_1
X_4001_ _4001_/A _4001_/B _4001_/C vssd1 vssd1 vccd1 vccd1 _4009_/C sky130_fd_sc_hd__nand3_2
XFILLER_77_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4903_ _4903_/A _4907_/A vssd1 vssd1 vccd1 vccd1 _4904_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4834_ _4952_/X vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__inv_2
X_4765_ _3886_/X _4763_/Y _4715_/X _4764_/Y vssd1 vssd1 vccd1 vccd1 _5005_/D sky130_fd_sc_hd__o211a_1
X_3716_ _3716_/A _3716_/B vssd1 vssd1 vccd1 vccd1 _3716_/Y sky130_fd_sc_hd__nand2_1
X_4696_ _4716_/A _4716_/B vssd1 vssd1 vccd1 vccd1 _4696_/X sky130_fd_sc_hd__or2_1
X_3647_ _5166_/Q _3601_/X _3644_/X _3646_/Y vssd1 vssd1 vccd1 vccd1 _5166_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3578_ _3573_/A _3576_/Y _3577_/X vssd1 vssd1 vccd1 vccd1 _3578_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2529_ _5278_/Q _2525_/X _2526_/X _2528_/Y vssd1 vssd1 vccd1 vccd1 _5278_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold14 hold14/A vssd1 vssd1 vccd1 vccd1 hold14/X sky130_fd_sc_hd__clkdlybuf4s25_1
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5248_ _5289_/CLK _5248_/D vssd1 vssd1 vccd1 vccd1 _5248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5179_ _5181_/CLK _5179_/D vssd1 vssd1 vccd1 vccd1 _5179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2880_ _2884_/A _2880_/B _2880_/C vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__and3_1
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4550_ _4639_/B _4641_/B _4639_/A vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__o21ba_1
X_4481_ _4481_/A _4481_/B vssd1 vssd1 vccd1 vccd1 _4481_/Y sky130_fd_sc_hd__nand2_1
X_3501_ _3485_/Y _3488_/Y _3507_/B vssd1 vssd1 vccd1 vccd1 _3503_/B sky130_fd_sc_hd__a21o_1
X_3432_ _3605_/A _3605_/B _3431_/X vssd1 vssd1 vccd1 vccd1 _3594_/A sky130_fd_sc_hd__o21bai_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ _3793_/B _5116_/Q vssd1 vssd1 vccd1 vccd1 _3364_/B sky130_fd_sc_hd__nand2_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _5203_/CLK _5102_/D vssd1 vssd1 vccd1 vccd1 _5102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _5200_/Q _3261_/X _3247_/X _3293_/X vssd1 vssd1 vccd1 vccd1 _5200_/D sky130_fd_sc_hd__o211a_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _5265_/CLK _5033_/D vssd1 vssd1 vccd1 vccd1 _5033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4817_ _4817_/A vssd1 vssd1 vccd1 vccd1 _4819_/A sky130_fd_sc_hd__inv_2
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4748_ _4748_/A _4748_/B vssd1 vssd1 vccd1 vccd1 _4750_/A sky130_fd_sc_hd__nor2_1
X_4679_ _4679_/A _4679_/B _4679_/C vssd1 vssd1 vccd1 vccd1 _4680_/C sky130_fd_sc_hd__and3_1
Xoutput26 _5173_/Q vssd1 vssd1 vccd1 vccd1 data_out[11] sky130_fd_sc_hd__buf_2
Xoutput37 _5183_/Q vssd1 vssd1 vccd1 vccd1 data_out[21] sky130_fd_sc_hd__buf_2
Xoutput48 _5193_/Q vssd1 vssd1 vccd1 vccd1 data_out[31] sky130_fd_sc_hd__buf_2
XFILLER_0_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3981_ _3981_/A _3981_/B vssd1 vssd1 vccd1 vccd1 _3986_/B sky130_fd_sc_hd__nor2_2
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2932_ _5236_/Q _2928_/X _2903_/X _2931_/X vssd1 vssd1 vccd1 vccd1 _5236_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_42_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5203_/CLK sky130_fd_sc_hd__clkbuf_16
X_2863_ _2856_/X _2862_/Y _2850_/X vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2794_ _5257_/Q _3668_/A _4115_/B vssd1 vssd1 vccd1 vccd1 _2794_/Y sky130_fd_sc_hd__o21ai_1
X_4602_ _4599_/A _4596_/B _4599_/B vssd1 vssd1 vccd1 vccd1 _4777_/B sky130_fd_sc_hd__o21ba_1
X_4533_ _5023_/Q vssd1 vssd1 vccd1 vccd1 _4535_/B sky130_fd_sc_hd__inv_2
X_4464_ _4464_/A vssd1 vssd1 vccd1 vccd1 _4471_/A sky130_fd_sc_hd__inv_2
X_4395_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__clkbuf_2
X_3415_ _3631_/B _3627_/A vssd1 vssd1 vccd1 vccd1 _3415_/Y sky130_fd_sc_hd__nor2_1
X_3346_ _5219_/Q vssd1 vssd1 vccd1 vccd1 _3774_/B sky130_fd_sc_hd__inv_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5016_ _5283_/CLK _5016_/D vssd1 vssd1 vccd1 vccd1 _5016_/Q sky130_fd_sc_hd__dfxtp_1
X_3277_ _3282_/B _3282_/A vssd1 vssd1 vccd1 vccd1 _3277_/X sky130_fd_sc_hd__or2_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_33_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5181_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_5_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_24_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _5265_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_40_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4180_ _4185_/A _4178_/Y _4179_/Y vssd1 vssd1 vccd1 vccd1 _4180_/Y sky130_fd_sc_hd__a21oi_1
X_3200_ _2603_/X _3197_/Y _2962_/X _3199_/Y vssd1 vssd1 vccd1 vccd1 _5218_/D sky130_fd_sc_hd__o211a_1
X_3131_ _3206_/B _3206_/A _3212_/B vssd1 vssd1 vccd1 vccd1 _3132_/C sky130_fd_sc_hd__or3_1
XFILLER_79_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3062_ _5135_/Q vssd1 vssd1 vccd1 vccd1 _3063_/B sky130_fd_sc_hd__inv_2
XFILLER_63_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3964_ _3964_/A _3964_/B _3996_/A vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__nand3_2
Xclkbuf_leaf_15_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5051_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2915_ _5239_/Q _2907_/X _2911_/Y _2913_/X _2914_/X vssd1 vssd1 vccd1 vccd1 _5239_/D
+ sky130_fd_sc_hd__o221a_1
X_3895_ _4980_/Q vssd1 vssd1 vccd1 vccd1 _3895_/Y sky130_fd_sc_hd__inv_2
X_2846_ _3738_/A vssd1 vssd1 vccd1 vccd1 _3601_/A sky130_fd_sc_hd__buf_2
X_2777_ _2777_/A vssd1 vssd1 vccd1 vccd1 _2896_/B sky130_fd_sc_hd__inv_2
X_4516_ _4535_/A vssd1 vssd1 vccd1 vccd1 _4516_/X sky130_fd_sc_hd__buf_2
X_4447_ _4447_/A _4447_/B vssd1 vssd1 vccd1 vccd1 _4448_/B sky130_fd_sc_hd__and2_1
X_4378_ _4378_/A _4378_/B _4383_/B _4378_/D vssd1 vssd1 vccd1 vccd1 _4379_/A sky130_fd_sc_hd__or4_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _5195_/Q _3307_/X _3327_/Y _3328_/X _3315_/X vssd1 vssd1 vccd1 vccd1 _5195_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2700_ _2700_/A _2700_/B vssd1 vssd1 vccd1 vccd1 _2917_/A sky130_fd_sc_hd__nand2_1
X_3680_ _5158_/Q _3671_/X _3644_/X _3679_/Y vssd1 vssd1 vccd1 vccd1 _5158_/D sky130_fd_sc_hd__o211a_1
X_2631_ _5277_/Q _4623_/A vssd1 vssd1 vccd1 vccd1 _2644_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2562_ _2573_/A _4782_/A vssd1 vssd1 vccd1 vccd1 _2562_/Y sky130_fd_sc_hd__nand2_1
X_4301_ _4301_/A _4434_/B vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__and2_1
X_5281_ _5281_/CLK _5281_/D vssd1 vssd1 vccd1 vccd1 _5281_/Q sky130_fd_sc_hd__dfxtp_1
X_4232_ _5066_/Q _5034_/Q vssd1 vssd1 vccd1 vccd1 _4476_/A sky130_fd_sc_hd__nor2_1
X_2493_ _2496_/A hold6/X vssd1 vssd1 vccd1 vccd1 _2493_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_4_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5251_/CLK sky130_fd_sc_hd__clkbuf_16
X_4163_ _4873_/A _4163_/B vssd1 vssd1 vccd1 vccd1 _4163_/X sky130_fd_sc_hd__or2_1
XFILLER_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4094_ _4327_/A _4099_/A _4093_/Y vssd1 vssd1 vccd1 vccd1 _5079_/D sky130_fd_sc_hd__a21oi_1
X_3114_ _3221_/A _3221_/B _3113_/X vssd1 vssd1 vccd1 vccd1 _3201_/B sky130_fd_sc_hd__a21oi_1
X_3045_ _5230_/Q vssd1 vssd1 vccd1 vccd1 _3744_/B sky130_fd_sc_hd__inv_2
XFILLER_23_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4996_ _4996_/CLK _4996_/D vssd1 vssd1 vccd1 vccd1 _4996_/Q sky130_fd_sc_hd__dfxtp_1
X_3947_ _4003_/A _4002_/A vssd1 vssd1 vccd1 vccd1 _3949_/A sky130_fd_sc_hd__nand2_1
XFILLER_11_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3878_ _5089_/Q vssd1 vssd1 vccd1 vccd1 _4890_/A sky130_fd_sc_hd__inv_2
X_2829_ _5253_/Q vssd1 vssd1 vccd1 vccd1 hold17/A sky130_fd_sc_hd__clkinv_2
XFILLER_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4850_ _4850_/A vssd1 vssd1 vccd1 vccd1 _4987_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3801_ _5113_/Q _3792_/X _3789_/X _3800_/Y vssd1 vssd1 vccd1 vccd1 _5113_/D sky130_fd_sc_hd__o211a_1
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4781_ _4781_/A _4781_/B _4781_/C vssd1 vssd1 vccd1 vccd1 _4781_/X sky130_fd_sc_hd__and3_1
X_3732_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3744_/A sky130_fd_sc_hd__clkbuf_2
X_3663_ _3663_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3664_/B sky130_fd_sc_hd__nand2_1
X_2614_ _5286_/Q vssd1 vssd1 vccd1 vccd1 _2815_/B sky130_fd_sc_hd__inv_2
X_3594_ _3594_/A _3594_/B vssd1 vssd1 vccd1 vccd1 _3602_/A sky130_fd_sc_hd__and2_1
X_2545_ _2791_/A vssd1 vssd1 vccd1 vccd1 _4089_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2476_ _4987_/Q vssd1 vssd1 vccd1 vccd1 _4841_/A sky130_fd_sc_hd__inv_2
X_5264_ _5265_/CLK _5264_/D vssd1 vssd1 vccd1 vccd1 _5264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5195_ _5195_/CLK _5195_/D vssd1 vssd1 vccd1 vccd1 _5195_/Q sky130_fd_sc_hd__dfxtp_2
X_4215_ _5044_/Q vssd1 vssd1 vccd1 vccd1 _4547_/B sky130_fd_sc_hd__inv_2
X_4146_ _4146_/A _5064_/Q vssd1 vssd1 vccd1 vccd1 _4146_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4077_ _4202_/A _4077_/B _4117_/C vssd1 vssd1 vccd1 vccd1 _4078_/C sky130_fd_sc_hd__nor3_1
XFILLER_55_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _5242_/Q vssd1 vssd1 vccd1 vccd1 _3712_/B sky130_fd_sc_hd__inv_2
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4979_ _5090_/CLK _4979_/D vssd1 vssd1 vccd1 vccd1 _4979_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_50_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4000_ _4000_/A _4000_/B vssd1 vssd1 vccd1 vccd1 _4001_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4902_ _4902_/A _4902_/B vssd1 vssd1 vccd1 vccd1 _4907_/A sky130_fd_sc_hd__nor2_1
X_4833_ _4387_/X _4828_/A _4991_/Q _4535_/Y _4772_/X vssd1 vssd1 vccd1 vccd1 _4991_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_60_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4764_ _4764_/A _4794_/B vssd1 vssd1 vccd1 vccd1 _4764_/Y sky130_fd_sc_hd__nand2_1
X_3715_ _5145_/Q _3711_/X _3708_/X _3714_/Y vssd1 vssd1 vccd1 vccd1 _5145_/D sky130_fd_sc_hd__o211a_1
X_4695_ _5019_/Q _4987_/Q _4693_/Y _4694_/X _4511_/X vssd1 vssd1 vccd1 vccd1 _5019_/D
+ sky130_fd_sc_hd__o221a_1
X_3646_ _3635_/A _3645_/X _3228_/B vssd1 vssd1 vccd1 vccd1 _3646_/Y sky130_fd_sc_hd__o21ai_1
X_3577_ _3577_/A vssd1 vssd1 vccd1 vccd1 _3577_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2528_ _2534_/A _4735_/A vssd1 vssd1 vccd1 vccd1 _2528_/Y sky130_fd_sc_hd__nand2_1
X_5247_ _5251_/CLK _5247_/D vssd1 vssd1 vccd1 vccd1 _5247_/Q sky130_fd_sc_hd__dfxtp_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_75_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5178_ _5181_/CLK _5178_/D vssd1 vssd1 vccd1 vccd1 _5178_/Q sky130_fd_sc_hd__dfxtp_1
X_4129_ _4294_/A _4129_/B _4144_/A vssd1 vssd1 vccd1 vccd1 _4133_/C sky130_fd_sc_hd__nor3_1
XFILLER_28_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3500_ _5223_/Q _3500_/B vssd1 vssd1 vccd1 vccd1 _3507_/B sky130_fd_sc_hd__nor2_1
X_4480_ _4387_/X _4477_/Y _4478_/X _4424_/X _4479_/Y vssd1 vssd1 vccd1 vccd1 _5034_/D
+ sky130_fd_sc_hd__o311a_1
X_3431_ _3611_/B _3608_/A vssd1 vssd1 vccd1 vccd1 _3431_/X sky130_fd_sc_hd__or2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3362_ _5116_/Q _3793_/B vssd1 vssd1 vccd1 vccd1 _3370_/B sky130_fd_sc_hd__or2_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _5201_/CLK _5101_/D vssd1 vssd1 vccd1 vccd1 _5101_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _3291_/X _3292_/Y _3272_/X vssd1 vssd1 vccd1 vccd1 _3293_/X sky130_fd_sc_hd__a21o_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _5068_/CLK _5032_/D vssd1 vssd1 vccd1 vccd1 _5032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4816_ _4816_/A _4826_/B vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4747_ _4745_/X _4746_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5009_/D sky130_fd_sc_hd__a21oi_1
XFILLER_31_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4678_ _4679_/A _4679_/B _4679_/C vssd1 vssd1 vccd1 vccd1 _4680_/B sky130_fd_sc_hd__a21oi_1
X_3629_ _5169_/Q _3580_/X _3627_/Y _3628_/X _3587_/X vssd1 vssd1 vccd1 vccd1 _5169_/D
+ sky130_fd_sc_hd__o221a_1
Xoutput49 _5165_/Q vssd1 vssd1 vccd1 vccd1 data_out[3] sky130_fd_sc_hd__buf_2
Xoutput27 _5174_/Q vssd1 vssd1 vccd1 vccd1 data_out[12] sky130_fd_sc_hd__buf_2
Xoutput38 _5184_/Q vssd1 vssd1 vccd1 vccd1 data_out[22] sky130_fd_sc_hd__buf_2
XFILLER_88_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3980_ _3980_/A vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__inv_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _2929_/X _2925_/A _2930_/X vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2862_ _2862_/A _2862_/B vssd1 vssd1 vccd1 vccd1 _2862_/Y sky130_fd_sc_hd__nand2_1
X_4601_ _4788_/A _4788_/B _4600_/Y vssd1 vssd1 vccd1 vccd1 _4777_/A sky130_fd_sc_hd__o21ai_1
X_2793_ _4772_/A vssd1 vssd1 vccd1 vccd1 _4115_/B sky130_fd_sc_hd__buf_4
X_4532_ _4987_/Q _5024_/Q _4530_/Y _4531_/X _4511_/X vssd1 vssd1 vccd1 vccd1 _5024_/D
+ sky130_fd_sc_hd__o221a_1
X_4463_ _4463_/A _4463_/B vssd1 vssd1 vccd1 vccd1 _4464_/A sky130_fd_sc_hd__or2_1
XFILLER_7_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3414_ _3414_/A _3414_/B vssd1 vssd1 vccd1 vccd1 _3627_/A sky130_fd_sc_hd__or2_1
X_4394_ _4387_/X _4390_/X _4392_/X _2808_/X _4393_/Y vssd1 vssd1 vccd1 vccd1 _5050_/D
+ sky130_fd_sc_hd__o311a_1
X_3345_ _3527_/B vssd1 vssd1 vccd1 vccd1 _3345_/Y sky130_fd_sc_hd__inv_2
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _3276_/A _3276_/B vssd1 vssd1 vccd1 vccd1 _3282_/A sky130_fd_sc_hd__and2_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ _5283_/CLK _5015_/D vssd1 vssd1 vccd1 vccd1 _5015_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3130_ _3208_/B _3130_/B vssd1 vssd1 vccd1 vccd1 _3212_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3061_ _3304_/A _3309_/A _3304_/B vssd1 vssd1 vccd1 vccd1 _3295_/A sky130_fd_sc_hd__a21oi_2
XFILLER_35_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3963_ _3995_/B _3995_/A vssd1 vssd1 vccd1 vccd1 _3964_/B sky130_fd_sc_hd__nor2_1
XFILLER_35_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2914_ _3259_/A vssd1 vssd1 vccd1 vccd1 _2914_/X sky130_fd_sc_hd__clkbuf_2
X_3894_ _4931_/A _4986_/Q vssd1 vssd1 vccd1 vccd1 _3897_/C sky130_fd_sc_hd__nand2_1
X_2845_ _5251_/Q _2814_/X _2842_/X _2844_/Y _2822_/X vssd1 vssd1 vccd1 vccd1 _5251_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_12_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4515_ _4987_/Q _5027_/Q _4469_/X _4514_/Y vssd1 vssd1 vccd1 vccd1 _5027_/D sky130_fd_sc_hd__o211a_1
X_2776_ _2766_/Y _2775_/Y _2702_/Y vssd1 vssd1 vccd1 vccd1 _2896_/A sky130_fd_sc_hd__o21bai_1
X_4446_ _4447_/A _4448_/A _4447_/B _4535_/A vssd1 vssd1 vccd1 vccd1 _4446_/X sky130_fd_sc_hd__a31o_1
X_4377_ _4378_/A _4378_/B _4383_/B _4378_/D vssd1 vssd1 vccd1 vccd1 _4377_/X sky130_fd_sc_hd__o22a_1
XFILLER_58_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3328_ _3331_/B _3327_/B _3312_/X vssd1 vssd1 vccd1 vccd1 _3328_/X sky130_fd_sc_hd__a21o_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3259_ _3259_/A vssd1 vssd1 vccd1 vccd1 _3259_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_54_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2630_ _2630_/A _2630_/B _2629_/Y vssd1 vssd1 vccd1 vccd1 _2783_/A sky130_fd_sc_hd__or3b_1
X_2561_ _5002_/Q vssd1 vssd1 vccd1 vccd1 _4782_/A sky130_fd_sc_hd__inv_2
X_2492_ _5020_/Q vssd1 vssd1 vccd1 vccd1 hold6/A sky130_fd_sc_hd__inv_2
X_4300_ _5073_/Q _5041_/Q vssd1 vssd1 vccd1 vccd1 _4434_/B sky130_fd_sc_hd__nand2_1
X_5280_ _5282_/CLK _5280_/D vssd1 vssd1 vccd1 vccd1 _5280_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4231_ _4455_/A _4457_/B _4455_/B vssd1 vssd1 vccd1 vccd1 _4431_/A sky130_fd_sc_hd__o21bai_2
XFILLER_4_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4162_ _4711_/A _4247_/A _4162_/C vssd1 vssd1 vccd1 vccd1 _4166_/A sky130_fd_sc_hd__or3_1
X_4093_ _4093_/A _4093_/B vssd1 vssd1 vccd1 vccd1 _4093_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3113_ _3229_/B _3113_/B _3113_/C vssd1 vssd1 vccd1 vccd1 _3113_/X sky130_fd_sc_hd__or3_1
X_3044_ _3044_/A _3076_/A vssd1 vssd1 vccd1 vccd1 _3265_/A sky130_fd_sc_hd__nand2_1
XFILLER_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4995_ _5265_/CLK _4995_/D vssd1 vssd1 vccd1 vccd1 _4995_/Q sky130_fd_sc_hd__dfxtp_1
X_3946_ _3945_/A _3945_/B _3945_/C vssd1 vssd1 vccd1 vccd1 _4002_/A sky130_fd_sc_hd__o21ai_1
XFILLER_11_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3877_ _3867_/X _4949_/X _3868_/X _3876_/Y vssd1 vssd1 vccd1 vccd1 _5090_/D sky130_fd_sc_hd__o211a_1
X_2828_ _2837_/C _2828_/B _2828_/C vssd1 vssd1 vccd1 vccd1 _2828_/X sky130_fd_sc_hd__and3_1
X_2759_ _5289_/Q _4940_/B vssd1 vssd1 vccd1 vccd1 _2761_/B sky130_fd_sc_hd__nor2_1
X_4429_ _4987_/Q _5043_/Q _3907_/X _4428_/Y vssd1 vssd1 vccd1 vccd1 _5043_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 _4984_/CLK sky130_fd_sc_hd__clkbuf_2
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3800_ _3810_/A _3800_/B vssd1 vssd1 vccd1 vccd1 _3800_/Y sky130_fd_sc_hd__nand2_1
X_4780_ _4781_/A _4781_/C _4781_/B vssd1 vssd1 vccd1 vccd1 _4780_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_20_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3731_ _5139_/Q _3725_/X _3722_/X _3730_/Y vssd1 vssd1 vccd1 vccd1 _5139_/D sky130_fd_sc_hd__o211a_1
X_3662_ _3837_/B _5099_/Q vssd1 vssd1 vccd1 vccd1 _3663_/A sky130_fd_sc_hd__nand2_1
X_3593_ _3593_/A _3593_/B vssd1 vssd1 vccd1 vccd1 _3597_/A sky130_fd_sc_hd__nor2_1
X_2613_ _5287_/Q hold6/A vssd1 vssd1 vccd1 vccd1 _2804_/A sky130_fd_sc_hd__nor2_1
X_2544_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_87_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5263_ _5263_/CLK _5263_/D vssd1 vssd1 vccd1 vccd1 _5263_/Q sky130_fd_sc_hd__dfxtp_1
X_4214_ _4413_/A _4415_/A vssd1 vssd1 vccd1 vccd1 _4324_/A sky130_fd_sc_hd__nor2_1
X_5194_ _5227_/CLK _5194_/D vssd1 vssd1 vccd1 vccd1 _5194_/Q sky130_fd_sc_hd__dfxtp_2
X_4145_ _4142_/Y _4235_/A _4144_/Y vssd1 vssd1 vccd1 vccd1 _5066_/D sky130_fd_sc_hd__a21oi_1
XFILLER_68_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4076_ _4074_/X _4075_/X _4057_/X _4058_/X _5083_/Q vssd1 vssd1 vccd1 vccd1 _4078_/B
+ sky130_fd_sc_hd__a41oi_1
XFILLER_70_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3027_ _5147_/Q _3709_/B vssd1 vssd1 vccd1 vccd1 _3111_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4978_ _5090_/CLK _4978_/D vssd1 vssd1 vccd1 vccd1 _4978_/Q sky130_fd_sc_hd__dfxtp_1
X_3929_ _4058_/A vssd1 vssd1 vccd1 vccd1 _4077_/B sky130_fd_sc_hd__inv_2
XFILLER_3_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4901_ _5091_/Q _4901_/B vssd1 vssd1 vccd1 vccd1 _4903_/A sky130_fd_sc_hd__nor2_1
X_4832_ _4992_/Q _4987_/Q _4830_/Y _4831_/X _4772_/X vssd1 vssd1 vccd1 vccd1 _4992_/D
+ sky130_fd_sc_hd__o221a_1
X_4763_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4763_/Y sky130_fd_sc_hd__xnor2_1
X_4694_ _4693_/B _4693_/A _4436_/X vssd1 vssd1 vccd1 vccd1 _4694_/X sky130_fd_sc_hd__a21o_1
X_3714_ _3716_/A _3714_/B vssd1 vssd1 vccd1 vccd1 _3714_/Y sky130_fd_sc_hd__nand2_1
X_3645_ _3645_/A _3645_/B _3649_/A vssd1 vssd1 vccd1 vccd1 _3645_/X sky130_fd_sc_hd__and3_1
XFILLER_20_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3576_ _3576_/A _3576_/B vssd1 vssd1 vccd1 vccd1 _3576_/Y sky130_fd_sc_hd__nand2_1
X_2527_ _5011_/Q vssd1 vssd1 vccd1 vccd1 _4735_/A sky130_fd_sc_hd__clkinv_2
X_5246_ _5289_/CLK _5246_/D vssd1 vssd1 vccd1 vccd1 _5246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold16 hold16/A vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_68_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5177_ _5213_/CLK _5177_/D vssd1 vssd1 vccd1 vccd1 _5177_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4128_ _4141_/A _4141_/B _4134_/C vssd1 vssd1 vccd1 vccd1 _4144_/A sky130_fd_sc_hd__nand3_2
XFILLER_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4059_ _4151_/A _4057_/X _4058_/X _3931_/A _5086_/Q vssd1 vssd1 vccd1 vccd1 _4060_/C
+ sky130_fd_sc_hd__a41oi_1
XFILLER_56_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3430_ _3430_/A vssd1 vssd1 vccd1 vccd1 _3608_/A sky130_fd_sc_hd__inv_2
X_3361_ _3562_/A vssd1 vssd1 vccd1 vccd1 _3453_/A sky130_fd_sc_hd__inv_2
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _5201_/CLK _5100_/D vssd1 vssd1 vccd1 vccd1 _5100_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _5068_/CLK _5031_/D vssd1 vssd1 vccd1 vccd1 _5031_/Q sky130_fd_sc_hd__dfxtp_1
X_3292_ _3292_/A _3292_/B vssd1 vssd1 vccd1 vccd1 _3292_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4815_ _4995_/Q _4987_/Q _4784_/X _4814_/X vssd1 vssd1 vccd1 vccd1 _4995_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4746_ _4746_/A _5009_/Q vssd1 vssd1 vccd1 vccd1 _4746_/Y sky130_fd_sc_hd__nand2_1
X_4677_ hold4/A _5054_/Q vssd1 vssd1 vccd1 vccd1 _4679_/C sky130_fd_sc_hd__xnor2_1
X_3628_ _3627_/B _3627_/A _3598_/X vssd1 vssd1 vccd1 vccd1 _3628_/X sky130_fd_sc_hd__a21o_1
Xoutput28 _5175_/Q vssd1 vssd1 vccd1 vccd1 data_out[13] sky130_fd_sc_hd__buf_2
Xoutput39 _5185_/Q vssd1 vssd1 vccd1 vccd1 data_out[23] sky130_fd_sc_hd__buf_2
X_3559_ _5182_/Q _3537_/X _3303_/X _3558_/X vssd1 vssd1 vccd1 vccd1 _5182_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5229_ _5259_/CLK _5229_/D vssd1 vssd1 vccd1 vccd1 _5229_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _3577_/A vssd1 vssd1 vccd1 vccd1 _2930_/X sky130_fd_sc_hd__buf_2
XFILLER_30_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _2858_/Y _2859_/X _2860_/X vssd1 vssd1 vccd1 vccd1 _5249_/D sky130_fd_sc_hd__o21a_1
X_4600_ _4793_/A _4790_/A vssd1 vssd1 vccd1 vccd1 _4600_/Y sky130_fd_sc_hd__nor2_1
X_2792_ _4103_/A vssd1 vssd1 vccd1 vccd1 _4772_/A sky130_fd_sc_hd__clkbuf_2
X_4531_ _4529_/X _5055_/Q _5023_/Q _4181_/X vssd1 vssd1 vccd1 vccd1 _4531_/X sky130_fd_sc_hd__a31o_1
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4462_ _4987_/Q _5037_/Q _3907_/X _4461_/X vssd1 vssd1 vccd1 vccd1 _5037_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3413_ _3822_/B _5105_/Q vssd1 vssd1 vccd1 vccd1 _3414_/B sky130_fd_sc_hd__and2_1
X_4393_ _4479_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4393_/Y sky130_fd_sc_hd__nand2_1
X_3344_ _3355_/B _3344_/B vssd1 vssd1 vccd1 vccd1 _3527_/B sky130_fd_sc_hd__nand2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _3275_/A vssd1 vssd1 vccd1 vccd1 _3279_/A sky130_fd_sc_hd__inv_2
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5014_ _5045_/CLK _5014_/D vssd1 vssd1 vccd1 vccd1 _5014_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4729_ _4726_/Y _4728_/X _2839_/X vssd1 vssd1 vccd1 vccd1 _5013_/D sky130_fd_sc_hd__o21a_1
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3060_ _3299_/B _3060_/B vssd1 vssd1 vccd1 vccd1 _3304_/B sky130_fd_sc_hd__nand2_1
X_3962_ _3996_/A _3964_/A _3995_/A _3995_/B vssd1 vssd1 vccd1 vccd1 _3975_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_16_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2913_ _2911_/B _2911_/A _2912_/X vssd1 vssd1 vccd1 vccd1 _2913_/X sky130_fd_sc_hd__a21o_1
X_3893_ _5095_/Q _4882_/B _5088_/Q _3891_/Y _3892_/X vssd1 vssd1 vccd1 vccd1 _3897_/A
+ sky130_fd_sc_hd__o221a_1
X_2844_ _2844_/A _2844_/B vssd1 vssd1 vccd1 vccd1 _2844_/Y sky130_fd_sc_hd__nor2_1
X_4514_ _4513_/Y _4507_/X _4987_/Q vssd1 vssd1 vccd1 vccd1 _4514_/Y sky130_fd_sc_hd__o21ai_1
X_2775_ _2922_/A _2922_/B _2693_/Y vssd1 vssd1 vccd1 vccd1 _2775_/Y sky130_fd_sc_hd__a21oi_1
X_4445_ _4445_/A _4445_/B vssd1 vssd1 vccd1 vccd1 _4448_/A sky130_fd_sc_hd__nor2_1
X_4376_ _5084_/Q _5052_/Q vssd1 vssd1 vccd1 vccd1 _4378_/B sky130_fd_sc_hd__nor2_1
X_3327_ _3331_/B _3327_/B vssd1 vssd1 vccd1 vccd1 _3327_/Y sky130_fd_sc_hd__nor2_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3258_ _3257_/B _3257_/A _3244_/X vssd1 vssd1 vccd1 vccd1 _3258_/X sky130_fd_sc_hd__a21o_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3189_ _3187_/Y _3188_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5220_/D sky130_fd_sc_hd__a21oi_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2560_ _5270_/Q _2544_/X _2547_/X _2559_/Y vssd1 vssd1 vccd1 vccd1 _5270_/D sky130_fd_sc_hd__o211a_1
X_2491_ _5288_/Q _2481_/X _2485_/X _2490_/Y vssd1 vssd1 vccd1 vccd1 _5288_/D sky130_fd_sc_hd__o211a_1
X_4230_ _5070_/Q _5038_/Q vssd1 vssd1 vccd1 vccd1 _4455_/B sky130_fd_sc_hd__and2_1
X_4161_ _5059_/Q vssd1 vssd1 vccd1 vccd1 _4247_/A sky130_fd_sc_hd__inv_2
XFILLER_67_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4092_ _4110_/A _4092_/B vssd1 vssd1 vccd1 vccd1 _4099_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3112_ _3236_/A _3233_/A vssd1 vssd1 vccd1 vccd1 _3113_/C sky130_fd_sc_hd__nand2_1
X_3043_ _5139_/Q _3730_/B vssd1 vssd1 vccd1 vccd1 _3076_/A sky130_fd_sc_hd__or2_1
XFILLER_55_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _4996_/CLK _4994_/D vssd1 vssd1 vccd1 vccd1 _4994_/Q sky130_fd_sc_hd__dfxtp_2
X_3945_ _3945_/A _3945_/B _3945_/C vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__or3_1
XFILLER_23_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3876_ _3879_/A _3876_/B vssd1 vssd1 vccd1 vccd1 _3876_/Y sky130_fd_sc_hd__nand2_1
X_2827_ _2837_/C _2828_/C _2828_/B vssd1 vssd1 vccd1 vccd1 _2827_/Y sky130_fd_sc_hd__a21oi_1
X_2758_ hold4/X vssd1 vssd1 vccd1 vccd1 _4940_/B sky130_fd_sc_hd__inv_2
X_4428_ _4421_/B _4427_/X _4987_/Q vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__o21ai_1
X_2689_ _2689_/A vssd1 vssd1 vccd1 vccd1 _2929_/A sky130_fd_sc_hd__inv_2
X_4359_ _4359_/A _4671_/B vssd1 vssd1 vccd1 vccd1 _4378_/A sky130_fd_sc_hd__nor2_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3730_ _3730_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _3730_/Y sky130_fd_sc_hd__nand2_1
X_3661_ _3839_/B _5098_/Q vssd1 vssd1 vccd1 vccd1 _3668_/B sky130_fd_sc_hd__nand2_1
XFILLER_70_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3592_ _5176_/Q _3537_/X _3589_/X _3591_/X vssd1 vssd1 vccd1 vccd1 _5176_/D sky130_fd_sc_hd__o211a_1
X_2612_ _5258_/Q _2584_/X _2609_/X _2611_/Y vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__o211a_1
X_2543_ _5274_/Q _2525_/X _2526_/X _2542_/Y vssd1 vssd1 vccd1 vccd1 _5274_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5262_ _5263_/CLK hold16/X vssd1 vssd1 vccd1 vccd1 _5262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4213_ _4213_/A vssd1 vssd1 vccd1 vccd1 _4415_/A sky130_fd_sc_hd__inv_2
X_5193_ _5193_/CLK _5193_/D vssd1 vssd1 vccd1 vccd1 _5193_/Q sky130_fd_sc_hd__dfxtp_1
X_4144_ _4144_/A _4144_/B vssd1 vssd1 vccd1 vccd1 _4144_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4075_ _4141_/B vssd1 vssd1 vccd1 vccd1 _4075_/X sky130_fd_sc_hd__clkbuf_2
X_3026_ _5243_/Q vssd1 vssd1 vccd1 vccd1 _3709_/B sky130_fd_sc_hd__inv_2
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ _5137_/CLK _4977_/D vssd1 vssd1 vccd1 vccd1 _4977_/Q sky130_fd_sc_hd__dfxtp_1
X_3928_ _4063_/C _4087_/B vssd1 vssd1 vccd1 vccd1 _4058_/A sky130_fd_sc_hd__nor2_1
X_3859_ _3844_/X _4944_/X _3845_/X _3858_/Y vssd1 vssd1 vccd1 vccd1 _5095_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4900_ _4900_/A vssd1 vssd1 vccd1 vccd1 _4900_/X sky130_fd_sc_hd__clkbuf_1
X_4831_ _4830_/B _4830_/A _4181_/X vssd1 vssd1 vccd1 vccd1 _4831_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_1_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4762_ _4516_/X _4758_/Y _4759_/X _4760_/X _4761_/Y vssd1 vssd1 vccd1 vccd1 _5006_/D
+ sky130_fd_sc_hd__o311a_1
X_3713_ _5146_/Q _3711_/X _3708_/X _3712_/Y vssd1 vssd1 vccd1 vccd1 _5146_/D sky130_fd_sc_hd__o211a_1
X_4693_ _4693_/A _4693_/B vssd1 vssd1 vccd1 vccd1 _4693_/Y sky130_fd_sc_hd__nor2_1
X_3644_ _3644_/A vssd1 vssd1 vccd1 vccd1 _3644_/X sky130_fd_sc_hd__buf_4
X_3575_ _5179_/Q _3512_/X _3572_/X _3574_/Y _3518_/X vssd1 vssd1 vccd1 vccd1 _5179_/D
+ sky130_fd_sc_hd__o221a_1
X_2526_ _4853_/A vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5245_ _5287_/CLK _5245_/D vssd1 vssd1 vccd1 vccd1 _5245_/Q sky130_fd_sc_hd__dfxtp_1
Xhold17 hold17/A vssd1 vssd1 vccd1 vccd1 hold17/X sky130_fd_sc_hd__clkdlybuf4s50_1
X_5176_ _5181_/CLK _5176_/D vssd1 vssd1 vccd1 vccd1 _5176_/Q sky130_fd_sc_hd__dfxtp_1
X_4127_ _4127_/A vssd1 vssd1 vccd1 vccd1 _4134_/C sky130_fd_sc_hd__inv_2
XFILLER_68_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4058_ _4058_/A vssd1 vssd1 vccd1 vccd1 _4058_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_45_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3009_ hold17/A _5157_/Q vssd1 vssd1 vccd1 vccd1 _3015_/A sky130_fd_sc_hd__and2_1
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3360_ _3371_/A _3370_/A vssd1 vssd1 vccd1 vccd1 _3562_/A sky130_fd_sc_hd__nor2_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _5265_/CLK _5030_/D vssd1 vssd1 vccd1 vccd1 _5030_/Q sky130_fd_sc_hd__dfxtp_1
X_3291_ _3292_/B _3292_/A vssd1 vssd1 vccd1 vccd1 _3291_/X sky130_fd_sc_hd__or2_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4814_ _4813_/X _4810_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _4814_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4745_ _4745_/A _4745_/B _4739_/Y vssd1 vssd1 vccd1 vccd1 _4745_/X sky130_fd_sc_hd__or3b_1
X_4676_ _4674_/B _4682_/B _4987_/Q vssd1 vssd1 vccd1 vccd1 _4679_/A sky130_fd_sc_hd__o21ai_1
X_3627_ _3627_/A _3627_/B vssd1 vssd1 vccd1 vccd1 _3627_/Y sky130_fd_sc_hd__nor2_1
Xoutput29 _5176_/Q vssd1 vssd1 vccd1 vccd1 data_out[14] sky130_fd_sc_hd__buf_2
X_3558_ _3557_/X _3544_/Y _3272_/X vssd1 vssd1 vccd1 vccd1 _3558_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2509_ _2516_/A _4650_/A vssd1 vssd1 vccd1 vccd1 _2509_/Y sky130_fd_sc_hd__nand2_1
X_3489_ _3764_/B _5127_/Q _3485_/Y _3488_/Y vssd1 vssd1 vccd1 vccd1 _3489_/Y sky130_fd_sc_hd__a22oi_1
X_5228_ _5228_/CLK _5228_/D vssd1 vssd1 vccd1 vccd1 _5228_/Q sky130_fd_sc_hd__dfxtp_1
X_5159_ _5263_/CLK _5159_/D vssd1 vssd1 vccd1 vccd1 _5159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5230_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_44_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_27_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5263_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_46_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2860_ _5249_/Q _3528_/B _4849_/A vssd1 vssd1 vccd1 vccd1 _2860_/X sky130_fd_sc_hd__o21a_1
XFILLER_62_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2791_ _2791_/A vssd1 vssd1 vccd1 vccd1 _4103_/A sky130_fd_sc_hd__clkbuf_4
X_4530_ _5055_/Q _5023_/Q _4529_/X vssd1 vssd1 vccd1 vccd1 _4530_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_7_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4461_ _4457_/A _4460_/Y _4407_/X vssd1 vssd1 vccd1 vccd1 _4461_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3412_ _5105_/Q _3822_/B vssd1 vssd1 vccd1 vccd1 _3414_/A sky130_fd_sc_hd__nor2_1
X_4392_ _4338_/A _4397_/C _4353_/C vssd1 vssd1 vccd1 vccd1 _4392_/X sky130_fd_sc_hd__o21a_1
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3343_ _3771_/B _5124_/Q vssd1 vssd1 vccd1 vccd1 _3344_/B sky130_fd_sc_hd__nand2_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _5204_/Q _3261_/X _3247_/X _3273_/X vssd1 vssd1 vccd1 vccd1 _5204_/D sky130_fd_sc_hd__o211a_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _5045_/CLK _5013_/D vssd1 vssd1 vccd1 vccd1 _5013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _5070_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_34_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2989_ _2983_/Y _2988_/Y _2839_/X vssd1 vssd1 vccd1 vccd1 _5227_/D sky130_fd_sc_hd__o21a_1
X_4728_ _4728_/A _4987_/Q _4728_/C vssd1 vssd1 vccd1 vccd1 _4728_/X sky130_fd_sc_hd__and3_1
X_4659_ _4702_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4660_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3961_ _4958_/Q _3961_/B vssd1 vssd1 vccd1 vccd1 _3995_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2912_ _3598_/A vssd1 vssd1 vccd1 vccd1 _2912_/X sky130_fd_sc_hd__buf_2
X_3892_ _4980_/Q _3876_/B _4925_/B _4985_/Q vssd1 vssd1 vccd1 vccd1 _3892_/X sky130_fd_sc_hd__o22a_1
X_2843_ _2843_/A _2843_/B vssd1 vssd1 vccd1 vccd1 _2844_/B sky130_fd_sc_hd__and2_1
X_2774_ _2933_/A _2933_/B _2774_/C vssd1 vssd1 vccd1 vccd1 _2922_/A sky130_fd_sc_hd__nand3_1
X_4513_ _4507_/A _4520_/C _4507_/C vssd1 vssd1 vccd1 vccd1 _4513_/Y sky130_fd_sc_hd__a21oi_1
X_4444_ _4450_/B _4450_/A vssd1 vssd1 vccd1 vccd1 _4447_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_7_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5283_/CLK sky130_fd_sc_hd__clkbuf_16
X_4375_ _4372_/Y _4374_/X _2839_/X vssd1 vssd1 vccd1 vccd1 _5053_/D sky130_fd_sc_hd__o21a_1
X_3326_ _3326_/A _3326_/B vssd1 vssd1 vccd1 vccd1 _3327_/B sky130_fd_sc_hd__nand2_1
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _3257_/A _3257_/B vssd1 vssd1 vccd1 vccd1 _3257_/Y sky130_fd_sc_hd__nor2_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3188_ _3505_/A _5220_/Q vssd1 vssd1 vccd1 vccd1 _3188_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2490_ _2496_/A _4537_/A vssd1 vssd1 vccd1 vccd1 _2490_/Y sky130_fd_sc_hd__nand2_1
X_4160_ _5060_/Q vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__inv_2
XFILLER_67_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3111_ _3111_/A _3111_/B vssd1 vssd1 vccd1 vccd1 _3233_/A sky130_fd_sc_hd__nor2_1
X_4091_ _4093_/A _4332_/A _4090_/Y vssd1 vssd1 vccd1 vccd1 _5080_/D sky130_fd_sc_hd__a21oi_1
X_3042_ _3733_/B _5138_/Q _3076_/B vssd1 vssd1 vccd1 vccd1 _3044_/A sky130_fd_sc_hd__or3b_1
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4993_ _4996_/CLK _4993_/D vssd1 vssd1 vccd1 vccd1 _4993_/Q sky130_fd_sc_hd__dfxtp_1
X_3944_ _3944_/A _3944_/B vssd1 vssd1 vccd1 vccd1 _3945_/C sky130_fd_sc_hd__nor2_1
X_3875_ _5090_/Q vssd1 vssd1 vccd1 vccd1 _3876_/B sky130_fd_sc_hd__inv_2
X_2826_ _2835_/B _2835_/C _2835_/A vssd1 vssd1 vccd1 vccd1 _2837_/C sky130_fd_sc_hd__o21ai_1
X_2757_ _5288_/Q _4537_/A vssd1 vssd1 vccd1 vccd1 _2761_/A sky130_fd_sc_hd__nor2_1
X_2688_ _2925_/B _2688_/B vssd1 vssd1 vccd1 vccd1 _2689_/A sky130_fd_sc_hd__nand2_1
X_4427_ _4427_/A _4427_/B _4427_/C vssd1 vssd1 vccd1 vccd1 _4427_/X sky130_fd_sc_hd__and3_1
X_4358_ _5052_/Q vssd1 vssd1 vccd1 vccd1 _4671_/B sky130_fd_sc_hd__inv_2
XFILLER_58_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4289_ _4289_/A _4289_/B vssd1 vssd1 vccd1 vccd1 _4290_/A sky130_fd_sc_hd__nor2_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _3309_/A _3309_/B vssd1 vssd1 vccd1 vccd1 _3311_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _5194_/Q vssd1 vssd1 vccd1 vccd1 _3839_/B sky130_fd_sc_hd__inv_2
X_3591_ _3585_/A _3590_/Y _3577_/X vssd1 vssd1 vccd1 vccd1 _3591_/X sky130_fd_sc_hd__a21o_1
X_2611_ _3676_/A _2990_/B vssd1 vssd1 vccd1 vccd1 _2611_/Y sky130_fd_sc_hd__nand2_1
X_2542_ _2555_/A _4754_/A vssd1 vssd1 vccd1 vccd1 _2542_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5261_ _5263_/CLK _5261_/D vssd1 vssd1 vccd1 vccd1 _5261_/Q sky130_fd_sc_hd__dfxtp_1
X_4212_ _4212_/A _4212_/B vssd1 vssd1 vccd1 vccd1 _4213_/A sky130_fd_sc_hd__nor2_1
X_5192_ _5193_/CLK _5192_/D vssd1 vssd1 vccd1 vccd1 _5192_/Q sky130_fd_sc_hd__dfxtp_1
X_4143_ _5066_/Q vssd1 vssd1 vccd1 vccd1 _4235_/A sky130_fd_sc_hd__inv_2
X_4074_ _4141_/A vssd1 vssd1 vccd1 vccd1 _4074_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3025_ _3229_/B _3113_/B vssd1 vssd1 vccd1 vccd1 _3025_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4976_ _5137_/CLK _4976_/D vssd1 vssd1 vccd1 vccd1 _4976_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3927_ _4092_/B vssd1 vssd1 vccd1 vccd1 _4087_/B sky130_fd_sc_hd__inv_2
X_3858_ _3861_/A _4925_/B vssd1 vssd1 vccd1 vccd1 _3858_/Y sky130_fd_sc_hd__nand2_1
X_3789_ _3802_/A vssd1 vssd1 vccd1 vccd1 _3789_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2809_ _2809_/A vssd1 vssd1 vccd1 vccd1 _3238_/A sky130_fd_sc_hd__buf_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4830_ _4830_/A _4830_/B vssd1 vssd1 vccd1 vccd1 _4830_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4761_ _4761_/A _4794_/B vssd1 vssd1 vccd1 vccd1 _4761_/Y sky130_fd_sc_hd__nand2_1
X_4692_ _4692_/A _4692_/B vssd1 vssd1 vccd1 vccd1 _4693_/B sky130_fd_sc_hd__nand2_1
X_3712_ _3716_/A _3712_/B vssd1 vssd1 vccd1 vccd1 _3712_/Y sky130_fd_sc_hd__nand2_1
X_3643_ _5167_/Q _3634_/X _3638_/X _3641_/Y _3642_/X vssd1 vssd1 vccd1 vccd1 _5167_/D
+ sky130_fd_sc_hd__o221a_1
X_3574_ _3574_/A _3574_/B vssd1 vssd1 vccd1 vccd1 _3574_/Y sky130_fd_sc_hd__nor2_1
X_2525_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2525_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5244_ _5254_/CLK _5244_/D vssd1 vssd1 vccd1 vccd1 _5244_/Q sky130_fd_sc_hd__dfxtp_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5175_ _5209_/CLK _5175_/D vssd1 vssd1 vccd1 vccd1 _5175_/Q sky130_fd_sc_hd__dfxtp_1
X_4126_ _4126_/A _4151_/B vssd1 vssd1 vccd1 vccd1 _4127_/A sky130_fd_sc_hd__nand2_1
XFILLER_56_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4057_ _4068_/A vssd1 vssd1 vccd1 vccd1 _4057_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_28_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3008_ _5157_/Q hold17/A vssd1 vssd1 vccd1 vccd1 _3010_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4959_ _4964_/CLK _4959_/D vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__dfxtp_1
XFILLER_79_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _5201_/Q _3252_/X _3288_/Y _3289_/X _3259_/X vssd1 vssd1 vccd1 vccd1 _5201_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4813_ _4813_/A _4813_/B vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__or2_1
X_4744_ _4744_/A _4744_/B vssd1 vssd1 vccd1 vccd1 _4745_/B sky130_fd_sc_hd__nor2_1
X_4675_ _4681_/A _4681_/C _4681_/B vssd1 vssd1 vccd1 vccd1 _4682_/B sky130_fd_sc_hd__a21oi_1
X_3626_ _3626_/A _3626_/B vssd1 vssd1 vccd1 vccd1 _3627_/B sky130_fd_sc_hd__nand2_1
X_3557_ _3557_/A _3557_/B vssd1 vssd1 vccd1 vccd1 _3557_/X sky130_fd_sc_hd__or2_1
X_2508_ _5016_/Q vssd1 vssd1 vccd1 vccd1 _4650_/A sky130_fd_sc_hd__inv_2
XFILLER_88_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3488_ _3514_/A vssd1 vssd1 vccd1 vccd1 _3488_/Y sky130_fd_sc_hd__inv_2
X_5227_ _5227_/CLK _5227_/D vssd1 vssd1 vccd1 vccd1 _5227_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _5259_/CLK _5158_/D vssd1 vssd1 vccd1 vccd1 _5158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4109_ _4111_/A _4216_/A _4108_/Y vssd1 vssd1 vccd1 vccd1 _5076_/D sky130_fd_sc_hd__a21oi_1
X_5089_ _5090_/CLK _5089_/D vssd1 vssd1 vccd1 vccd1 _5089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_2_0_0_clk clkbuf_2_1_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_clk/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2790_ _2978_/A vssd1 vssd1 vccd1 vccd1 _3668_/A sky130_fd_sc_hd__buf_4
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _4460_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _4460_/Y sky130_fd_sc_hd__nand2_1
X_4391_ _4396_/B _4391_/B vssd1 vssd1 vccd1 vccd1 _4397_/C sky130_fd_sc_hd__nor2_1
X_3411_ _5201_/Q vssd1 vssd1 vccd1 vccd1 _3822_/B sky130_fd_sc_hd__inv_2
X_3342_ _5124_/Q _3771_/B vssd1 vssd1 vccd1 vccd1 _3355_/B sky130_fd_sc_hd__or2_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3273_ _3267_/A _3271_/Y _3272_/X vssd1 vssd1 vccd1 vccd1 _3273_/X sky130_fd_sc_hd__a21o_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ _5281_/CLK _5012_/D vssd1 vssd1 vccd1 vccd1 _5012_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2988_ _2991_/B _2986_/X _2987_/Y vssd1 vssd1 vccd1 vccd1 _2988_/Y sky130_fd_sc_hd__a21oi_1
X_4727_ _4727_/A _4727_/B vssd1 vssd1 vccd1 vccd1 _4728_/C sky130_fd_sc_hd__nand2_1
X_4658_ _5018_/Q _5050_/Q vssd1 vssd1 vccd1 vccd1 _4666_/A sky130_fd_sc_hd__nor2_1
X_3609_ _3608_/B _3608_/A _3598_/X vssd1 vssd1 vccd1 vccd1 _3609_/X sky130_fd_sc_hd__a21o_1
XFILLER_1_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4589_ _4589_/A _4589_/B vssd1 vssd1 vccd1 vccd1 _4590_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3960_ _3961_/B _4958_/Q vssd1 vssd1 vccd1 vccd1 _3995_/A sky130_fd_sc_hd__and2_1
XFILLER_35_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2911_ _2911_/A _2911_/B vssd1 vssd1 vccd1 vccd1 _2911_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3891_ _4978_/Q vssd1 vssd1 vccd1 vccd1 _3891_/Y sky130_fd_sc_hd__inv_2
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2842_ _2843_/A _2844_/A _2843_/B _2803_/A vssd1 vssd1 vccd1 vccd1 _2842_/X sky130_fd_sc_hd__a31o_1
X_2773_ _2773_/A vssd1 vssd1 vccd1 vccd1 _2774_/C sky130_fd_sc_hd__inv_2
X_4512_ _4987_/Q _5028_/Q _4509_/Y _4510_/X _4511_/X vssd1 vssd1 vccd1 vccd1 _5028_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_7_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4443_ _4441_/X _4442_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5041_/D sky130_fd_sc_hd__a21oi_1
X_4374_ _4378_/A _4373_/Y _4987_/Q _4368_/B vssd1 vssd1 vccd1 vccd1 _4374_/X sky130_fd_sc_hd__o211a_1
X_3325_ _3754_/B _5131_/Q vssd1 vssd1 vccd1 vccd1 _3326_/A sky130_fd_sc_hd__nand2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3256_ _3723_/B _5142_/Q _3255_/X vssd1 vssd1 vccd1 vccd1 _3257_/B sky130_fd_sc_hd__o21a_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3187_ _3187_/A _3504_/C _3187_/C vssd1 vssd1 vccd1 vccd1 _3187_/Y sky130_fd_sc_hd__nand3_1
XFILLER_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3110_ _3110_/A _3110_/B vssd1 vssd1 vccd1 vccd1 _3236_/A sky130_fd_sc_hd__nor2_1
X_4090_ _4081_/B _4065_/C _4093_/B vssd1 vssd1 vccd1 vccd1 _4090_/Y sky130_fd_sc_hd__o21ai_1
X_3041_ _3730_/B _5139_/Q vssd1 vssd1 vccd1 vccd1 _3076_/B sky130_fd_sc_hd__nand2_1
XFILLER_36_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4992_ _4996_/CLK _4992_/D vssd1 vssd1 vccd1 vccd1 _4992_/Q sky130_fd_sc_hd__dfxtp_2
X_3943_ _4962_/Q hold19/A vssd1 vssd1 vccd1 vccd1 _3944_/B sky130_fd_sc_hd__and2_1
X_3874_ _3867_/X _4948_/X _3868_/X _3873_/Y vssd1 vssd1 vccd1 vccd1 _5091_/D sky130_fd_sc_hd__o211a_1
X_2825_ _2841_/A _2825_/B vssd1 vssd1 vccd1 vccd1 _2835_/C sky130_fd_sc_hd__and2_1
X_2756_ _2804_/A _2752_/Y _2755_/Y vssd1 vssd1 vccd1 vccd1 _2798_/A sky130_fd_sc_hd__o21ai_1
X_2687_ _4603_/A _5268_/Q vssd1 vssd1 vccd1 vccd1 _2688_/B sky130_fd_sc_hd__nand2_1
X_4426_ _4387_/X _4422_/Y _4423_/X _4424_/X _4425_/Y vssd1 vssd1 vccd1 vccd1 _5044_/D
+ sky130_fd_sc_hd__o311a_1
X_4357_ _5084_/Q _5052_/Q _4383_/B _4378_/D vssd1 vssd1 vccd1 vccd1 _4373_/A sky130_fd_sc_hd__o22ai_2
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ _4288_/A _4612_/B vssd1 vssd1 vccd1 vccd1 _4289_/B sky130_fd_sc_hd__nor2_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3308_ _3747_/B _5133_/Q vssd1 vssd1 vccd1 vccd1 _3309_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _2803_/X _3236_/Y _2962_/X _3238_/Y vssd1 vssd1 vccd1 vccd1 _5210_/D sky130_fd_sc_hd__o211a_1
XFILLER_73_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3590_ _3590_/A _3590_/B vssd1 vssd1 vccd1 vccd1 _3590_/Y sky130_fd_sc_hd__nand2_1
X_2610_ _4991_/Q vssd1 vssd1 vccd1 vccd1 _2990_/B sky130_fd_sc_hd__inv_2
X_2541_ _4629_/A vssd1 vssd1 vccd1 vccd1 _4754_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5260_ _5263_/CLK hold10/X vssd1 vssd1 vccd1 vccd1 _5260_/Q sky130_fd_sc_hd__dfxtp_1
X_4211_ _4211_/A _4211_/B vssd1 vssd1 vccd1 vccd1 _4413_/A sky130_fd_sc_hd__nand2_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5191_ _5193_/CLK _5191_/D vssd1 vssd1 vccd1 vccd1 _5191_/Q sky130_fd_sc_hd__dfxtp_1
X_4142_ _4146_/A _4142_/B vssd1 vssd1 vccd1 vccd1 _4142_/Y sky130_fd_sc_hd__nand2_1
X_4073_ _4073_/A _4073_/B vssd1 vssd1 vccd1 vccd1 _5084_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3024_ _3024_/A vssd1 vssd1 vccd1 vccd1 _3113_/B sky130_fd_sc_hd__inv_2
XFILLER_36_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4975_ _5201_/CLK _4975_/D vssd1 vssd1 vccd1 vccd1 _4975_/Q sky130_fd_sc_hd__dfxtp_1
X_3926_ _3926_/A _4096_/B vssd1 vssd1 vccd1 vccd1 _4092_/B sky130_fd_sc_hd__and2_1
X_3857_ _5095_/Q vssd1 vssd1 vccd1 vccd1 _4925_/B sky130_fd_sc_hd__inv_2
XFILLER_50_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2808_ _4784_/A vssd1 vssd1 vccd1 vccd1 _2808_/X sky130_fd_sc_hd__buf_2
X_3788_ _5118_/Q _3779_/X _3776_/X _3787_/Y vssd1 vssd1 vccd1 vccd1 _5118_/D sky130_fd_sc_hd__o211a_1
X_2739_ _2739_/A vssd1 vssd1 vccd1 vccd1 _2739_/Y sky130_fd_sc_hd__inv_2
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4409_ _4987_/Q _5047_/Q _3907_/X _4408_/X vssd1 vssd1 vccd1 vccd1 _5047_/D sky130_fd_sc_hd__o211a_1
XFILLER_86_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4760_ _4760_/A vssd1 vssd1 vccd1 vccd1 _4760_/X sky130_fd_sc_hd__buf_2
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4691_ _4691_/A vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__inv_2
X_3711_ _3725_/A vssd1 vssd1 vccd1 vccd1 _3711_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3642_ _4183_/A vssd1 vssd1 vccd1 vccd1 _3642_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3573_ _3573_/A _3573_/B vssd1 vssd1 vccd1 vccd1 _3574_/B sky130_fd_sc_hd__and2_1
X_2524_ _5279_/Q _2506_/X _2507_/X _2523_/Y vssd1 vssd1 vccd1 vccd1 hold2/A sky130_fd_sc_hd__o211a_1
X_5243_ _5251_/CLK _5243_/D vssd1 vssd1 vccd1 vccd1 _5243_/Q sky130_fd_sc_hd__dfxtp_1
Xhold19 hold19/A vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__clkdlybuf4s25_1
X_5174_ _5209_/CLK _5174_/D vssd1 vssd1 vccd1 vccd1 _5174_/Q sky130_fd_sc_hd__dfxtp_1
X_4125_ _4125_/A vssd1 vssd1 vccd1 vccd1 _4129_/B sky130_fd_sc_hd__inv_2
XFILLER_68_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _4163_/B vssd1 vssd1 vccd1 vccd1 _4151_/A sky130_fd_sc_hd__clkbuf_2
X_3007_ _3002_/Y _3142_/A _3143_/B vssd1 vssd1 vccd1 vccd1 _3186_/B sky130_fd_sc_hd__a21oi_1
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4958_ _4964_/CLK hold22/X vssd1 vssd1 vccd1 vccd1 _4958_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4889_ _5089_/Q _5088_/Q vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__nor2_1
X_3909_ _3886_/X _4951_/S _3907_/X _3908_/Y vssd1 vssd1 vccd1 vccd1 _5087_/D sky130_fd_sc_hd__o211a_1
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4812_ _3861_/A _4809_/Y _4810_/X _4760_/X _4811_/Y vssd1 vssd1 vccd1 vccd1 _4996_/D
+ sky130_fd_sc_hd__o311a_1
X_4743_ _5010_/Q _4987_/Q _4741_/Y _4742_/X _4713_/X vssd1 vssd1 vccd1 vccd1 _5010_/D
+ sky130_fd_sc_hd__o221a_1
X_4674_ _4674_/A _4674_/B vssd1 vssd1 vccd1 vccd1 _4681_/B sky130_fd_sc_hd__or2_1
X_3625_ _3824_/B _5104_/Q _3631_/A vssd1 vssd1 vccd1 vccd1 _3626_/A sky130_fd_sc_hd__a21o_1
X_3556_ _5183_/Q _3512_/X _3554_/Y _3555_/X _3518_/X vssd1 vssd1 vccd1 vccd1 _5183_/D
+ sky130_fd_sc_hd__o221a_1
X_2507_ _4853_/A vssd1 vssd1 vccd1 vccd1 _2507_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3487_ _5126_/Q _3767_/B vssd1 vssd1 vccd1 vccd1 _3514_/A sky130_fd_sc_hd__nor2_1
X_5226_ _5228_/CLK _5226_/D vssd1 vssd1 vccd1 vccd1 _5226_/Q sky130_fd_sc_hd__dfxtp_1
X_5157_ _5259_/CLK _5157_/D vssd1 vssd1 vccd1 vccd1 _5157_/Q sky130_fd_sc_hd__dfxtp_1
X_4108_ _4097_/A _4065_/C _4093_/B vssd1 vssd1 vccd1 vccd1 _4108_/Y sky130_fd_sc_hd__o21ai_1
X_5088_ _5090_/CLK _5088_/D vssd1 vssd1 vccd1 vccd1 _5088_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4039_ _5064_/Q vssd1 vssd1 vccd1 vccd1 _4272_/A sky130_fd_sc_hd__inv_2
XFILLER_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4390_ _4396_/B _4391_/B _4345_/A _4340_/A vssd1 vssd1 vccd1 vccd1 _4390_/X sky130_fd_sc_hd__o211a_1
X_3410_ _3626_/B _3410_/B vssd1 vssd1 vccd1 vccd1 _3631_/B sky130_fd_sc_hd__nand2_1
X_3341_ _5220_/Q vssd1 vssd1 vccd1 vccd1 _3771_/B sky130_fd_sc_hd__inv_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _3577_/A vssd1 vssd1 vccd1 vccd1 _3272_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5011_ _5283_/CLK _5011_/D vssd1 vssd1 vccd1 vccd1 _5011_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2987_ _2991_/B _2986_/X _3832_/A vssd1 vssd1 vccd1 vccd1 _2987_/Y sky130_fd_sc_hd__o21ai_1
X_4726_ _4987_/Q _4726_/B vssd1 vssd1 vccd1 vccd1 _4726_/Y sky130_fd_sc_hd__nor2_1
X_4657_ _4666_/B _4657_/B vssd1 vssd1 vccd1 vccd1 _4704_/B sky130_fd_sc_hd__nand2_1
X_3608_ _3608_/A _3608_/B vssd1 vssd1 vccd1 vccd1 _3608_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4588_ _4573_/A _4810_/C _4573_/B vssd1 vssd1 vccd1 vccd1 _4797_/B sky130_fd_sc_hd__o21ba_1
X_3539_ _3538_/X _3533_/B _3228_/B vssd1 vssd1 vccd1 vccd1 _3539_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_76_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5209_ _5209_/CLK _5209_/D vssd1 vssd1 vccd1 vccd1 _5209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2910_ _2917_/A _2917_/B _2700_/A vssd1 vssd1 vccd1 vccd1 _2911_/B sky130_fd_sc_hd__o21a_1
XFILLER_31_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3890_ _4985_/Q vssd1 vssd1 vccd1 vccd1 _4882_/B sky130_fd_sc_hd__inv_2
X_2841_ _2841_/A _2843_/B _2841_/C vssd1 vssd1 vccd1 vccd1 _2843_/A sky130_fd_sc_hd__nand3_1
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2772_ _2942_/A _2772_/B vssd1 vssd1 vccd1 vccd1 _2933_/A sky130_fd_sc_hd__nand2_1
X_4511_ _4772_/A vssd1 vssd1 vccd1 vccd1 _4511_/X sky130_fd_sc_hd__buf_2
X_4442_ _4746_/A _5041_/Q vssd1 vssd1 vccd1 vccd1 _4442_/Y sky130_fd_sc_hd__nand2_1
X_4373_ _4373_/A _4373_/B vssd1 vssd1 vccd1 vccd1 _4373_/Y sky130_fd_sc_hd__nand2_1
X_3324_ _3756_/B _5130_/Q vssd1 vssd1 vccd1 vccd1 _3331_/B sky130_fd_sc_hd__nand2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3255_ _3262_/B _3262_/A vssd1 vssd1 vccd1 vccd1 _3255_/X sky130_fd_sc_hd__or2_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3186_ _3186_/A _3186_/B _3186_/C vssd1 vssd1 vccd1 vccd1 _3187_/A sky130_fd_sc_hd__or3_1
XFILLER_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4709_ _4709_/A _4709_/B vssd1 vssd1 vccd1 vccd1 _4710_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3040_ _5235_/Q vssd1 vssd1 vccd1 vccd1 _3730_/B sky130_fd_sc_hd__inv_2
XFILLER_48_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4991_ _5058_/CLK _4991_/D vssd1 vssd1 vccd1 vccd1 _4991_/Q sky130_fd_sc_hd__dfxtp_1
X_3942_ _4962_/Q hold19/A vssd1 vssd1 vccd1 vccd1 _3944_/A sky130_fd_sc_hd__nor2_1
X_3873_ _3879_/A _4902_/A vssd1 vssd1 vccd1 vccd1 _3873_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2824_ _2824_/A _2824_/B vssd1 vssd1 vccd1 vccd1 _2841_/A sky130_fd_sc_hd__nand2_1
X_2755_ _2755_/A _2755_/B vssd1 vssd1 vccd1 vccd1 _2755_/Y sky130_fd_sc_hd__nand2_1
X_2686_ _5268_/Q _4603_/A vssd1 vssd1 vccd1 vccd1 _2925_/B sky130_fd_sc_hd__or2_1
X_4425_ _4479_/A _4547_/B vssd1 vssd1 vccd1 vccd1 _4425_/Y sky130_fd_sc_hd__nand2_1
X_4356_ _4382_/A _4381_/A _4383_/A vssd1 vssd1 vccd1 vccd1 _4378_/D sky130_fd_sc_hd__a21oi_1
XFILLER_86_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3307_/X sky130_fd_sc_hd__clkbuf_2
X_4287_ _5036_/Q vssd1 vssd1 vccd1 vccd1 _4612_/B sky130_fd_sc_hd__inv_2
XFILLER_58_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _3238_/A _3797_/B vssd1 vssd1 vccd1 vccd1 _3238_/Y sky130_fd_sc_hd__nand2_1
X_3169_ _3167_/Y _3168_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5224_/D sky130_fd_sc_hd__a21oi_1
XFILLER_54_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2540_ _5007_/Q vssd1 vssd1 vccd1 vccd1 _4629_/A sky130_fd_sc_hd__inv_2
X_4210_ _4210_/A _4540_/B vssd1 vssd1 vccd1 vccd1 _4211_/B sky130_fd_sc_hd__nand2_1
X_5190_ _5195_/CLK _5190_/D vssd1 vssd1 vccd1 vccd1 _5190_/Q sky130_fd_sc_hd__dfxtp_1
X_4141_ _4141_/A _4141_/B _4141_/C vssd1 vssd1 vccd1 vccd1 _4146_/A sky130_fd_sc_hd__and3_1
X_4072_ _4087_/B _4065_/B _4117_/C _4144_/B vssd1 vssd1 vccd1 vccd1 _4073_/B sky130_fd_sc_hd__o31ai_1
XFILLER_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3023_ _3023_/A _3032_/A vssd1 vssd1 vccd1 vccd1 _3024_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4974_ _5064_/CLK hold20/X vssd1 vssd1 vccd1 vccd1 _4974_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3925_ _4216_/A _4322_/A vssd1 vssd1 vccd1 vccd1 _4096_/B sky130_fd_sc_hd__nor2_1
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3856_ _3844_/X _4943_/X _3845_/X _3855_/Y vssd1 vssd1 vccd1 vccd1 _5096_/D sky130_fd_sc_hd__o211a_1
X_3787_ _3797_/A _3787_/B vssd1 vssd1 vccd1 vccd1 _3787_/Y sky130_fd_sc_hd__nand2_1
X_2807_ _3815_/A vssd1 vssd1 vccd1 vccd1 _4784_/A sky130_fd_sc_hd__clkbuf_2
X_2738_ _2738_/A _2738_/B vssd1 vssd1 vccd1 vccd1 _2739_/A sky130_fd_sc_hd__nor2_1
X_4408_ _4406_/X _4402_/A _4407_/X vssd1 vssd1 vccd1 vccd1 _4408_/X sky130_fd_sc_hd__a21o_1
XFILLER_59_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2669_ _2669_/A _4997_/Q vssd1 vssd1 vccd1 vccd1 _2770_/A sky130_fd_sc_hd__nand2_1
XFILLER_86_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4339_ _4339_/A _4656_/B vssd1 vssd1 vccd1 vccd1 _4340_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3710_ _5147_/Q _3698_/X _3708_/X _3709_/Y vssd1 vssd1 vccd1 vccd1 _5147_/D sky130_fd_sc_hd__o211a_1
X_4690_ _4690_/A _4690_/B vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__nor2_1
X_3641_ _3641_/A _3641_/B vssd1 vssd1 vccd1 vccd1 _3641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3572_ _3573_/A _3574_/A _3573_/B _2898_/X vssd1 vssd1 vccd1 vccd1 _3572_/X sky130_fd_sc_hd__a31o_1
X_2523_ _2534_/A _4547_/A vssd1 vssd1 vccd1 vccd1 _2523_/Y sky130_fd_sc_hd__nand2_1
X_5242_ _5289_/CLK _5242_/D vssd1 vssd1 vccd1 vccd1 _5242_/Q sky130_fd_sc_hd__dfxtp_1
X_5173_ _5209_/CLK _5173_/D vssd1 vssd1 vccd1 vccd1 _5173_/Q sky130_fd_sc_hd__dfxtp_1
X_4124_ _5069_/Q vssd1 vssd1 vccd1 vccd1 _4294_/A sky130_fd_sc_hd__inv_2
Xinput1 enable_in vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_28_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4055_ _4069_/A _4162_/C vssd1 vssd1 vccd1 vccd1 _4163_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3006_ _3688_/B _5155_/Q vssd1 vssd1 vccd1 vccd1 _3143_/B sky130_fd_sc_hd__and2_1
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4957_ _4964_/CLK _4957_/D vssd1 vssd1 vccd1 vccd1 hold22/A sky130_fd_sc_hd__dfxtp_1
X_3908_ _4479_/A _4871_/B vssd1 vssd1 vccd1 vccd1 _3908_/Y sky130_fd_sc_hd__nand2_1
X_4888_ _5088_/Q _4892_/A vssd1 vssd1 vccd1 vccd1 _4888_/Y sky130_fd_sc_hd__nor2_1
X_3839_ _4940_/A _3839_/B vssd1 vssd1 vccd1 vccd1 _3839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5207_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4811_ _4811_/A _4820_/B vssd1 vssd1 vccd1 vccd1 _4811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4742_ _4741_/B _4741_/A _4711_/X vssd1 vssd1 vccd1 vccd1 _4742_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _5021_/Q _5053_/Q vssd1 vssd1 vccd1 vccd1 _4674_/A sky130_fd_sc_hd__nor2_1
X_3624_ _3388_/Y _3635_/A _3406_/Y vssd1 vssd1 vccd1 vccd1 _3631_/A sky130_fd_sc_hd__o21ai_1
X_3555_ _3544_/Y _3472_/Y _3458_/A _2803_/A vssd1 vssd1 vccd1 vccd1 _3555_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3486_ _5222_/Q vssd1 vssd1 vccd1 vccd1 _3767_/B sky130_fd_sc_hd__inv_2
XFILLER_0_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2506_ _2584_/A vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5225_ _5228_/CLK _5225_/D vssd1 vssd1 vccd1 vccd1 _5225_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5156_ _5259_/CLK _5156_/D vssd1 vssd1 vccd1 vccd1 _5156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4107_ _4110_/A _4107_/B vssd1 vssd1 vccd1 vccd1 _4111_/A sky130_fd_sc_hd__nand2_1
X_5087_ _5282_/CLK _5087_/D vssd1 vssd1 vccd1 vccd1 _5087_/Q sky130_fd_sc_hd__dfxtp_1
X_4038_ _5065_/Q vssd1 vssd1 vccd1 vccd1 _4278_/A sky130_fd_sc_hd__inv_2
XFILLER_56_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3340_ _5126_/Q vssd1 vssd1 vccd1 vccd1 _3513_/B sky130_fd_sc_hd__inv_2
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _3271_/A _3271_/B vssd1 vssd1 vccd1 vccd1 _3271_/Y sky130_fd_sc_hd__nand2_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ _5278_/CLK _5010_/D vssd1 vssd1 vccd1 vccd1 _5010_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2986_ _2985_/Y _2986_/B vssd1 vssd1 vccd1 vccd1 _2986_/X sky130_fd_sc_hd__and2b_1
X_4725_ _5014_/Q _4987_/Q _4723_/Y _4724_/X _4713_/X vssd1 vssd1 vccd1 vccd1 _5014_/D
+ sky130_fd_sc_hd__o221a_1
X_4656_ _4656_/A _4656_/B vssd1 vssd1 vccd1 vccd1 _4657_/B sky130_fd_sc_hd__nand2_1
X_3607_ _3607_/A _3607_/B vssd1 vssd1 vccd1 vccd1 _3608_/B sky130_fd_sc_hd__nand2_1
X_4587_ _4994_/Q _5026_/Q _4810_/B _4813_/A _4807_/A vssd1 vssd1 vccd1 vccd1 _4797_/A
+ sky130_fd_sc_hd__o2111ai_2
X_3538_ _3538_/A _3538_/B _3538_/C vssd1 vssd1 vccd1 vccd1 _3538_/X sky130_fd_sc_hd__and3_1
XFILLER_1_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3469_ _5215_/Q vssd1 vssd1 vccd1 vccd1 _3784_/B sky130_fd_sc_hd__inv_2
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5208_ _5209_/CLK _5208_/D vssd1 vssd1 vccd1 vccd1 _5208_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5139_ _5251_/CLK _5139_/D vssd1 vssd1 vccd1 vccd1 _5139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _2834_/Y _2837_/X _2839_/X vssd1 vssd1 vccd1 vccd1 _5252_/D sky130_fd_sc_hd__o21a_1
XFILLER_31_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2771_ _2771_/A _2943_/A vssd1 vssd1 vccd1 vccd1 _2772_/B sky130_fd_sc_hd__nor2_1
X_4510_ _4509_/B _4509_/A _4436_/X vssd1 vssd1 vccd1 vccd1 _4510_/X sky130_fd_sc_hd__a21o_1
XFILLER_11_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4441_ _4745_/A _4441_/B _4434_/A vssd1 vssd1 vccd1 vccd1 _4441_/X sky130_fd_sc_hd__or3b_1
X_4372_ _4987_/Q _4537_/B vssd1 vssd1 vccd1 vccd1 _4372_/Y sky130_fd_sc_hd__nor2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _5226_/Q vssd1 vssd1 vccd1 vccd1 _3756_/B sky130_fd_sc_hd__inv_2
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3254_ _3254_/A _3254_/B vssd1 vssd1 vccd1 vccd1 _3262_/A sky130_fd_sc_hd__and2_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3185_ _5221_/Q _2972_/X _3183_/Y _3184_/X _2980_/X vssd1 vssd1 vccd1 vccd1 _5221_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2969_ _2969_/A _2969_/B vssd1 vssd1 vccd1 vccd1 _2969_/Y sky130_fd_sc_hd__nor2_1
X_4708_ _4708_/A _4696_/X vssd1 vssd1 vccd1 vccd1 _4709_/A sky130_fd_sc_hd__or2b_1
X_4639_ _4639_/A _4639_/B vssd1 vssd1 vccd1 vccd1 _4731_/A sky130_fd_sc_hd__nor2_1
XFILLER_78_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4990_ _5201_/CLK _4990_/D vssd1 vssd1 vccd1 vccd1 _4990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3941_ _4966_/Q hold18/A vssd1 vssd1 vccd1 vccd1 _3945_/B sky130_fd_sc_hd__and2b_1
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3872_ _5091_/Q vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__inv_2
X_2823_ _5254_/Q _2814_/X _2819_/Y _2820_/X _2822_/X vssd1 vssd1 vccd1 vccd1 _5254_/D
+ sky130_fd_sc_hd__o221a_1
X_2754_ _5288_/Q _5021_/Q vssd1 vssd1 vccd1 vccd1 _2755_/B sky130_fd_sc_hd__nand2_1
X_2685_ _2677_/Y _2679_/Y _2773_/A vssd1 vssd1 vccd1 vccd1 _2685_/Y sky130_fd_sc_hd__a21oi_1
X_4424_ _4784_/A vssd1 vssd1 vccd1 vccd1 _4424_/X sky130_fd_sc_hd__clkbuf_4
X_4355_ _5083_/Q _5051_/Q vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__nor2_1
X_3306_ _5198_/Q _3261_/X _3303_/X _3305_/Y vssd1 vssd1 vccd1 vccd1 _5198_/D sky130_fd_sc_hd__o211a_1
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ _5068_/Q _5036_/Q vssd1 vssd1 vccd1 vccd1 _4289_/A sky130_fd_sc_hd__nor2_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _5210_/Q vssd1 vssd1 vccd1 vccd1 _3797_/B sky130_fd_sc_hd__inv_2
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3168_ _3505_/A _5224_/Q vssd1 vssd1 vccd1 vccd1 _3168_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3099_ _3714_/B _5145_/Q vssd1 vssd1 vccd1 vccd1 _3100_/A sky130_fd_sc_hd__nand2_1
XFILLER_81_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4140_ _5063_/Q _5062_/Q _5061_/Q vssd1 vssd1 vccd1 vccd1 _4141_/C sky130_fd_sc_hd__and3_1
X_4071_ _4130_/B _5083_/Q _4058_/X _5084_/Q vssd1 vssd1 vccd1 vccd1 _4073_/A sky130_fd_sc_hd__a31oi_1
X_3022_ _3703_/B _5149_/Q vssd1 vssd1 vccd1 vccd1 _3032_/A sky130_fd_sc_hd__and2_1
XFILLER_55_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4973_ _5064_/CLK _4973_/D vssd1 vssd1 vccd1 vccd1 hold20/A sky130_fd_sc_hd__dfxtp_1
X_3924_ _5075_/Q vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__inv_2
X_3855_ _3861_/A _4931_/A vssd1 vssd1 vccd1 vccd1 _3855_/Y sky130_fd_sc_hd__nand2_1
X_3786_ _3826_/A vssd1 vssd1 vccd1 vccd1 _3797_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2806_ _2806_/A _2806_/B _2806_/C vssd1 vssd1 vccd1 vccd1 _2806_/X sky130_fd_sc_hd__and3_1
X_2737_ _2731_/Y _2722_/A _2733_/B vssd1 vssd1 vccd1 vccd1 _2738_/A sky130_fd_sc_hd__o21ai_1
X_2668_ _5264_/Q vssd1 vssd1 vccd1 vccd1 _2669_/A sky130_fd_sc_hd__inv_2
X_4407_ _4501_/A vssd1 vssd1 vccd1 vccd1 _4407_/X sky130_fd_sc_hd__buf_2
X_2599_ _5260_/Q _2584_/X _2585_/X _2598_/Y vssd1 vssd1 vccd1 vccd1 hold10/A sky130_fd_sc_hd__o211a_1
X_4338_ _4338_/A vssd1 vssd1 vccd1 vccd1 _4340_/A sky130_fd_sc_hd__inv_2
XFILLER_59_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4269_ _4269_/A _4486_/B vssd1 vssd1 vccd1 vccd1 _4490_/B sky130_fd_sc_hd__nand2_1
XFILLER_75_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _3640_/A vssd1 vssd1 vccd1 vccd1 _3641_/B sky130_fd_sc_hd__inv_2
X_3571_ _3571_/A _3571_/B vssd1 vssd1 vccd1 vccd1 _3574_/A sky130_fd_sc_hd__nor2_1
X_2522_ _5012_/Q vssd1 vssd1 vccd1 vccd1 _4547_/A sky130_fd_sc_hd__inv_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5241_ _5289_/CLK _5241_/D vssd1 vssd1 vccd1 vccd1 _5241_/Q sky130_fd_sc_hd__dfxtp_1
X_5172_ _5206_/CLK _5172_/D vssd1 vssd1 vccd1 vccd1 _5172_/Q sky130_fd_sc_hd__dfxtp_1
X_4123_ _4313_/A _4065_/C _4122_/Y vssd1 vssd1 vccd1 vccd1 _5071_/D sky130_fd_sc_hd__a21oi_1
X_4054_ _4169_/D _4179_/A _4169_/B _4168_/A vssd1 vssd1 vccd1 vccd1 _4162_/C sky130_fd_sc_hd__a31oi_4
Xinput2 oversample_in[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
XFILLER_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3005_ _3005_/A vssd1 vssd1 vccd1 vccd1 _3142_/A sky130_fd_sc_hd__inv_2
XFILLER_24_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ _4964_/CLK _4956_/D vssd1 vssd1 vccd1 vccd1 _4956_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3907_/X sky130_fd_sc_hd__clkbuf_4
X_4887_ _4887_/A _4887_/B vssd1 vssd1 vccd1 vccd1 _4892_/A sky130_fd_sc_hd__and2_1
X_3838_ _5099_/Q _3832_/X _3829_/X _3837_/Y vssd1 vssd1 vccd1 vccd1 _5099_/D sky130_fd_sc_hd__o211a_1
X_3769_ _3771_/A _3769_/B vssd1 vssd1 vccd1 vccd1 _3769_/Y sky130_fd_sc_hd__nand2_1
XFILLER_10_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _4810_/A _4810_/B _4810_/C vssd1 vssd1 vccd1 vccd1 _4810_/X sky130_fd_sc_hd__and3_1
XFILLER_61_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4741_ _4741_/A _4741_/B vssd1 vssd1 vccd1 vccd1 _4741_/Y sky130_fd_sc_hd__nor2_1
X_4672_ _4687_/A vssd1 vssd1 vccd1 vccd1 _4681_/C sky130_fd_sc_hd__inv_2
X_3623_ _5170_/Q _3601_/X _3589_/X _3622_/X vssd1 vssd1 vccd1 vccd1 _5170_/D sky130_fd_sc_hd__o211a_1
X_3554_ _3544_/Y _3458_/A _3472_/Y vssd1 vssd1 vccd1 vccd1 _3554_/Y sky130_fd_sc_hd__a21oi_1
X_3485_ _5222_/Q _3513_/B _3515_/A _3515_/B vssd1 vssd1 vccd1 vccd1 _3485_/Y sky130_fd_sc_hd__o22ai_4
X_2505_ _3738_/A vssd1 vssd1 vccd1 vccd1 _2584_/A sky130_fd_sc_hd__buf_2
X_5224_ _5228_/CLK _5224_/D vssd1 vssd1 vccd1 vccd1 _5224_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5155_ _5259_/CLK _5155_/D vssd1 vssd1 vccd1 vccd1 _5155_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5086_ _5086_/CLK _5086_/D vssd1 vssd1 vccd1 vccd1 _5086_/Q sky130_fd_sc_hd__dfxtp_1
X_4106_ _4322_/A _4106_/B vssd1 vssd1 vccd1 vccd1 _4107_/B sky130_fd_sc_hd__nor2_1
X_4037_ _4053_/A vssd1 vssd1 vccd1 vccd1 _4141_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4939_ _4939_/A vssd1 vssd1 vccd1 vccd1 _4939_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_20_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3270_ _5205_/Q _3252_/X _3268_/Y _3269_/X _3259_/X vssd1 vssd1 vccd1 vccd1 _5205_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4724_ _4723_/B _4723_/A _4711_/X vssd1 vssd1 vccd1 vccd1 _4724_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2985_ _4992_/Q _2985_/B vssd1 vssd1 vccd1 vccd1 _2985_/Y sky130_fd_sc_hd__nor2_1
X_4655_ _4655_/A vssd1 vssd1 vccd1 vccd1 _4666_/B sky130_fd_sc_hd__inv_2
X_3606_ _3611_/B _3611_/A vssd1 vssd1 vccd1 vccd1 _3607_/A sky130_fd_sc_hd__or2_1
X_4586_ _4816_/A _4819_/B _4826_/B vssd1 vssd1 vccd1 vccd1 _4807_/A sky130_fd_sc_hd__nand3_1
X_3537_ _3601_/A vssd1 vssd1 vccd1 vccd1 _3537_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_88_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3468_ _3551_/B _3468_/B vssd1 vssd1 vccd1 vccd1 _3473_/B sky130_fd_sc_hd__or2_1
X_3399_ _5101_/Q _3833_/B vssd1 vssd1 vccd1 vccd1 _3400_/A sky130_fd_sc_hd__nor2_1
X_5207_ _5207_/CLK _5207_/D vssd1 vssd1 vccd1 vccd1 _5207_/Q sky130_fd_sc_hd__dfxtp_1
X_5138_ _5251_/CLK _5138_/D vssd1 vssd1 vccd1 vccd1 _5138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5069_ _5070_/CLK _5069_/D vssd1 vssd1 vccd1 vccd1 _5069_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2770_ _2770_/A vssd1 vssd1 vccd1 vccd1 _2943_/A sky130_fd_sc_hd__inv_2
X_4440_ _4440_/A _4440_/B vssd1 vssd1 vccd1 vccd1 _4441_/B sky130_fd_sc_hd__nor2_1
X_4371_ _4369_/Y _4679_/B _4873_/A vssd1 vssd1 vccd1 vccd1 _5054_/D sky130_fd_sc_hd__a21oi_1
X_3322_ _5196_/Q _3307_/X _3320_/X _3321_/Y _3315_/X vssd1 vssd1 vccd1 vccd1 _5196_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _3253_/A _3253_/B vssd1 vssd1 vccd1 vccd1 _3257_/A sky130_fd_sc_hd__nor2_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ _3187_/C _3140_/B _3015_/B _2866_/X vssd1 vssd1 vccd1 vccd1 _3184_/X sky130_fd_sc_hd__a31o_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2968_ _2977_/A _2968_/B vssd1 vssd1 vccd1 vccd1 _2969_/B sky130_fd_sc_hd__or2_1
X_4707_ _4705_/X _4706_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5017_/D sky130_fd_sc_hd__a21oi_1
X_2899_ _2900_/A _2901_/A _2900_/B _2898_/X vssd1 vssd1 vccd1 vccd1 _2899_/X sky130_fd_sc_hd__a31o_1
X_4638_ _4623_/A _4623_/B _4636_/Y _4634_/A _4637_/X vssd1 vssd1 vccd1 vccd1 _4719_/B
+ sky130_fd_sc_hd__o221a_1
X_4569_ _4801_/A _4569_/B vssd1 vssd1 vccd1 vccd1 _4591_/B sky130_fd_sc_hd__nor2_1
XFILLER_76_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3940_ hold18/A _4966_/Q vssd1 vssd1 vccd1 vccd1 _3945_/A sky130_fd_sc_hd__and2b_1
XFILLER_51_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3871_ _3867_/X _4947_/X _3868_/X _3870_/Y vssd1 vssd1 vccd1 vccd1 _5092_/D sky130_fd_sc_hd__o211a_1
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2822_ _3259_/A vssd1 vssd1 vccd1 vccd1 _2822_/X sky130_fd_sc_hd__clkbuf_2
X_2753_ _5288_/Q _5021_/Q vssd1 vssd1 vccd1 vccd1 _2755_/A sky130_fd_sc_hd__or2_1
X_2684_ _2684_/A _2935_/A vssd1 vssd1 vccd1 vccd1 _2773_/A sky130_fd_sc_hd__nand2_1
X_4423_ _4423_/A _4423_/B vssd1 vssd1 vccd1 vccd1 _4423_/X sky130_fd_sc_hd__and2_1
X_4354_ _4344_/A _4340_/A _4349_/Y _4353_/X vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__o211a_1
XFILLER_86_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _3295_/A _3304_/X _4940_/A vssd1 vssd1 vccd1 vccd1 _3305_/Y sky130_fd_sc_hd__o21ai_1
X_4285_ _4285_/A _4285_/B vssd1 vssd1 vccd1 vccd1 _4471_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _3236_/A _3236_/B vssd1 vssd1 vccd1 vccd1 _3236_/Y sky130_fd_sc_hd__xnor2_1
X_3167_ _3167_/A _3167_/B _3504_/C vssd1 vssd1 vccd1 vccd1 _3167_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3098_ _5145_/Q _3714_/B vssd1 vssd1 vccd1 vccd1 _3101_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4070_ _4086_/A vssd1 vssd1 vccd1 vccd1 _4130_/B sky130_fd_sc_hd__clkbuf_2
X_3021_ _5149_/Q _3703_/B vssd1 vssd1 vccd1 vccd1 _3023_/A sky130_fd_sc_hd__nor2_1
X_4972_ _5080_/CLK _4972_/D vssd1 vssd1 vccd1 vccd1 _4972_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3923_ _5076_/Q vssd1 vssd1 vccd1 vccd1 _4216_/A sky130_fd_sc_hd__inv_2
X_3854_ _5096_/Q vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__inv_2
X_2805_ _2806_/A _2806_/B _2806_/C vssd1 vssd1 vccd1 vccd1 _2805_/Y sky130_fd_sc_hd__a21oi_1
X_3785_ _5119_/Q _3779_/X _3776_/X _3784_/Y vssd1 vssd1 vccd1 vccd1 _5119_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2736_ _2857_/A vssd1 vssd1 vccd1 vccd1 _2736_/Y sky130_fd_sc_hd__inv_2
X_2667_ _2667_/A _5263_/Q vssd1 vssd1 vccd1 vccd1 _2767_/A sky130_fd_sc_hd__nand2_1
X_4406_ _4406_/A _4406_/B _4335_/A vssd1 vssd1 vccd1 vccd1 _4406_/X sky130_fd_sc_hd__or3b_1
X_2598_ _3676_/A _4579_/A vssd1 vssd1 vccd1 vccd1 _2598_/Y sky130_fd_sc_hd__nand2_1
X_4337_ _4339_/A _4656_/B vssd1 vssd1 vccd1 vccd1 _4338_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4268_ _5063_/Q _5031_/Q vssd1 vssd1 vccd1 vccd1 _4486_/B sky130_fd_sc_hd__nand2_1
X_3219_ _3218_/X _3203_/Y _2930_/X vssd1 vssd1 vccd1 vccd1 _3219_/X sky130_fd_sc_hd__a21o_1
X_4199_ _5053_/Q vssd1 vssd1 vccd1 vccd1 _4537_/B sky130_fd_sc_hd__inv_2
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _3576_/B _3576_/A vssd1 vssd1 vccd1 vccd1 _3573_/A sky130_fd_sc_hd__or2_1
X_2521_ _5280_/Q _2506_/X _2507_/X hold1/X vssd1 vssd1 vccd1 vccd1 _5280_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _5254_/CLK _5240_/D vssd1 vssd1 vccd1 vccd1 _5240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5171_ _5206_/CLK _5171_/D vssd1 vssd1 vccd1 vccd1 _5171_/Q sky130_fd_sc_hd__dfxtp_1
X_4122_ _4313_/A _4065_/C _4093_/B vssd1 vssd1 vccd1 vccd1 _4122_/Y sky130_fd_sc_hd__o21ai_1
X_4053_ _4053_/A vssd1 vssd1 vccd1 vccd1 _4069_/A sky130_fd_sc_hd__inv_2
XFILLER_56_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 oversample_in[1] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_3004_ _5154_/Q _3690_/B vssd1 vssd1 vccd1 vccd1 _3005_/A sky130_fd_sc_hd__nor2_1
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4955_ _4964_/CLK _4955_/D vssd1 vssd1 vccd1 vccd1 _4956_/D sky130_fd_sc_hd__dfxtp_1
X_3906_ _5093_/Q _3887_/Y _3889_/X _3897_/X _3905_/Y vssd1 vssd1 vccd1 vccd1 _4951_/S
+ sky130_fd_sc_hd__o2111a_4
XFILLER_32_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4886_ _4881_/Y _4882_/Y _4883_/Y _4884_/Y _4885_/X vssd1 vssd1 vccd1 vccd1 _4887_/B
+ sky130_fd_sc_hd__o2111a_1
X_3837_ _3837_/A _3837_/B vssd1 vssd1 vccd1 vccd1 _3837_/Y sky130_fd_sc_hd__nand2_1
X_3768_ _5126_/Q _3766_/X _3763_/X _3767_/Y vssd1 vssd1 vccd1 vccd1 _5126_/D sky130_fd_sc_hd__o211a_1
X_2719_ _2890_/A _2893_/B _2643_/A vssd1 vssd1 vccd1 vccd1 _2719_/X sky130_fd_sc_hd__or3b_1
X_3699_ _3703_/A _3699_/B vssd1 vssd1 vccd1 vccd1 _3699_/Y sky130_fd_sc_hd__nand2_1
XFILLER_74_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4740_ _4637_/A _4637_/B _4739_/Y vssd1 vssd1 vccd1 vccd1 _4741_/B sky130_fd_sc_hd__o21a_1
X_4671_ hold6/A _4671_/B vssd1 vssd1 vccd1 vccd1 _4687_/A sky130_fd_sc_hd__nor2_1
X_3622_ _3616_/X _3621_/Y _3577_/X vssd1 vssd1 vccd1 vccd1 _3622_/X sky130_fd_sc_hd__a21o_1
X_3553_ _5184_/Q _3537_/X _3303_/X _3552_/X vssd1 vssd1 vccd1 vccd1 _5184_/D sky130_fd_sc_hd__o211a_1
X_3484_ _3538_/A _3538_/C _3483_/X vssd1 vssd1 vccd1 vccd1 _3515_/B sky130_fd_sc_hd__a21oi_2
X_2504_ _5284_/Q _2481_/X _2485_/X _2503_/Y vssd1 vssd1 vccd1 vccd1 hold13/A sky130_fd_sc_hd__o211a_1
X_5223_ _5228_/CLK _5223_/D vssd1 vssd1 vccd1 vccd1 _5223_/Q sky130_fd_sc_hd__dfxtp_1
X_5154_ _5259_/CLK _5154_/D vssd1 vssd1 vccd1 vccd1 _5154_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4105_ _4105_/A vssd1 vssd1 vccd1 vccd1 _5077_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_29_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5085_ _5086_/CLK _5085_/D vssd1 vssd1 vccd1 vccd1 _5085_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4036_ _4987_/Q _5060_/Q _5059_/Q vssd1 vssd1 vccd1 vccd1 _4053_/A sky130_fd_sc_hd__and3_1
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4938_ _4975_/Q _4976_/Q vssd1 vssd1 vccd1 vccd1 _4939_/A sky130_fd_sc_hd__and2_1
X_4869_ _4873_/A input2/X vssd1 vssd1 vccd1 vccd1 _4870_/A sky130_fd_sc_hd__or2_1
XFILLER_20_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2984_ _2990_/B _5258_/Q vssd1 vssd1 vccd1 vccd1 _2991_/B sky130_fd_sc_hd__nand2_1
X_4723_ _4723_/A _4723_/B vssd1 vssd1 vccd1 vccd1 _4723_/Y sky130_fd_sc_hd__nor2_1
X_4654_ _4656_/A _4656_/B vssd1 vssd1 vccd1 vccd1 _4655_/A sky130_fd_sc_hd__nor2_1
X_3605_ _3605_/A _3605_/B vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__nor2_1
X_4585_ _4993_/Q _5025_/Q vssd1 vssd1 vccd1 vccd1 _4826_/B sky130_fd_sc_hd__nand2_1
X_3536_ _5187_/Q _3512_/X _3534_/Y _3535_/X _3518_/X vssd1 vssd1 vccd1 vccd1 _5187_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_88_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5206_ _5206_/CLK _5206_/D vssd1 vssd1 vccd1 vccd1 _5206_/Q sky130_fd_sc_hd__dfxtp_1
X_3467_ _3475_/B _3467_/B vssd1 vssd1 vccd1 vccd1 _3468_/B sky130_fd_sc_hd__or2_1
XFILLER_69_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3398_ _5197_/Q vssd1 vssd1 vccd1 vccd1 _3833_/B sky130_fd_sc_hd__inv_2
X_5137_ _5137_/CLK _5137_/D vssd1 vssd1 vccd1 vccd1 _5137_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5068_ _5068_/CLK _5068_/D vssd1 vssd1 vccd1 vccd1 _5068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4019_ _4019_/A _4019_/B vssd1 vssd1 vccd1 vccd1 _4020_/A sky130_fd_sc_hd__nand2_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4711_/A _5054_/Q vssd1 vssd1 vccd1 vccd1 _4679_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3321_ _3310_/A _3317_/X _3319_/Y _3504_/C vssd1 vssd1 vccd1 vccd1 _3321_/Y sky130_fd_sc_hd__o31ai_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3252_/X sky130_fd_sc_hd__clkbuf_2
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3183_ _3187_/C _3015_/B _3140_/B vssd1 vssd1 vccd1 vccd1 _3183_/Y sky130_fd_sc_hd__a21oi_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2967_ _2967_/A _2963_/C vssd1 vssd1 vccd1 vccd1 _2969_/A sky130_fd_sc_hd__or2b_1
X_2898_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2898_/X sky130_fd_sc_hd__clkbuf_4
X_4706_ _4746_/A _5017_/Q vssd1 vssd1 vccd1 vccd1 _4706_/Y sky130_fd_sc_hd__nand2_1
X_4637_ _4637_/A _4637_/B _4637_/C vssd1 vssd1 vccd1 vccd1 _4637_/X sky130_fd_sc_hd__or3_1
XFILLER_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4568_ _4997_/Q _5029_/Q vssd1 vssd1 vccd1 vccd1 _4800_/C sky130_fd_sc_hd__nand2_1
X_4499_ _4387_/X _4496_/Y _4497_/X _4424_/X _4498_/Y vssd1 vssd1 vccd1 vccd1 _5030_/D
+ sky130_fd_sc_hd__o311a_1
X_3519_ _5190_/Q _3512_/X _3516_/Y _3517_/X _3518_/X vssd1 vssd1 vccd1 vccd1 _5190_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_20_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _5063_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_4_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_63_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3870_ _3879_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3870_/Y sky130_fd_sc_hd__nand2_1
X_2821_ _4103_/A vssd1 vssd1 vccd1 vccd1 _3259_/A sky130_fd_sc_hd__clkbuf_4
X_2752_ _2806_/A _2806_/B _2804_/B vssd1 vssd1 vccd1 vccd1 _2752_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4422_ _4423_/B _4423_/A vssd1 vssd1 vccd1 vccd1 _4422_/Y sky130_fd_sc_hd__nor2_1
X_2683_ _2683_/A _2683_/B vssd1 vssd1 vccd1 vccd1 _2935_/A sky130_fd_sc_hd__nor2_1
X_4353_ _4396_/C _4396_/B _4353_/C vssd1 vssd1 vccd1 vccd1 _4353_/X sky130_fd_sc_hd__or3_1
X_4284_ _5067_/Q _5035_/Q vssd1 vssd1 vccd1 vccd1 _4285_/B sky130_fd_sc_hd__nand2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3304_ _3304_/A _3304_/B _3309_/A vssd1 vssd1 vccd1 vccd1 _3304_/X sky130_fd_sc_hd__and3_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _5211_/Q _3190_/X _3233_/Y _3234_/X _3194_/X vssd1 vssd1 vccd1 vccd1 _5211_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3166_ _3170_/A _3166_/B _3166_/C vssd1 vssd1 vccd1 vccd1 _3167_/A sky130_fd_sc_hd__nand3b_1
XFILLER_66_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3097_ _5241_/Q vssd1 vssd1 vccd1 vccd1 _3714_/B sky130_fd_sc_hd__inv_2
XFILLER_62_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3999_ _3994_/Y _4009_/B _3996_/Y vssd1 vssd1 vccd1 vccd1 _4001_/A sky130_fd_sc_hd__a21o_1
XFILLER_10_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5201_/CLK sky130_fd_sc_hd__clkbuf_16
X_3020_ _3032_/B _3020_/B vssd1 vssd1 vccd1 vccd1 _3229_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4971_ _5080_/CLK _4971_/D vssd1 vssd1 vccd1 vccd1 _4972_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3922_ _4110_/B _5078_/Q _5077_/Q vssd1 vssd1 vccd1 vccd1 _3926_/A sky130_fd_sc_hd__and3_1
X_3853_ _3881_/A vssd1 vssd1 vccd1 vccd1 _3861_/A sky130_fd_sc_hd__clkbuf_4
X_2804_ _2804_/A _2804_/B vssd1 vssd1 vccd1 vccd1 _2806_/C sky130_fd_sc_hd__nor2_1
X_3784_ _3784_/A _3784_/B vssd1 vssd1 vccd1 vccd1 _3784_/Y sky130_fd_sc_hd__nand2_1
X_2735_ _2780_/A _2720_/Y _2734_/X vssd1 vssd1 vccd1 vccd1 _2824_/A sky130_fd_sc_hd__o21bai_1
X_2666_ _2963_/A _2963_/C _2963_/B vssd1 vssd1 vccd1 vccd1 _2953_/A sky130_fd_sc_hd__a21oi_4
X_4405_ _4987_/Q _5048_/Q _4403_/Y _4404_/X _4183_/X vssd1 vssd1 vccd1 vccd1 _5048_/D
+ sky130_fd_sc_hd__o221a_1
X_4336_ _5049_/Q vssd1 vssd1 vccd1 vccd1 _4656_/B sky130_fd_sc_hd__inv_2
X_2597_ _4993_/Q vssd1 vssd1 vccd1 vccd1 _4579_/A sky130_fd_sc_hd__clkinv_2
XFILLER_59_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4267_ _4267_/A _4594_/B vssd1 vssd1 vccd1 vccd1 _4269_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4198_ _5085_/Q vssd1 vssd1 vccd1 vccd1 _4362_/B sky130_fd_sc_hd__inv_2
XFILLER_74_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3218_ _3218_/A _3218_/B vssd1 vssd1 vccd1 vccd1 _3218_/X sky130_fd_sc_hd__or2_1
X_3149_ _5254_/Q vssd1 vssd1 vccd1 vccd1 _3679_/B sky130_fd_sc_hd__inv_2
XFILLER_82_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2520_ _2534_/A _4726_/B vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__nand2_1
X_5170_ _5206_/CLK _5170_/D vssd1 vssd1 vccd1 vccd1 _5170_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4121_ _4873_/A _4121_/B _4121_/C vssd1 vssd1 vccd1 vccd1 _5072_/D sky130_fd_sc_hd__nor3_1
XFILLER_68_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4052_ _4077_/B _4052_/B _4117_/C vssd1 vssd1 vccd1 vccd1 _4060_/B sky130_fd_sc_hd__nor3_1
XFILLER_68_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3003_ _5250_/Q vssd1 vssd1 vccd1 vccd1 _3690_/B sky130_fd_sc_hd__inv_2
Xinput4 oversample_in[2] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4954_ _4964_/CLK _4954_/D vssd1 vssd1 vccd1 vccd1 _4954_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3905_ _3861_/B _4984_/Q _3898_/Y _3900_/X _3904_/X vssd1 vssd1 vccd1 vccd1 _3905_/Y
+ sky130_fd_sc_hd__a2111oi_1
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4885_ _4977_/Q _4890_/B _4890_/A _4978_/Q vssd1 vssd1 vccd1 vccd1 _4885_/X sky130_fd_sc_hd__o2bb2a_1
X_3836_ _5100_/Q _3832_/X _3829_/X _3835_/Y vssd1 vssd1 vccd1 vccd1 _5100_/D sky130_fd_sc_hd__o211a_1
X_3767_ _3771_/A _3767_/B vssd1 vssd1 vccd1 vccd1 _3767_/Y sky130_fd_sc_hd__nand2_1
X_2718_ _2889_/B _2718_/B vssd1 vssd1 vccd1 vccd1 _2893_/B sky130_fd_sc_hd__nand2_1
X_3698_ _3725_/A vssd1 vssd1 vccd1 vccd1 _3698_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2649_ _4598_/A _5267_/Q vssd1 vssd1 vccd1 vccd1 _2683_/B sky130_fd_sc_hd__and2_1
XFILLER_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4319_ _4434_/B _4319_/B vssd1 vssd1 vccd1 vccd1 _4319_/X sky130_fd_sc_hd__or2_1
XFILLER_55_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4670_ _5020_/Q _5052_/Q _4690_/B _4687_/D vssd1 vssd1 vccd1 vccd1 _4681_/A sky130_fd_sc_hd__o22ai_1
XFILLER_14_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3621_ _3621_/A _3621_/B vssd1 vssd1 vccd1 vccd1 _3621_/Y sky130_fd_sc_hd__nand2_1
X_3552_ _3548_/B _3551_/Y _3272_/X vssd1 vssd1 vccd1 vccd1 _3552_/X sky130_fd_sc_hd__a21o_1
X_2503_ _2516_/A _4656_/A vssd1 vssd1 vccd1 vccd1 _2503_/Y sky130_fd_sc_hd__nand2_1
X_3483_ _3527_/B _3483_/B _3354_/Y vssd1 vssd1 vccd1 vccd1 _3483_/X sky130_fd_sc_hd__or3b_1
X_5222_ _5228_/CLK _5222_/D vssd1 vssd1 vccd1 vccd1 _5222_/Q sky130_fd_sc_hd__dfxtp_2
X_5153_ _5289_/CLK _5153_/D vssd1 vssd1 vccd1 vccd1 _5153_/Q sky130_fd_sc_hd__dfxtp_1
X_4104_ _4104_/A _4104_/B _4760_/A vssd1 vssd1 vccd1 vccd1 _4105_/A sky130_fd_sc_hd__and3_1
XFILLER_84_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5084_ _5086_/CLK _5084_/D vssd1 vssd1 vccd1 vccd1 _5084_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4035_ _4169_/D _4179_/A _4169_/B _4168_/A vssd1 vssd1 vccd1 vccd1 _4141_/A sky130_fd_sc_hd__a31o_2
XFILLER_37_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4937_ _4937_/A vssd1 vssd1 vccd1 vccd1 _4937_/X sky130_fd_sc_hd__clkbuf_1
X_4868_ _4868_/A vssd1 vssd1 vccd1 vccd1 _4978_/D sky130_fd_sc_hd__clkbuf_1
X_3819_ _3832_/A vssd1 vssd1 vccd1 vccd1 _3819_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4799_ _4800_/A _4800_/C _4800_/B vssd1 vssd1 vccd1 vccd1 _4799_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_87_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2983_ _3754_/B _3228_/B vssd1 vssd1 vccd1 vccd1 _2983_/Y sky130_fd_sc_hd__nor2_1
X_4722_ _4728_/A _4722_/B vssd1 vssd1 vccd1 vccd1 _4723_/B sky130_fd_sc_hd__nand2_1
X_4653_ _4708_/A _4710_/A vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__nor2_1
X_3604_ _5174_/Q _3601_/X _3589_/X _3603_/X vssd1 vssd1 vccd1 vccd1 _5174_/D sky130_fd_sc_hd__o211a_1
X_4584_ _4994_/Q _5026_/Q vssd1 vssd1 vccd1 vccd1 _4819_/B sky130_fd_sc_hd__nand2_1
X_3535_ _3534_/B _3534_/A _3312_/X vssd1 vssd1 vccd1 vccd1 _3535_/X sky130_fd_sc_hd__a21o_1
X_3466_ _3780_/B _5121_/Q vssd1 vssd1 vccd1 vccd1 _3467_/B sky130_fd_sc_hd__and2_1
X_5205_ _5206_/CLK _5205_/D vssd1 vssd1 vccd1 vccd1 _5205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3397_ _5197_/Q _3389_/Y _3655_/A _3650_/B vssd1 vssd1 vccd1 vccd1 _3645_/A sky130_fd_sc_hd__o22ai_2
XFILLER_69_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5136_ _5201_/CLK _5136_/D vssd1 vssd1 vccd1 vccd1 _5136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5067_ _5068_/CLK _5067_/D vssd1 vssd1 vccd1 vccd1 _5067_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4018_ _4018_/A vssd1 vssd1 vccd1 vccd1 _4021_/A sky130_fd_sc_hd__inv_2
XFILLER_37_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3320_ _3310_/A _3317_/X _3319_/Y vssd1 vssd1 vccd1 vccd1 _3320_/X sky130_fd_sc_hd__o21a_1
XFILLER_3_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3634_/A sky130_fd_sc_hd__clkbuf_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3182_ _3186_/B _3186_/C _3186_/A vssd1 vssd1 vccd1 vccd1 _3187_/C sky130_fd_sc_hd__o21ai_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2966_ _4994_/Q _2966_/B vssd1 vssd1 vccd1 vccd1 _2967_/A sky130_fd_sc_hd__nor2_1
X_2897_ _2904_/B _2904_/A vssd1 vssd1 vccd1 vccd1 _2900_/A sky130_fd_sc_hd__nand2_1
X_4705_ _4745_/A _4705_/B _4705_/C vssd1 vssd1 vccd1 vccd1 _4705_/X sky130_fd_sc_hd__or3_1
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4636_ _4748_/B _4630_/A _4748_/A vssd1 vssd1 vccd1 vccd1 _4636_/Y sky130_fd_sc_hd__o21bai_1
X_4567_ _4998_/Q _5030_/Q vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4498_ _4754_/B _4569_/B vssd1 vssd1 vccd1 vccd1 _4498_/Y sky130_fd_sc_hd__nand2_1
X_3518_ _4183_/A vssd1 vssd1 vccd1 vccd1 _3518_/X sky130_fd_sc_hd__clkbuf_2
X_3449_ _3449_/A vssd1 vssd1 vccd1 vccd1 _3573_/B sky130_fd_sc_hd__inv_2
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _5219_/CLK _5119_/D vssd1 vssd1 vccd1 vccd1 _5119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2820_ _2819_/B _2819_/A _2603_/A vssd1 vssd1 vccd1 vccd1 _2820_/X sky130_fd_sc_hd__a21o_1
X_2751_ _5020_/Q _2751_/B vssd1 vssd1 vccd1 vccd1 _2804_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2682_ _2938_/A vssd1 vssd1 vccd1 vccd1 _2684_/A sky130_fd_sc_hd__inv_2
XFILLER_69_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4421_ _4421_/A _4421_/B vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__nor2_1
X_4352_ _4352_/A _4352_/B vssd1 vssd1 vccd1 vccd1 _4396_/C sky130_fd_sc_hd__nand2_1
X_4283_ _4283_/A _4607_/B vssd1 vssd1 vccd1 vccd1 _4285_/A sky130_fd_sc_hd__nand2_1
X_3303_ _3644_/A vssd1 vssd1 vccd1 vccd1 _3303_/X sky130_fd_sc_hd__buf_2
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _3233_/B _3233_/A _2912_/X vssd1 vssd1 vccd1 vccd1 _3234_/X sky130_fd_sc_hd__a21o_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3165_ _3165_/A _3165_/B vssd1 vssd1 vccd1 vccd1 _3166_/C sky130_fd_sc_hd__nor2_1
X_3096_ _5240_/Q _5144_/Q vssd1 vssd1 vccd1 vccd1 _3248_/B sky130_fd_sc_hd__xor2_1
XFILLER_54_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3998_ _4000_/A _3968_/Y _3997_/Y _4000_/B vssd1 vssd1 vccd1 vccd1 _4005_/A sky130_fd_sc_hd__o211ai_2
X_2949_ _2948_/Y _2768_/A _2943_/B vssd1 vssd1 vccd1 vccd1 _2949_/Y sky130_fd_sc_hd__a21oi_2
X_4619_ _4619_/A _4619_/B vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4970_ _5064_/CLK hold5/X vssd1 vssd1 vccd1 vccd1 _4970_/Q sky130_fd_sc_hd__dfxtp_1
X_3921_ _4106_/B vssd1 vssd1 vccd1 vccd1 _4110_/B sky130_fd_sc_hd__inv_2
XFILLER_63_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3852_ _4711_/A vssd1 vssd1 vccd1 vccd1 _3881_/A sky130_fd_sc_hd__buf_4
X_2803_ _2803_/A vssd1 vssd1 vccd1 vccd1 _2803_/X sky130_fd_sc_hd__buf_2
X_3783_ _5120_/Q _3779_/X _3776_/X _3782_/Y vssd1 vssd1 vccd1 vccd1 _5120_/D sky130_fd_sc_hd__o211a_1
X_2734_ _2869_/C _2738_/B _2733_/X vssd1 vssd1 vccd1 vccd1 _2734_/X sky130_fd_sc_hd__or3b_1
X_2665_ _2957_/B _2665_/B vssd1 vssd1 vccd1 vccd1 _2963_/B sky130_fd_sc_hd__nand2_1
X_4404_ _4403_/B _4403_/A _3886_/A vssd1 vssd1 vccd1 vccd1 _4404_/X sky130_fd_sc_hd__a21o_1
X_2596_ _3705_/A vssd1 vssd1 vccd1 vccd1 _3676_/A sky130_fd_sc_hd__clkbuf_2
X_4335_ _4335_/A _4403_/A vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__nor2_1
XFILLER_5_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4266_ _5031_/Q vssd1 vssd1 vccd1 vccd1 _4594_/B sky130_fd_sc_hd__inv_2
X_4197_ _4197_/A vssd1 vssd1 vccd1 vccd1 _5055_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_67_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3217_ _5215_/Q _3190_/X _3215_/Y _3216_/X _3194_/X vssd1 vssd1 vccd1 vccd1 _5215_/D
+ sky130_fd_sc_hd__o221a_1
X_3148_ _5254_/Q _3174_/B _3016_/X _3147_/Y vssd1 vssd1 vccd1 vccd1 _3148_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3079_ _5236_/Q vssd1 vssd1 vccd1 vccd1 _3728_/B sky130_fd_sc_hd__inv_2
XFILLER_54_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4120_ _5071_/Q _4074_/X _4075_/X _4057_/X _5072_/Q vssd1 vssd1 vccd1 vccd1 _4121_/B
+ sky130_fd_sc_hd__a41oi_1
X_4051_ _4064_/A vssd1 vssd1 vccd1 vccd1 _4117_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_83_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3002_ _3143_/A vssd1 vssd1 vccd1 vccd1 _3002_/Y sky130_fd_sc_hd__inv_2
XFILLER_49_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput5 oversample_in[3] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_4953_ _4964_/CLK _4953_/D vssd1 vssd1 vccd1 vccd1 _4954_/D sky130_fd_sc_hd__dfxtp_1
X_3904_ _5096_/Q _3901_/Y _5091_/Q _3902_/Y _3903_/X vssd1 vssd1 vccd1 vccd1 _3904_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4884_ _5090_/Q _4979_/Q vssd1 vssd1 vccd1 vccd1 _4884_/Y sky130_fd_sc_hd__xnor2_1
X_3835_ _3837_/A _3835_/B vssd1 vssd1 vccd1 vccd1 _3835_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3766_ _3792_/A vssd1 vssd1 vccd1 vccd1 _3766_/X sky130_fd_sc_hd__clkbuf_2
X_2717_ _4754_/A _5274_/Q vssd1 vssd1 vccd1 vccd1 _2718_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3697_ _5152_/Q _3685_/X _3695_/X _3696_/Y vssd1 vssd1 vccd1 vccd1 _5152_/D sky130_fd_sc_hd__o211a_1
X_2648_ _2697_/B _2698_/A _5003_/Q _2647_/Y vssd1 vssd1 vccd1 vccd1 _2777_/A sky130_fd_sc_hd__a31o_1
X_2579_ _2594_/A _4801_/A vssd1 vssd1 vccd1 vccd1 _2579_/Y sky130_fd_sc_hd__nand2_1
X_4318_ _4445_/B _4312_/A _4445_/A vssd1 vssd1 vccd1 vccd1 _4318_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4249_ _4249_/A _4258_/A vssd1 vssd1 vccd1 vccd1 _4507_/C sky130_fd_sc_hd__and2_1
XFILLER_74_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3620_ _5171_/Q _3580_/X _3618_/Y _3619_/X _3587_/X vssd1 vssd1 vccd1 vccd1 _5171_/D
+ sky130_fd_sc_hd__o221a_1
X_3551_ _3551_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3551_/Y sky130_fd_sc_hd__nand2_1
X_2502_ _5017_/Q vssd1 vssd1 vccd1 vccd1 _4656_/A sky130_fd_sc_hd__inv_2
X_3482_ _3531_/B _3531_/A _3538_/B vssd1 vssd1 vccd1 vccd1 _3483_/B sky130_fd_sc_hd__or3_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5221_ _5227_/CLK _5221_/D vssd1 vssd1 vccd1 vccd1 _5221_/Q sky130_fd_sc_hd__dfxtp_1
X_5152_ _5289_/CLK _5152_/D vssd1 vssd1 vccd1 vccd1 _5152_/Q sky130_fd_sc_hd__dfxtp_1
X_4103_ _4103_/A vssd1 vssd1 vccd1 vccd1 _4760_/A sky130_fd_sc_hd__buf_4
X_5083_ _5086_/CLK _5083_/D vssd1 vssd1 vccd1 vccd1 _5083_/Q sky130_fd_sc_hd__dfxtp_1
X_4034_ _4033_/A _4033_/C _4506_/A vssd1 vssd1 vccd1 vccd1 _4168_/A sky130_fd_sc_hd__a21oi_2
XFILLER_71_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _4936_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4937_/A sky130_fd_sc_hd__and2_1
XFILLER_52_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4867_ _4873_/A input3/X vssd1 vssd1 vccd1 vccd1 _4868_/A sky130_fd_sc_hd__or2_1
X_3818_ _5107_/Q _3805_/X _3816_/X _3817_/Y vssd1 vssd1 vccd1 vccd1 _5107_/D sky130_fd_sc_hd__o211a_1
X_4798_ _4803_/B _4803_/A vssd1 vssd1 vccd1 vccd1 _4800_/A sky130_fd_sc_hd__or2_1
X_3749_ _3815_/A vssd1 vssd1 vccd1 vccd1 _3802_/A sky130_fd_sc_hd__buf_2
XFILLER_79_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2982_ _5227_/Q vssd1 vssd1 vccd1 vccd1 _3754_/B sky130_fd_sc_hd__inv_2
XFILLER_34_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4721_ _4727_/B _4727_/A vssd1 vssd1 vccd1 vccd1 _4728_/A sky130_fd_sc_hd__or2_1
X_4652_ _4652_/A vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__inv_2
X_3603_ _3595_/X _3602_/Y _3577_/X vssd1 vssd1 vccd1 vccd1 _3603_/X sky130_fd_sc_hd__a21o_1
X_4583_ _4823_/A _4826_/C _4825_/B vssd1 vssd1 vccd1 vccd1 _4816_/A sky130_fd_sc_hd__nand3b_1
X_3534_ _3534_/A _3534_/B vssd1 vssd1 vccd1 vccd1 _3534_/Y sky130_fd_sc_hd__nor2_1
X_3465_ _5121_/Q _3780_/B vssd1 vssd1 vccd1 vccd1 _3475_/B sky130_fd_sc_hd__nor2_1
XFILLER_69_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5204_ _5206_/CLK _5204_/D vssd1 vssd1 vccd1 vccd1 _5204_/Q sky130_fd_sc_hd__dfxtp_1
X_3396_ _3835_/B _5100_/Q _3657_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3650_/B sky130_fd_sc_hd__a22oi_2
XFILLER_84_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5135_ _5203_/CLK _5135_/D vssd1 vssd1 vccd1 vccd1 _5135_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5066_ _5068_/CLK _5066_/D vssd1 vssd1 vccd1 vccd1 _5066_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4017_ _4033_/A _5057_/Q _4017_/C vssd1 vssd1 vccd1 vccd1 _4179_/B sky130_fd_sc_hd__nand3_1
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4919_ _4921_/C _4925_/A vssd1 vssd1 vccd1 vccd1 _4920_/A sky130_fd_sc_hd__and2_1
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _5208_/Q _2928_/X _3247_/X _3249_/X vssd1 vssd1 vccd1 vccd1 _5208_/D sky130_fd_sc_hd__o211a_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3181_ _3181_/A _3191_/B vssd1 vssd1 vccd1 vccd1 _3186_/C sky130_fd_sc_hd__nor2_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4704_ _4704_/A _4704_/B vssd1 vssd1 vccd1 vccd1 _4705_/C sky130_fd_sc_hd__and2_1
X_2965_ _5230_/Q _2928_/X _2962_/X _2964_/Y vssd1 vssd1 vccd1 vccd1 _5230_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2896_ _2896_/A _2896_/B vssd1 vssd1 vccd1 vccd1 _2904_/B sky130_fd_sc_hd__nand2_1
X_4635_ _4737_/A _4737_/B _4634_/X vssd1 vssd1 vccd1 vccd1 _4719_/A sky130_fd_sc_hd__o21bai_1
X_4566_ _4566_/A vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__inv_2
X_3517_ _3516_/B _3516_/A _3312_/X vssd1 vssd1 vccd1 vccd1 _3517_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4497_ _4497_/A _4497_/B _4497_/C vssd1 vssd1 vccd1 vccd1 _4497_/X sky130_fd_sc_hd__and3_1
X_3448_ _3583_/B _3585_/B _3583_/A vssd1 vssd1 vccd1 vccd1 _3541_/B sky130_fd_sc_hd__o21ba_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _5202_/Q vssd1 vssd1 vccd1 vccd1 _3820_/B sky130_fd_sc_hd__inv_2
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5118_ _5219_/CLK _5118_/D vssd1 vssd1 vccd1 vccd1 _5118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5049_ _5051_/CLK _5049_/D vssd1 vssd1 vccd1 vccd1 _5049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2750_ _5287_/Q vssd1 vssd1 vccd1 vccd1 _2751_/B sky130_fd_sc_hd__inv_2
X_2681_ _2681_/A _2681_/B vssd1 vssd1 vccd1 vccd1 _2938_/A sky130_fd_sc_hd__nand2_2
X_4420_ _4873_/A _4420_/B vssd1 vssd1 vccd1 vccd1 _5045_/D sky130_fd_sc_hd__nor2_1
X_4351_ _4351_/A vssd1 vssd1 vccd1 vccd1 _4352_/B sky130_fd_sc_hd__inv_2
X_4282_ _5035_/Q vssd1 vssd1 vccd1 vccd1 _4607_/B sky130_fd_sc_hd__inv_2
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3302_ _5199_/Q _3252_/X _3298_/X _3301_/Y _3259_/X vssd1 vssd1 vccd1 vccd1 _5199_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _3233_/A _3233_/B vssd1 vssd1 vccd1 vccd1 _3233_/Y sky130_fd_sc_hd__nor2_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _3148_/Y _3151_/Y _3170_/B vssd1 vssd1 vccd1 vccd1 _3166_/B sky130_fd_sc_hd__a21o_1
X_3095_ _3254_/A _3254_/B _3094_/X vssd1 vssd1 vccd1 vccd1 _3240_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3997_ _3994_/Y _4009_/B _3996_/Y vssd1 vssd1 vccd1 vccd1 _3997_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_22_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2948_ _2656_/Y _2953_/A _2767_/A vssd1 vssd1 vccd1 vccd1 _2948_/Y sky130_fd_sc_hd__o21ai_1
X_2879_ _2884_/A _2880_/C _2880_/B vssd1 vssd1 vccd1 vccd1 _2879_/Y sky130_fd_sc_hd__a21oi_1
X_4618_ _5005_/Q _5037_/Q vssd1 vssd1 vccd1 vccd1 _4619_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4549_ _5012_/Q _5044_/Q vssd1 vssd1 vccd1 vccd1 _4639_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _4304_/A _4299_/A _4309_/A _4313_/A vssd1 vssd1 vccd1 vccd1 _4106_/B sky130_fd_sc_hd__or4_2
XFILLER_44_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3851_ _4841_/A vssd1 vssd1 vccd1 vccd1 _4711_/A sky130_fd_sc_hd__buf_4
XFILLER_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3782_ _3784_/A _3782_/B vssd1 vssd1 vccd1 vccd1 _3782_/Y sky130_fd_sc_hd__nand2_1
X_2802_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2803_/A sky130_fd_sc_hd__buf_4
X_2733_ _2731_/Y _2733_/B vssd1 vssd1 vccd1 vccd1 _2733_/X sky130_fd_sc_hd__and2b_1
X_2664_ _4574_/A _5262_/Q vssd1 vssd1 vccd1 vccd1 _2665_/B sky130_fd_sc_hd__nand2_1
X_4403_ _4403_/A _4403_/B vssd1 vssd1 vccd1 vccd1 _4403_/Y sky130_fd_sc_hd__nor2_1
X_2595_ _5261_/Q _2584_/X _2585_/X _2594_/Y vssd1 vssd1 vccd1 vccd1 _5261_/D sky130_fd_sc_hd__o211a_1
X_4334_ _4334_/A vssd1 vssd1 vccd1 vccd1 _4403_/A sky130_fd_sc_hd__inv_2
X_4265_ _4494_/A _4494_/B _4264_/Y vssd1 vssd1 vccd1 vccd1 _4484_/B sky130_fd_sc_hd__a21oi_1
X_4196_ _4196_/A _4760_/A _4196_/C vssd1 vssd1 vccd1 vccd1 _4197_/A sky130_fd_sc_hd__and3_1
X_3216_ _3203_/Y _3119_/A _3122_/A _2866_/X vssd1 vssd1 vccd1 vccd1 _3216_/X sky130_fd_sc_hd__a31o_1
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3147_ _3196_/A _3196_/C _3146_/X vssd1 vssd1 vccd1 vccd1 _3147_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3078_ _3276_/A _3276_/B _3077_/X vssd1 vssd1 vccd1 vccd1 _3265_/B sky130_fd_sc_hd__a21oi_1
XFILLER_35_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4141_/A _4141_/B _4068_/A vssd1 vssd1 vccd1 vccd1 _4064_/A sky130_fd_sc_hd__nand3_2
XFILLER_49_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3001_ _5155_/Q _3688_/B vssd1 vssd1 vccd1 vccd1 _3143_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput6 oversample_in[4] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4952_ _4873_/B _4976_/Q _4952_/S vssd1 vssd1 vccd1 vccd1 _4952_/X sky130_fd_sc_hd__mux2_1
X_4883_ _5093_/Q _4982_/Q vssd1 vssd1 vccd1 vccd1 _4883_/Y sky130_fd_sc_hd__xnor2_1
X_3903_ _4902_/A _4981_/Q _5093_/Q _3887_/Y vssd1 vssd1 vccd1 vccd1 _3903_/X sky130_fd_sc_hd__a22o_1
X_3834_ _5101_/Q _3832_/X _3829_/X _3833_/Y vssd1 vssd1 vccd1 vccd1 _5101_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3765_ _5127_/Q _3753_/X _3763_/X _3764_/Y vssd1 vssd1 vccd1 vccd1 _5127_/D sky130_fd_sc_hd__o211a_1
X_3696_ _3703_/A _3696_/B vssd1 vssd1 vccd1 vccd1 _3696_/Y sky130_fd_sc_hd__nand2_1
X_2716_ _2716_/A _2716_/B vssd1 vssd1 vccd1 vccd1 _2890_/A sky130_fd_sc_hd__or2_1
XFILLER_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2647_ _5271_/Q _4612_/A vssd1 vssd1 vccd1 vccd1 _2647_/Y sky130_fd_sc_hd__nor2_1
X_2578_ _4998_/Q vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__inv_2
X_4317_ _4431_/A _4431_/B _4316_/Y vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__o21ai_2
X_4248_ _5059_/Q _5027_/Q vssd1 vssd1 vccd1 vccd1 _4258_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4179_ _4179_/A _4179_/B vssd1 vssd1 vccd1 vccd1 _4179_/Y sky130_fd_sc_hd__nand2_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3550_ _3547_/X _2496_/A _3548_/Y _3549_/Y vssd1 vssd1 vccd1 vccd1 _5185_/D sky130_fd_sc_hd__a31oi_1
X_2501_ _5285_/Q _2481_/X _2485_/X _2500_/Y vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__o211a_1
X_3481_ _3481_/A _3481_/B vssd1 vssd1 vccd1 vccd1 _3538_/B sky130_fd_sc_hd__nand2_1
X_5220_ _5228_/CLK _5220_/D vssd1 vssd1 vccd1 vccd1 _5220_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5151_ _5289_/CLK _5151_/D vssd1 vssd1 vccd1 vccd1 _5151_/Q sky130_fd_sc_hd__dfxtp_1
X_5082_ _5086_/CLK _5082_/D vssd1 vssd1 vccd1 vccd1 _5082_/Q sky130_fd_sc_hd__dfxtp_1
X_4102_ _4097_/A _4064_/A _4210_/A vssd1 vssd1 vccd1 vccd1 _4104_/A sky130_fd_sc_hd__o21ai_1
X_4033_ _4033_/A _4506_/A _4033_/C vssd1 vssd1 vccd1 vccd1 _4169_/B sky130_fd_sc_hd__nand3_2
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _5097_/Q _4935_/B vssd1 vssd1 vccd1 vccd1 _4936_/A sky130_fd_sc_hd__xor2_1
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4866_ _4866_/A vssd1 vssd1 vccd1 vccd1 _4979_/D sky130_fd_sc_hd__clkbuf_1
X_3817_ _3824_/A _3817_/B vssd1 vssd1 vccd1 vccd1 _3817_/Y sky130_fd_sc_hd__nand2_1
X_4797_ _4797_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4803_/A sky130_fd_sc_hd__and2_1
X_3748_ _5133_/Q _3739_/X _3735_/X _3747_/Y vssd1 vssd1 vccd1 vccd1 _5133_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3679_ _3690_/A _3679_/B vssd1 vssd1 vccd1 vccd1 _3679_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2981_ _5228_/Q _2972_/X _2976_/X _2979_/Y _2980_/X vssd1 vssd1 vccd1 vccd1 _5228_/D
+ sky130_fd_sc_hd__o221a_1
Xclkbuf_leaf_41_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5206_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4720_ _4643_/B _4734_/B _4550_/X vssd1 vssd1 vccd1 vccd1 _4727_/A sky130_fd_sc_hd__o21ba_1
X_4651_ _4651_/A _4651_/B vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__nor2_1
Xinput20 phase_in[7] vssd1 vssd1 vccd1 vccd1 _4959_/D sky130_fd_sc_hd__clkbuf_1
X_3602_ _3602_/A _3602_/B vssd1 vssd1 vccd1 vccd1 _3602_/Y sky130_fd_sc_hd__nand2_1
X_4582_ _4829_/B _4828_/A vssd1 vssd1 vccd1 vccd1 _4825_/B sky130_fd_sc_hd__nand2_1
X_3533_ _3533_/A _3533_/B vssd1 vssd1 vccd1 vccd1 _3534_/B sky130_fd_sc_hd__nor2_1
X_3464_ _5217_/Q vssd1 vssd1 vccd1 vccd1 _3780_/B sky130_fd_sc_hd__inv_2
X_5203_ _5203_/CLK _5203_/D vssd1 vssd1 vccd1 vccd1 _5203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3395_ _5099_/Q _5195_/Q vssd1 vssd1 vccd1 vccd1 _3663_/B sky130_fd_sc_hd__or2b_1
X_5134_ _5207_/CLK _5134_/D vssd1 vssd1 vccd1 vccd1 _5134_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5065_ _5068_/CLK _5065_/D vssd1 vssd1 vccd1 vccd1 _5065_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4016_ _4016_/A _4022_/A _4016_/C vssd1 vssd1 vccd1 vccd1 _4017_/C sky130_fd_sc_hd__nand3_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5219_/CLK sky130_fd_sc_hd__clkbuf_16
X_4918_ _4918_/A _5094_/Q vssd1 vssd1 vccd1 vccd1 _4925_/A sky130_fd_sc_hd__nand2_1
XFILLER_32_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4849_ _4849_/A input1/X vssd1 vssd1 vccd1 vccd1 _4850_/A sky130_fd_sc_hd__and2_1
XFILLER_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_23_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _4996_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _3196_/A _3196_/C vssd1 vssd1 vccd1 vccd1 _3191_/B sky130_fd_sc_hd__and2_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2964_ _2953_/A _2963_/X _4940_/A vssd1 vssd1 vccd1 vccd1 _2964_/Y sky130_fd_sc_hd__o21ai_2
Xclkbuf_leaf_14_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5086_/CLK sky130_fd_sc_hd__clkbuf_16
X_4703_ _4516_/X _4698_/X _4700_/X _4424_/X _4702_/Y vssd1 vssd1 vccd1 vccd1 _5018_/D
+ sky130_fd_sc_hd__o311a_1
X_2895_ _5242_/Q _2847_/X _2609_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _5242_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4634_ _4634_/A _4634_/B vssd1 vssd1 vccd1 vccd1 _4634_/X sky130_fd_sc_hd__or2_1
X_4565_ _4779_/A _4781_/C _4564_/Y vssd1 vssd1 vccd1 vccd1 _4566_/A sky130_fd_sc_hd__o21a_1
X_3516_ _3516_/A _3516_/B vssd1 vssd1 vccd1 vccd1 _3516_/Y sky130_fd_sc_hd__nor2_1
X_4496_ _4497_/A _4497_/C _4497_/B vssd1 vssd1 vccd1 vccd1 _4496_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_89_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3447_ _3581_/A _3581_/B _3446_/X vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__o21bai_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3378_ _3436_/A _3434_/A _3593_/A vssd1 vssd1 vccd1 vccd1 _3581_/A sky130_fd_sc_hd__a21o_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_84_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5117_ _5181_/CLK _5117_/D vssd1 vssd1 vccd1 vccd1 _5117_/Q sky130_fd_sc_hd__dfxtp_1
X_5048_ _5283_/CLK _5048_/D vssd1 vssd1 vccd1 vccd1 _5048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2680_ _4794_/A _5266_/Q vssd1 vssd1 vccd1 vccd1 _2681_/B sky130_fd_sc_hd__nand2_1
X_4350_ _4332_/A _4650_/B _4402_/B vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__o21ai_1
X_3301_ _3301_/A _3301_/B vssd1 vssd1 vccd1 vccd1 _3301_/Y sky130_fd_sc_hd__nor2_1
X_4281_ _4474_/A _4474_/B _4280_/X vssd1 vssd1 vccd1 vccd1 _4463_/B sky130_fd_sc_hd__a21oi_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _3110_/B _3236_/B _3110_/A vssd1 vssd1 vccd1 vccd1 _3233_/B sky130_fd_sc_hd__o21ba_1
Xclkbuf_leaf_3_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5282_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3163_ _5255_/Q _3163_/B vssd1 vssd1 vccd1 vccd1 _3170_/B sky130_fd_sc_hd__nor2_1
XFILLER_66_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3094_ _3253_/A _3253_/B _3262_/B vssd1 vssd1 vccd1 vccd1 _3094_/X sky130_fd_sc_hd__or3_1
XFILLER_35_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3996_ _3996_/A vssd1 vssd1 vccd1 vccd1 _3996_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2947_ _5233_/Q _2907_/X _2945_/Y _2946_/X _2914_/X vssd1 vssd1 vccd1 vccd1 _5233_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2878_ _2875_/X _2876_/Y _2877_/Y vssd1 vssd1 vccd1 vccd1 _2884_/A sky130_fd_sc_hd__a21o_1
X_4617_ _4617_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4759_/B sky130_fd_sc_hd__nor2_1
X_4548_ _4735_/A _4548_/B vssd1 vssd1 vccd1 vccd1 _4641_/B sky130_fd_sc_hd__nor2_1
X_4479_ _4479_/A _4563_/B vssd1 vssd1 vccd1 vccd1 _4479_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3850_ _4942_/X _3844_/X _3845_/X _3849_/Y vssd1 vssd1 vccd1 vccd1 _5097_/D sky130_fd_sc_hd__o211a_1
X_3781_ _5121_/Q _3779_/X _3776_/X _3780_/Y vssd1 vssd1 vccd1 vccd1 _5121_/D sky130_fd_sc_hd__o211a_1
X_2801_ _2798_/Y _2800_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5256_/D sky130_fd_sc_hd__a21oi_1
XFILLER_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2732_ _4547_/A _5279_/Q vssd1 vssd1 vccd1 vccd1 _2733_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2663_ _2966_/B _4994_/Q vssd1 vssd1 vccd1 vccd1 _2963_/C sky130_fd_sc_hd__nand2_1
X_4402_ _4402_/A _4402_/B vssd1 vssd1 vccd1 vccd1 _4403_/B sky130_fd_sc_hd__nand2_1
X_2594_ _2594_/A hold7/X vssd1 vssd1 vccd1 vccd1 _2594_/Y sky130_fd_sc_hd__nand2_1
X_4333_ _4351_/A _4333_/B vssd1 vssd1 vccd1 vccd1 _4334_/A sky130_fd_sc_hd__nor2_1
XFILLER_5_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4264_ _4493_/A _4497_/B vssd1 vssd1 vccd1 vccd1 _4264_/Y sky130_fd_sc_hd__nand2_1
X_3215_ _3203_/Y _3122_/A _3119_/A vssd1 vssd1 vccd1 vccd1 _3215_/Y sky130_fd_sc_hd__a21oi_1
X_4195_ _4195_/A _5055_/Q vssd1 vssd1 vccd1 vccd1 _4196_/C sky130_fd_sc_hd__nand2_1
XFILLER_67_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3146_ _3146_/A _3181_/A vssd1 vssd1 vccd1 vccd1 _3146_/X sky130_fd_sc_hd__or2_1
XFILLER_82_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3077_ _3282_/B _3275_/A vssd1 vssd1 vccd1 vccd1 _3077_/X sky130_fd_sc_hd__or2_1
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3979_ _4001_/C _3979_/B vssd1 vssd1 vccd1 vccd1 _3979_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 oversample_in[5] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
X_3000_ _5251_/Q vssd1 vssd1 vccd1 vccd1 _3688_/B sky130_fd_sc_hd__inv_2
XFILLER_49_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4951_ _4888_/Y _4890_/B _4951_/S vssd1 vssd1 vccd1 vccd1 _4951_/X sky130_fd_sc_hd__mux2_1
XFILLER_17_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3902_ _4981_/Q vssd1 vssd1 vccd1 vccd1 _3902_/Y sky130_fd_sc_hd__inv_2
X_4882_ _4931_/A _4882_/B vssd1 vssd1 vccd1 vccd1 _4882_/Y sky130_fd_sc_hd__nor2_1
X_3833_ _3837_/A _3833_/B vssd1 vssd1 vccd1 vccd1 _3833_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3764_ _3771_/A _3764_/B vssd1 vssd1 vccd1 vccd1 _3764_/Y sky130_fd_sc_hd__nand2_1
X_3695_ _3735_/A vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2715_ _2874_/A vssd1 vssd1 vccd1 vccd1 _2715_/Y sky130_fd_sc_hd__inv_2
X_2646_ _5270_/Q vssd1 vssd1 vccd1 vccd1 _2698_/A sky130_fd_sc_hd__inv_2
X_2577_ _3705_/A vssd1 vssd1 vccd1 vccd1 _2594_/A sky130_fd_sc_hd__clkbuf_2
X_4316_ _4316_/A _4316_/B vssd1 vssd1 vccd1 vccd1 _4316_/Y sky130_fd_sc_hd__nor2_1
X_4247_ _4247_/A _4574_/B vssd1 vssd1 vccd1 vccd1 _4249_/A sky130_fd_sc_hd__nand2_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4178_ _4185_/B _4178_/B vssd1 vssd1 vccd1 vccd1 _4178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ _3696_/B _5152_/Q vssd1 vssd1 vccd1 vccd1 _3130_/B sky130_fd_sc_hd__nand2_1
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3480_ _3777_/B _5122_/Q vssd1 vssd1 vccd1 vccd1 _3481_/B sky130_fd_sc_hd__nand2_1
X_2500_ _2516_/A _4702_/A vssd1 vssd1 vccd1 vccd1 _2500_/Y sky130_fd_sc_hd__nand2_1
XFILLER_69_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5150_ _5289_/CLK _5150_/D vssd1 vssd1 vccd1 vccd1 _5150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5081_ _5086_/CLK _5081_/D vssd1 vssd1 vccd1 vccd1 _5081_/Q sky130_fd_sc_hd__dfxtp_1
X_4101_ _5077_/Q vssd1 vssd1 vccd1 vccd1 _4210_/A sky130_fd_sc_hd__inv_2
X_4032_ _5058_/Q vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__inv_2
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4934_ _4934_/A vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__clkbuf_1
X_4865_ _4873_/A input4/X vssd1 vssd1 vccd1 vccd1 _4866_/A sky130_fd_sc_hd__or2_1
X_3816_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3816_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_4796_ _4796_/A vssd1 vssd1 vccd1 vccd1 _4803_/B sky130_fd_sc_hd__inv_2
X_3747_ _3758_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3747_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3678_ _3705_/A vssd1 vssd1 vccd1 vccd1 _3690_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2629_ _2745_/A _2835_/B vssd1 vssd1 vccd1 vccd1 _2629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5279_ _5282_/CLK hold2/X vssd1 vssd1 vccd1 vccd1 _5279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2980_ _3259_/A vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_21_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4650_ _4650_/A _4650_/B vssd1 vssd1 vccd1 vccd1 _4651_/B sky130_fd_sc_hd__nor2_1
Xinput21 phase_in[8] vssd1 vssd1 vccd1 vccd1 _4957_/D sky130_fd_sc_hd__clkbuf_1
Xinput10 oversample_in[8] vssd1 vssd1 vccd1 vccd1 _4853_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3601_ _3601_/A vssd1 vssd1 vccd1 vccd1 _3601_/X sky130_fd_sc_hd__clkbuf_2
X_4581_ _4991_/Q _5023_/Q vssd1 vssd1 vccd1 vccd1 _4828_/A sky130_fd_sc_hd__nand2_1
X_3532_ _3538_/B _3532_/B vssd1 vssd1 vccd1 vccd1 _3533_/B sky130_fd_sc_hd__nor2_1
X_3463_ _3548_/C _3463_/B vssd1 vssd1 vccd1 vccd1 _3551_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5202_ _5203_/CLK _5202_/D vssd1 vssd1 vccd1 vccd1 _5202_/Q sky130_fd_sc_hd__dfxtp_1
X_3394_ _5099_/Q _3837_/B _5194_/Q _3393_/Y vssd1 vssd1 vccd1 vccd1 _3657_/A sky130_fd_sc_hd__o2bb2ai_1
X_5133_ _5230_/CLK _5133_/D vssd1 vssd1 vccd1 vccd1 _5133_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5064_ _5064_/CLK _5064_/D vssd1 vssd1 vccd1 vccd1 _5064_/Q sky130_fd_sc_hd__dfxtp_1
X_4015_ _4033_/C _4015_/B vssd1 vssd1 vccd1 vccd1 _4016_/C sky130_fd_sc_hd__nand2_1
XFILLER_80_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4917_ _5094_/Q _4918_/A vssd1 vssd1 vccd1 vccd1 _4921_/C sky130_fd_sc_hd__or2_1
XFILLER_52_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4848_ _4848_/A vssd1 vssd1 vccd1 vccd1 _4988_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_20_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4779_ _4779_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4781_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2963_ _2963_/A _2963_/B _2963_/C vssd1 vssd1 vccd1 vccd1 _2963_/X sky130_fd_sc_hd__and3_1
XFILLER_15_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4702_ _4702_/A _4794_/B vssd1 vssd1 vccd1 vccd1 _4702_/Y sky130_fd_sc_hd__nand2_1
X_2894_ _2889_/A _2893_/Y _2850_/X vssd1 vssd1 vccd1 vccd1 _2894_/X sky130_fd_sc_hd__a21o_1
XFILLER_8_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4633_ _4748_/A _4748_/B _4753_/A vssd1 vssd1 vccd1 vccd1 _4634_/B sky130_fd_sc_hd__or3_1
X_4564_ _4779_/B vssd1 vssd1 vccd1 vccd1 _4564_/Y sky130_fd_sc_hd__inv_2
X_3515_ _3515_/A _3515_/B vssd1 vssd1 vccd1 vccd1 _3516_/B sky130_fd_sc_hd__nor2_1
X_4495_ _4500_/B _4500_/A vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__or2_1
X_3446_ _3583_/A _3583_/B _3590_/B vssd1 vssd1 vccd1 vccd1 _3446_/X sky130_fd_sc_hd__or3_1
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ _5111_/Q _3806_/B vssd1 vssd1 vccd1 vccd1 _3593_/A sky130_fd_sc_hd__nor2_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5116_ _5213_/CLK _5116_/D vssd1 vssd1 vccd1 vccd1 _5116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5047_ _5074_/CLK _5047_/D vssd1 vssd1 vccd1 vccd1 _5047_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3300_ _3300_/A vssd1 vssd1 vccd1 vccd1 _3301_/B sky130_fd_sc_hd__inv_2
X_4280_ _4476_/B _4476_/A _4481_/B vssd1 vssd1 vccd1 vccd1 _4280_/X sky130_fd_sc_hd__or3_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _3228_/Y _3230_/X _2839_/X vssd1 vssd1 vccd1 vccd1 _5212_/D sky130_fd_sc_hd__o21a_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3162_ _5159_/Q vssd1 vssd1 vccd1 vccd1 _3163_/B sky130_fd_sc_hd__inv_2
XFILLER_39_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _3093_/A _3093_/B vssd1 vssd1 vccd1 vccd1 _3262_/B sky130_fd_sc_hd__or2_1
XFILLER_81_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3995_ _3995_/A _3995_/B _3995_/C _3995_/D vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__or4_2
XFILLER_50_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2946_ _2945_/B _2945_/A _2912_/X vssd1 vssd1 vccd1 vccd1 _2946_/X sky130_fd_sc_hd__a21o_1
X_2877_ _2880_/C _2877_/B vssd1 vssd1 vccd1 vccd1 _2877_/Y sky130_fd_sc_hd__nand2_1
X_4616_ _4613_/A _4769_/B _4613_/B vssd1 vssd1 vccd1 vccd1 _4756_/B sky130_fd_sc_hd__o21ba_1
X_4547_ _4547_/A _4547_/B vssd1 vssd1 vccd1 vccd1 _4639_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4478_ _4478_/A _4478_/B _4478_/C vssd1 vssd1 vccd1 vccd1 _4478_/X sky130_fd_sc_hd__and3_1
X_3429_ _3429_/A _3429_/B vssd1 vssd1 vccd1 vccd1 _3430_/A sky130_fd_sc_hd__nor2_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3780_ _3784_/A _3780_/B vssd1 vssd1 vccd1 vccd1 _3780_/Y sky130_fd_sc_hd__nand2_1
X_2800_ _3505_/A _5256_/Q vssd1 vssd1 vccd1 vccd1 _2800_/Y sky130_fd_sc_hd__nand2_1
X_2731_ _5279_/Q _4547_/A vssd1 vssd1 vccd1 vccd1 _2731_/Y sky130_fd_sc_hd__nor2_1
X_4401_ _4406_/A _4406_/B _4335_/A vssd1 vssd1 vccd1 vccd1 _4402_/A sky130_fd_sc_hd__o21bai_1
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2662_ _2966_/B _4994_/Q _2977_/A _2968_/B vssd1 vssd1 vccd1 vccd1 _2963_/A sky130_fd_sc_hd__o22ai_2
X_2593_ _4994_/Q vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__inv_2
X_4332_ _4332_/A _4650_/B vssd1 vssd1 vccd1 vccd1 _4333_/B sky130_fd_sc_hd__nor2_1
X_4263_ _4263_/A _4263_/B vssd1 vssd1 vccd1 vccd1 _4497_/B sky130_fd_sc_hd__nor2_1
X_3214_ _5216_/Q _2928_/X _2962_/X _3213_/X vssd1 vssd1 vccd1 vccd1 _5216_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4194_ _5055_/Q _4195_/A vssd1 vssd1 vccd1 vccd1 _4196_/A sky130_fd_sc_hd__or2_1
X_3145_ _3196_/B _3145_/B vssd1 vssd1 vccd1 vccd1 _3181_/A sky130_fd_sc_hd__or2_1
XFILLER_67_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3076_ _3076_/A _3076_/B vssd1 vssd1 vccd1 vccd1 _3275_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3978_ _3937_/Y _3980_/A _3986_/A _3986_/C vssd1 vssd1 vccd1 vccd1 _3992_/A sky130_fd_sc_hd__a22oi_4
XFILLER_50_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2929_ _2929_/A _2929_/B vssd1 vssd1 vccd1 vccd1 _2929_/X sky130_fd_sc_hd__or2_1
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 oversample_in[6] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4950_ _4895_/X _4894_/B _4951_/S vssd1 vssd1 vccd1 vccd1 _4950_/X sky130_fd_sc_hd__mux2_1
X_4881_ _5096_/Q _4985_/Q vssd1 vssd1 vccd1 vccd1 _4881_/Y sky130_fd_sc_hd__nor2_1
X_3901_ _4986_/Q vssd1 vssd1 vccd1 vccd1 _3901_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3832_ _3832_/A vssd1 vssd1 vccd1 vccd1 _3832_/X sky130_fd_sc_hd__clkbuf_4
X_3763_ _3802_/A vssd1 vssd1 vccd1 vccd1 _3763_/X sky130_fd_sc_hd__clkbuf_2
X_3694_ _5153_/Q _3685_/X _3682_/X _3693_/Y vssd1 vssd1 vccd1 vccd1 _5153_/D sky130_fd_sc_hd__o211a_1
X_2714_ _2706_/B _2708_/A _5005_/Q _2704_/Y vssd1 vssd1 vccd1 vccd1 _2874_/A sky130_fd_sc_hd__a31o_1
X_2645_ _4612_/A _5271_/Q vssd1 vssd1 vccd1 vccd1 _2697_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4315_ _4445_/A _4445_/B _4450_/B vssd1 vssd1 vccd1 vccd1 _4316_/B sky130_fd_sc_hd__or3_1
X_2576_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__clkbuf_2
X_4246_ _5027_/Q vssd1 vssd1 vccd1 vccd1 _4574_/B sky130_fd_sc_hd__inv_2
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4177_ _4177_/A _4192_/B vssd1 vssd1 vccd1 vccd1 _4178_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3128_ _3135_/A vssd1 vssd1 vccd1 vccd1 _3208_/B sky130_fd_sc_hd__inv_2
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_82_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3059_ _3744_/B _5134_/Q vssd1 vssd1 vccd1 vccd1 _3060_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5080_ _5080_/CLK _5080_/D vssd1 vssd1 vccd1 vccd1 _5080_/Q sky130_fd_sc_hd__dfxtp_1
X_4100_ _4208_/A _4104_/B _4099_/Y vssd1 vssd1 vccd1 vccd1 _5078_/D sky130_fd_sc_hd__a21oi_1
X_4031_ _4033_/A _4017_/C _5057_/Q vssd1 vssd1 vccd1 vccd1 _4179_/A sky130_fd_sc_hd__a21o_1
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4933_ _4933_/A _4936_/B vssd1 vssd1 vccd1 vccd1 _4934_/A sky130_fd_sc_hd__and2_1
X_4864_ _4864_/A vssd1 vssd1 vccd1 vccd1 _4980_/D sky130_fd_sc_hd__clkbuf_1
X_3815_ _3815_/A vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__clkbuf_2
X_4795_ _3886_/X _4793_/Y _4784_/X _4794_/Y vssd1 vssd1 vccd1 vccd1 _4999_/D sky130_fd_sc_hd__o211a_1
X_3746_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3758_/A sky130_fd_sc_hd__clkbuf_2
X_3677_ _5159_/Q _3671_/X _3644_/X _3676_/Y vssd1 vssd1 vccd1 vccd1 _5159_/D sky130_fd_sc_hd__o211a_1
X_2628_ _2741_/A _2626_/Y _2741_/B vssd1 vssd1 vccd1 vccd1 _2835_/B sky130_fd_sc_hd__o21ba_1
X_2559_ _2573_/A _4607_/A vssd1 vssd1 vccd1 vccd1 _2559_/Y sky130_fd_sc_hd__nand2_1
X_5278_ _5278_/CLK _5278_/D vssd1 vssd1 vccd1 vccd1 _5278_/Q sky130_fd_sc_hd__dfxtp_1
X_4229_ _4229_/A vssd1 vssd1 vccd1 vccd1 _4457_/B sky130_fd_sc_hd__inv_2
XFILLER_75_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput22 phase_in[9] vssd1 vssd1 vccd1 vccd1 _4955_/D sky130_fd_sc_hd__clkbuf_1
Xinput11 oversample_in[9] vssd1 vssd1 vccd1 vccd1 _4851_/B sky130_fd_sc_hd__clkbuf_2
X_4580_ _4992_/Q _5024_/Q vssd1 vssd1 vccd1 vccd1 _4829_/B sky130_fd_sc_hd__nand2_1
X_3600_ _5175_/Q _3580_/X _3597_/Y _3599_/X _3587_/X vssd1 vssd1 vccd1 vccd1 _5175_/D
+ sky130_fd_sc_hd__o221a_1
X_3531_ _3531_/A _3531_/B vssd1 vssd1 vccd1 vccd1 _3534_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3462_ _3782_/B _5120_/Q vssd1 vssd1 vccd1 vccd1 _3463_/B sky130_fd_sc_hd__nand2_1
X_3393_ _5098_/Q vssd1 vssd1 vccd1 vccd1 _3393_/Y sky130_fd_sc_hd__inv_2
X_5201_ _5201_/CLK _5201_/D vssd1 vssd1 vccd1 vccd1 _5201_/Q sky130_fd_sc_hd__dfxtp_1
X_5132_ _5227_/CLK _5132_/D vssd1 vssd1 vccd1 vccd1 _5132_/Q sky130_fd_sc_hd__dfxtp_1
X_5063_ _5063_/CLK _5063_/D vssd1 vssd1 vccd1 vccd1 _5063_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4014_ _4020_/B _4009_/C _4009_/B vssd1 vssd1 vccd1 vccd1 _4033_/C sky130_fd_sc_hd__a21o_1
XFILLER_37_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4916_ _4916_/A vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__clkbuf_1
X_4847_ _4844_/Y _4847_/B _4847_/C vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__and3b_1
XFILLER_32_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4778_ _4785_/B _4785_/A vssd1 vssd1 vccd1 vccd1 _4781_/A sky130_fd_sc_hd__or2_1
X_3729_ _5140_/Q _3725_/X _3722_/X _3728_/Y vssd1 vssd1 vccd1 vccd1 _5140_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2962_ _3644_/A vssd1 vssd1 vccd1 vccd1 _2962_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4701_ _4701_/A vssd1 vssd1 vccd1 vccd1 _4794_/B sky130_fd_sc_hd__buf_2
XFILLER_30_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2893_ _2893_/A _2893_/B vssd1 vssd1 vccd1 vccd1 _2893_/Y sky130_fd_sc_hd__nand2_1
X_4632_ _4632_/A _4632_/B vssd1 vssd1 vccd1 vccd1 _4753_/A sky130_fd_sc_hd__nand2_1
X_4563_ _4782_/A _4563_/B vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__nor2_1
X_4494_ _4494_/A _4494_/B vssd1 vssd1 vccd1 vccd1 _4500_/A sky130_fd_sc_hd__and2_1
X_3514_ _3514_/A _3514_/B vssd1 vssd1 vccd1 vccd1 _3516_/A sky130_fd_sc_hd__nor2_1
X_3445_ _3585_/B _3445_/B vssd1 vssd1 vccd1 vccd1 _3590_/B sky130_fd_sc_hd__nand2_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _3806_/B _5111_/Q vssd1 vssd1 vccd1 vccd1 _3434_/A sky130_fd_sc_hd__nand2_1
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5115_ _5213_/CLK _5115_/D vssd1 vssd1 vccd1 vccd1 _5115_/Q sky130_fd_sc_hd__dfxtp_1
X_5046_ _5076_/CLK _5046_/D vssd1 vssd1 vccd1 vccd1 _5046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3230_ _3230_/A _3230_/B _3230_/C vssd1 vssd1 vccd1 vccd1 _3230_/X sky130_fd_sc_hd__and3_1
XFILLER_79_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _3157_/Y _3159_/Y _3160_/Y vssd1 vssd1 vccd1 vccd1 _5225_/D sky130_fd_sc_hd__a21oi_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3092_ _3723_/B _5142_/Q vssd1 vssd1 vccd1 vccd1 _3093_/B sky130_fd_sc_hd__and2_1
XFILLER_81_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3994_ _3994_/A _3995_/D vssd1 vssd1 vccd1 vccd1 _3994_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _2945_/A _2945_/B vssd1 vssd1 vccd1 vccd1 _2945_/Y sky130_fd_sc_hd__nor2_1
X_2876_ _2876_/A vssd1 vssd1 vccd1 vccd1 _2876_/Y sky130_fd_sc_hd__inv_2
X_4615_ _4767_/A _4767_/B _4614_/Y vssd1 vssd1 vccd1 vccd1 _4756_/A sky130_fd_sc_hd__o21bai_1
X_4546_ _4727_/B _4723_/A vssd1 vssd1 vccd1 vccd1 _4546_/Y sky130_fd_sc_hd__nor2_1
XFILLER_89_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4477_ _4478_/A _4478_/C _4478_/B vssd1 vssd1 vccd1 vccd1 _4477_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3428_ _3810_/B _5109_/Q vssd1 vssd1 vccd1 vccd1 _3429_/B sky130_fd_sc_hd__and2_1
XFILLER_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _3790_/B _5117_/Q vssd1 vssd1 vccd1 vccd1 _3370_/A sky130_fd_sc_hd__and2_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5029_ _5265_/CLK _5029_/D vssd1 vssd1 vccd1 vccd1 _5029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2730_ _2857_/B _2857_/A _2862_/B vssd1 vssd1 vccd1 vccd1 _2738_/B sky130_fd_sc_hd__or3_1
XFILLER_8_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2661_ _5260_/Q _4579_/A _2975_/A _2986_/B vssd1 vssd1 vccd1 vccd1 _2968_/B sky130_fd_sc_hd__a22oi_2
X_4400_ _4397_/X _4399_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5049_/D sky130_fd_sc_hd__a21oi_1
X_2592_ _5262_/Q _2584_/X _2585_/X _2591_/Y vssd1 vssd1 vccd1 vccd1 hold16/A sky130_fd_sc_hd__o211a_1
X_4331_ _5048_/Q vssd1 vssd1 vccd1 vccd1 _4650_/B sky130_fd_sc_hd__inv_2
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4262_ _4262_/A _4497_/C vssd1 vssd1 vccd1 vccd1 _4493_/A sky130_fd_sc_hd__and2_1
X_3213_ _3208_/A _3212_/Y _2930_/X vssd1 vssd1 vccd1 vccd1 _3213_/X sky130_fd_sc_hd__a21o_1
X_4193_ _4395_/A _4193_/B vssd1 vssd1 vccd1 vccd1 _4195_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3144_ _3144_/A vssd1 vssd1 vccd1 vccd1 _3145_/B sky130_fd_sc_hd__inv_2
X_3075_ _5234_/Q _5138_/Q vssd1 vssd1 vccd1 vccd1 _3282_/B sky130_fd_sc_hd__xor2_1
XFILLER_54_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3977_ _4001_/C _4000_/B _3979_/B vssd1 vssd1 vccd1 vccd1 _3986_/C sky130_fd_sc_hd__nand3_4
XFILLER_10_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2928_ _3601_/A vssd1 vssd1 vccd1 vccd1 _2928_/X sky130_fd_sc_hd__buf_2
XFILLER_50_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2859_ _2856_/X _2729_/A _2857_/Y _2603_/A vssd1 vssd1 vccd1 vccd1 _2859_/X sky130_fd_sc_hd__a31o_1
X_4529_ _4529_/A _4529_/B vssd1 vssd1 vccd1 vccd1 _4529_/X sky130_fd_sc_hd__or2_1
XFILLER_49_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 oversample_in[7] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_64_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4880_ _4880_/A _4880_/B _4880_/C vssd1 vssd1 vccd1 vccd1 _4887_/A sky130_fd_sc_hd__and3_1
X_3900_ _3898_/B _4982_/Q _5094_/Q _3899_/Y vssd1 vssd1 vccd1 vccd1 _3900_/X sky130_fd_sc_hd__a22o_1
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3831_ _5102_/Q _3819_/X _3829_/X _3830_/Y vssd1 vssd1 vccd1 vccd1 _5102_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3762_ _5128_/Q _3753_/X _3750_/X _3761_/Y vssd1 vssd1 vccd1 vccd1 _5128_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3693_ _3703_/A _3693_/B vssd1 vssd1 vccd1 vccd1 _3693_/Y sky130_fd_sc_hd__nand2_1
X_2713_ _2777_/A _2703_/Y _2712_/Y vssd1 vssd1 vccd1 vccd1 _2713_/Y sky130_fd_sc_hd__o21bai_1
X_2644_ _2644_/A _2644_/B _2643_/Y vssd1 vssd1 vccd1 vccd1 _2780_/A sky130_fd_sc_hd__or3b_1
X_2575_ _2836_/A vssd1 vssd1 vccd1 vccd1 _3718_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4314_ _4447_/B _4314_/B vssd1 vssd1 vccd1 vccd1 _4450_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4245_ _4258_/B _4259_/A vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__nor2_1
X_4176_ _5056_/Q _4176_/B vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__or2_1
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3127_ _5152_/Q _3696_/B vssd1 vssd1 vccd1 vccd1 _3135_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ _3058_/A vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__inv_2
XFILLER_82_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4030_ _4179_/B _4185_/B _4030_/C vssd1 vssd1 vccd1 vccd1 _4169_/D sky130_fd_sc_hd__nand3_2
XFILLER_37_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4932_ _4932_/A _4935_/B vssd1 vssd1 vccd1 vccd1 _4933_/A sky130_fd_sc_hd__nor2_1
X_4863_ _4873_/A input5/X vssd1 vssd1 vccd1 vccd1 _4864_/A sky130_fd_sc_hd__or2_1
X_3814_ _5108_/Q _3805_/X _3802_/X _3813_/Y vssd1 vssd1 vccd1 vccd1 _5108_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4794_ _4794_/A _4794_/B vssd1 vssd1 vccd1 vccd1 _4794_/Y sky130_fd_sc_hd__nand2_1
X_3745_ _5134_/Q _3739_/X _3735_/X _3744_/Y vssd1 vssd1 vccd1 vccd1 _5134_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3676_ _3676_/A _3676_/B vssd1 vssd1 vccd1 vccd1 _3676_/Y sky130_fd_sc_hd__nand2_1
X_2627_ _4650_/A _5283_/Q vssd1 vssd1 vccd1 vccd1 _2741_/B sky130_fd_sc_hd__and2_1
X_2558_ _5003_/Q vssd1 vssd1 vccd1 vccd1 _4607_/A sky130_fd_sc_hd__inv_2
XFILLER_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2489_ _5021_/Q vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__clkinv_2
X_5277_ _5278_/CLK _5277_/D vssd1 vssd1 vccd1 vccd1 _5277_/Q sky130_fd_sc_hd__dfxtp_1
X_4228_ _4294_/A _4556_/B vssd1 vssd1 vccd1 vccd1 _4229_/A sky130_fd_sc_hd__nor2_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4159_ _4159_/A vssd1 vssd1 vccd1 vccd1 _5061_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_55_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_35_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5215_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_62_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_26_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5259_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput12 phase_in[0] vssd1 vssd1 vccd1 vccd1 _4973_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 rst vssd1 vssd1 vccd1 vccd1 _4873_/A sky130_fd_sc_hd__buf_12
X_3530_ _3528_/Y _3529_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5188_/D sky130_fd_sc_hd__a21oi_1
X_3461_ _3475_/A vssd1 vssd1 vccd1 vccd1 _3548_/C sky130_fd_sc_hd__inv_2
XFILLER_6_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5200_ _5203_/CLK _5200_/D vssd1 vssd1 vccd1 vccd1 _5200_/Q sky130_fd_sc_hd__dfxtp_1
X_3392_ _5195_/Q vssd1 vssd1 vccd1 vccd1 _3837_/B sky130_fd_sc_hd__inv_2
X_5131_ _5227_/CLK _5131_/D vssd1 vssd1 vccd1 vccd1 _5131_/Q sky130_fd_sc_hd__dfxtp_1
X_5062_ _5063_/CLK _5062_/D vssd1 vssd1 vccd1 vccd1 _5062_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4013_ _3982_/X _4012_/Y _4027_/A _4026_/A _4022_/B vssd1 vssd1 vccd1 vccd1 _4016_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_65_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _5068_/CLK sky130_fd_sc_hd__clkbuf_16
X_4915_ _4915_/A _4915_/B vssd1 vssd1 vccd1 vccd1 _4916_/A sky130_fd_sc_hd__and2_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4846_ _4846_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4847_/C sky130_fd_sc_hd__nand2_1
XFILLER_32_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _4777_/A _4777_/B vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__and2_1
X_3728_ _3730_/A _3728_/B vssd1 vssd1 vccd1 vccd1 _3728_/Y sky130_fd_sc_hd__nand2_1
X_3659_ _5164_/Q _3634_/X _3656_/X _3658_/X _3642_/X vssd1 vssd1 vccd1 vccd1 _5164_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2961_ _4089_/A vssd1 vssd1 vccd1 vccd1 _3644_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_42_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4700_ _4655_/A _4705_/B _4662_/B vssd1 vssd1 vccd1 vccd1 _4700_/X sky130_fd_sc_hd__o21a_1
XFILLER_8_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2892_ _5243_/Q _2814_/X _2890_/Y _2891_/X _2822_/X vssd1 vssd1 vccd1 vccd1 _5243_/D
+ sky130_fd_sc_hd__o221a_1
X_4631_ _4754_/A _4631_/B vssd1 vssd1 vccd1 vccd1 _4632_/B sky130_fd_sc_hd__nand2_1
X_4562_ _5001_/Q _5033_/Q vssd1 vssd1 vccd1 vccd1 _4781_/C sky130_fd_sc_hd__nand2_1
X_4493_ _4493_/A vssd1 vssd1 vccd1 vccd1 _4500_/B sky130_fd_sc_hd__inv_2
X_3513_ _5222_/Q _3513_/B vssd1 vssd1 vccd1 vccd1 _3514_/B sky130_fd_sc_hd__nor2_1
X_3444_ _3803_/B _5112_/Q vssd1 vssd1 vccd1 vccd1 _3445_/B sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_6_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5278_/CLK sky130_fd_sc_hd__clkbuf_16
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3375_ _5207_/Q vssd1 vssd1 vccd1 vccd1 _3806_/B sky130_fd_sc_hd__inv_2
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _5213_/CLK _5114_/D vssd1 vssd1 vccd1 vccd1 _5114_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _5045_/CLK _5045_/D vssd1 vssd1 vccd1 vccd1 _5045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4829_ _4829_/A _4829_/B vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _5225_/Q _3668_/A _4115_/B vssd1 vssd1 vccd1 vccd1 _3160_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_66_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3091_ _3091_/A vssd1 vssd1 vccd1 vccd1 _3253_/B sky130_fd_sc_hd__inv_2
XFILLER_39_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_81_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3993_ _3993_/A _3993_/B vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__or2_1
X_2944_ _2944_/A vssd1 vssd1 vccd1 vccd1 _2945_/B sky130_fd_sc_hd__inv_2
X_2875_ _2890_/A _2893_/B _2893_/A vssd1 vssd1 vccd1 vccd1 _2875_/X sky130_fd_sc_hd__or3_1
X_4614_ _4774_/A _4766_/A vssd1 vssd1 vccd1 vccd1 _4614_/Y sky130_fd_sc_hd__nand2_1
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _4723_/A sky130_fd_sc_hd__inv_2
XFILLER_89_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4476_ _4476_/A _4476_/B vssd1 vssd1 vccd1 vccd1 _4478_/B sky130_fd_sc_hd__nor2_1
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3427_ _5109_/Q _3810_/B vssd1 vssd1 vccd1 vccd1 _3429_/A sky130_fd_sc_hd__nor2_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ _5117_/Q _3790_/B vssd1 vssd1 vccd1 vccd1 _3371_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3289_ _3288_/B _3288_/A _3244_/X vssd1 vssd1 vccd1 vccd1 _3289_/X sky130_fd_sc_hd__a21o_1
X_5028_ _5058_/CLK _5028_/D vssd1 vssd1 vccd1 vccd1 _5028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2660_ _2985_/B _4992_/Q vssd1 vssd1 vccd1 vccd1 _2986_/B sky130_fd_sc_hd__nand2_1
X_2591_ _2594_/A _4574_/A vssd1 vssd1 vccd1 vccd1 _2591_/Y sky130_fd_sc_hd__nand2_1
X_4330_ _5080_/Q _5048_/Q vssd1 vssd1 vccd1 vccd1 _4351_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4261_ _4261_/A _4589_/B vssd1 vssd1 vccd1 vccd1 _4262_/A sky130_fd_sc_hd__nand2_1
X_3212_ _3212_/A _3212_/B vssd1 vssd1 vccd1 vccd1 _3212_/Y sky130_fd_sc_hd__nand2_1
X_4192_ _4192_/A _4192_/B vssd1 vssd1 vccd1 vccd1 _4193_/B sky130_fd_sc_hd__nand2_1
XFILLER_27_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3143_ _3143_/A _3143_/B vssd1 vssd1 vccd1 vccd1 _3144_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3074_ _3071_/B _3287_/B _3071_/A vssd1 vssd1 vccd1 vccd1 _3276_/B sky130_fd_sc_hd__o21ba_1
XFILLER_39_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3976_ _3993_/A _3993_/B vssd1 vssd1 vccd1 vccd1 _3979_/B sky130_fd_sc_hd__nor2_1
XFILLER_10_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2927_ _5237_/Q _2907_/X _2924_/X _2926_/Y _2914_/X vssd1 vssd1 vccd1 vccd1 _5237_/D
+ sky130_fd_sc_hd__o221a_1
X_2858_ _2856_/X _2729_/A _2857_/Y vssd1 vssd1 vccd1 vccd1 _2858_/Y sky130_fd_sc_hd__a21oi_1
X_2789_ _2836_/A vssd1 vssd1 vccd1 vccd1 _2978_/A sky130_fd_sc_hd__buf_2
X_4528_ _5056_/Q _5024_/Q vssd1 vssd1 vccd1 vccd1 _4529_/A sky130_fd_sc_hd__nor2_1
X_4459_ _4987_/Q _5038_/Q _4456_/X _4458_/Y _4438_/X vssd1 vssd1 vccd1 vccd1 _5038_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_58_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _3837_/A _3830_/B vssd1 vssd1 vccd1 vccd1 _3830_/Y sky130_fd_sc_hd__nand2_1
X_3761_ _3771_/A _3761_/B vssd1 vssd1 vccd1 vccd1 _3761_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2712_ _2901_/A _2904_/A vssd1 vssd1 vccd1 vccd1 _2712_/Y sky130_fd_sc_hd__nand2_1
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3692_ _3705_/A vssd1 vssd1 vccd1 vccd1 _3703_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2643_ _2643_/A _2876_/A vssd1 vssd1 vccd1 vccd1 _2643_/Y sky130_fd_sc_hd__nand2_1
X_2574_ _5266_/Q _2564_/X _2565_/X _2573_/Y vssd1 vssd1 vccd1 vccd1 _5266_/D sky130_fd_sc_hd__o211a_1
X_4313_ _4313_/A _4631_/B vssd1 vssd1 vccd1 vccd1 _4314_/B sky130_fd_sc_hd__nand2_1
XFILLER_87_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4244_ _4244_/A _4572_/B vssd1 vssd1 vccd1 vccd1 _4259_/A sky130_fd_sc_hd__nor2_1
X_4175_ _4021_/Y _4016_/A _4023_/Y vssd1 vssd1 vccd1 vccd1 _4176_/B sky130_fd_sc_hd__o21a_1
XFILLER_67_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3126_ _5248_/Q vssd1 vssd1 vccd1 vccd1 _3696_/B sky130_fd_sc_hd__inv_2
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3057_ _5133_/Q _3747_/B vssd1 vssd1 vccd1 vccd1 _3058_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3959_ hold22/A vssd1 vssd1 vccd1 vccd1 _3961_/B sky130_fd_sc_hd__inv_2
XFILLER_2_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4931_ _4931_/A _4931_/B vssd1 vssd1 vccd1 vccd1 _4935_/B sky130_fd_sc_hd__nor2_1
X_4862_ _4862_/A vssd1 vssd1 vccd1 vccd1 _4981_/D sky130_fd_sc_hd__clkbuf_1
X_3813_ _3824_/A _3813_/B vssd1 vssd1 vccd1 vccd1 _3813_/Y sky130_fd_sc_hd__nand2_1
X_4793_ _4793_/A _4793_/B vssd1 vssd1 vccd1 vccd1 _4793_/Y sky130_fd_sc_hd__xnor2_1
X_3744_ _3744_/A _3744_/B vssd1 vssd1 vccd1 vccd1 _3744_/Y sky130_fd_sc_hd__nand2_1
X_3675_ _5160_/Q _3671_/X _3644_/X _3674_/Y vssd1 vssd1 vccd1 vccd1 _5160_/D sky130_fd_sc_hd__o211a_1
X_2626_ _5282_/Q hold15/A vssd1 vssd1 vccd1 vccd1 _2626_/Y sky130_fd_sc_hd__nor2_1
X_2557_ _2557_/A vssd1 vssd1 vccd1 vccd1 _2573_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_5276_ _5278_/CLK _5276_/D vssd1 vssd1 vccd1 vccd1 _5276_/Q sky130_fd_sc_hd__dfxtp_1
X_2488_ _2557_/A vssd1 vssd1 vccd1 vccd1 _2496_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_87_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4227_ _5037_/Q vssd1 vssd1 vccd1 vccd1 _4556_/B sky130_fd_sc_hd__inv_2
X_4158_ _4158_/A _4760_/A _4158_/C vssd1 vssd1 vccd1 vccd1 _4159_/A sky130_fd_sc_hd__and3_1
XFILLER_46_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4089_ _4089_/A vssd1 vssd1 vccd1 vccd1 _4093_/B sky130_fd_sc_hd__clkbuf_2
X_3109_ _3109_/A vssd1 vssd1 vccd1 vccd1 _3110_/B sky130_fd_sc_hd__inv_2
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 phase_in[10] vssd1 vssd1 vccd1 vccd1 _4953_/D sky130_fd_sc_hd__clkbuf_1
X_3460_ _5120_/Q _3782_/B vssd1 vssd1 vccd1 vccd1 _3475_/A sky130_fd_sc_hd__nor2_1
X_3391_ _5100_/Q _3835_/B vssd1 vssd1 vccd1 vccd1 _3655_/A sky130_fd_sc_hd__nor2_1
X_5130_ _5227_/CLK _5130_/D vssd1 vssd1 vccd1 vccd1 _5130_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5061_ _5063_/CLK _5061_/D vssd1 vssd1 vccd1 vccd1 _5061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4012_ _4020_/C _4012_/B vssd1 vssd1 vccd1 vccd1 _4012_/Y sky130_fd_sc_hd__nand2_1
XFILLER_80_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4914_ _4918_/A _4914_/B vssd1 vssd1 vccd1 vccd1 _4915_/B sky130_fd_sc_hd__nor2_1
X_4845_ _4989_/Q _4844_/Y _4839_/A _4847_/B vssd1 vssd1 vccd1 vccd1 _4989_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4776_ _5003_/Q _4987_/Q _4715_/X _4775_/X vssd1 vssd1 vccd1 vccd1 _5003_/D sky130_fd_sc_hd__o211a_1
X_3727_ _5141_/Q _3725_/X _3722_/X _3726_/Y vssd1 vssd1 vccd1 vccd1 _5141_/D sky130_fd_sc_hd__o211a_1
X_3658_ _3655_/A _3655_/B _3657_/X vssd1 vssd1 vccd1 vccd1 _3658_/X sky130_fd_sc_hd__o21ba_1
X_3589_ _3644_/A vssd1 vssd1 vccd1 vccd1 _3589_/X sky130_fd_sc_hd__clkbuf_2
X_2609_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2609_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_0_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5259_ _5259_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _5259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2960_ _2803_/X _2956_/Y _2957_/X _2808_/X _2959_/Y vssd1 vssd1 vccd1 vccd1 _5231_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_63_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2891_ _2890_/B _2890_/A _2603_/A vssd1 vssd1 vccd1 vccd1 _2891_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4630_ _4630_/A vssd1 vssd1 vccd1 vccd1 _4632_/A sky130_fd_sc_hd__inv_2
X_4561_ _5002_/Q _5034_/Q vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__nor2_1
X_4492_ _4987_/Q _5031_/Q _4469_/X _4491_/X vssd1 vssd1 vccd1 vccd1 _5031_/D sky130_fd_sc_hd__o211a_1
X_3512_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3512_/X sky130_fd_sc_hd__clkbuf_2
X_3443_ _5112_/Q _3803_/B vssd1 vssd1 vccd1 vccd1 _3585_/B sky130_fd_sc_hd__or2_1
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _5110_/Q _3808_/B vssd1 vssd1 vccd1 vccd1 _3436_/A sky130_fd_sc_hd__nor2_1
X_5113_ _5209_/CLK _5113_/D vssd1 vssd1 vccd1 vccd1 _5113_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5044_ _5076_/CLK _5044_/D vssd1 vssd1 vccd1 vccd1 _5044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _4828_/A vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__inv_2
X_4759_ _4759_/A _4759_/B vssd1 vssd1 vccd1 vccd1 _4759_/X sky130_fd_sc_hd__and2_1
XFILLER_0_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3090_ _3086_/B _3267_/B _3086_/A vssd1 vssd1 vccd1 vccd1 _3254_/B sky130_fd_sc_hd__o21ba_1
Xhold2 hold2/A vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_66_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3992_ _3992_/A _3992_/B vssd1 vssd1 vccd1 vccd1 _4007_/A sky130_fd_sc_hd__nor2_1
X_2943_ _2943_/A _2943_/B vssd1 vssd1 vccd1 vccd1 _2944_/A sky130_fd_sc_hd__nor2_1
X_2874_ _2874_/A _2874_/B vssd1 vssd1 vccd1 vccd1 _2893_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4613_ _4613_/A _4613_/B vssd1 vssd1 vccd1 vccd1 _4766_/A sky130_fd_sc_hd__nor2_1
X_4544_ _4552_/A _4544_/B vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4475_ _4481_/B _4481_/A vssd1 vssd1 vccd1 vccd1 _4478_/A sky130_fd_sc_hd__or2_1
X_3426_ _5205_/Q vssd1 vssd1 vccd1 vccd1 _3810_/B sky130_fd_sc_hd__inv_2
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3357_ _5213_/Q vssd1 vssd1 vccd1 vccd1 _3790_/B sky130_fd_sc_hd__inv_2
XFILLER_38_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ _5058_/CLK _5027_/D vssd1 vssd1 vccd1 vccd1 _5027_/Q sky130_fd_sc_hd__dfxtp_1
X_3288_ _3288_/A _3288_/B vssd1 vssd1 vccd1 vccd1 _3288_/Y sky130_fd_sc_hd__nor2_1
XFILLER_45_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _4995_/Q vssd1 vssd1 vccd1 vccd1 _4574_/A sky130_fd_sc_hd__inv_2
X_4260_ _5029_/Q vssd1 vssd1 vccd1 vccd1 _4589_/B sky130_fd_sc_hd__inv_2
XFILLER_86_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4191_ _4191_/A _4191_/B vssd1 vssd1 vccd1 vccd1 _4192_/A sky130_fd_sc_hd__nand2_1
X_3211_ _3207_/X _2496_/A _3208_/Y _3210_/Y vssd1 vssd1 vccd1 vccd1 _5217_/D sky130_fd_sc_hd__a31oi_1
X_3142_ _3142_/A _3142_/B vssd1 vssd1 vccd1 vccd1 _3196_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073_ _3047_/Y _3295_/A _3064_/Y _3072_/Y vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__o211ai_1
XFILLER_35_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3975_ _3975_/A _3994_/A _3975_/C vssd1 vssd1 vccd1 vccd1 _4000_/B sky130_fd_sc_hd__nand3_2
X_2926_ _2926_/A _2926_/B vssd1 vssd1 vccd1 vccd1 _2926_/Y sky130_fd_sc_hd__nor2_1
X_2857_ _2857_/A _2857_/B vssd1 vssd1 vccd1 vccd1 _2857_/Y sky130_fd_sc_hd__nor2_1
X_2788_ _2761_/C _2761_/B _2761_/A _2787_/Y vssd1 vssd1 vccd1 vccd1 _2788_/Y sky130_fd_sc_hd__o22ai_1
X_4527_ _4987_/Q _5025_/Q _4525_/Y _4526_/X _4511_/X vssd1 vssd1 vccd1 vccd1 _5025_/D
+ sky130_fd_sc_hd__o221a_1
X_4458_ _4458_/A _4458_/B vssd1 vssd1 vccd1 vccd1 _4458_/Y sky130_fd_sc_hd__nor2_1
X_3409_ _3824_/B _5104_/Q vssd1 vssd1 vccd1 vccd1 _3410_/B sky130_fd_sc_hd__nand2_1
X_4389_ _4396_/A _4396_/C vssd1 vssd1 vccd1 vccd1 _4391_/B sky130_fd_sc_hd__and2_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3760_ _3773_/A vssd1 vssd1 vccd1 vccd1 _3771_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2711_ _2711_/A vssd1 vssd1 vccd1 vccd1 _2904_/A sky130_fd_sc_hd__inv_2
X_3691_ _5154_/Q _3685_/X _3682_/X _3690_/Y vssd1 vssd1 vccd1 vccd1 _5154_/D sky130_fd_sc_hd__o211a_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2642_ _2639_/Y _2889_/B _2716_/B vssd1 vssd1 vccd1 vccd1 _2876_/A sky130_fd_sc_hd__a21oi_1
X_2573_ _2573_/A _4794_/A vssd1 vssd1 vccd1 vccd1 _2573_/Y sky130_fd_sc_hd__nand2_1
X_4312_ _4312_/A vssd1 vssd1 vccd1 vccd1 _4447_/B sky130_fd_sc_hd__inv_2
X_4243_ _5028_/Q vssd1 vssd1 vccd1 vccd1 _4572_/B sky130_fd_sc_hd__inv_2
XFILLER_87_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4174_ _4171_/Y _4173_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5058_/D sky130_fd_sc_hd__a21oi_1
XFILLER_67_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _5153_/Q _3693_/B vssd1 vssd1 vccd1 vccd1 _3206_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3056_ _5229_/Q vssd1 vssd1 vccd1 vccd1 _3747_/B sky130_fd_sc_hd__inv_2
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3958_ _3958_/A _3995_/C vssd1 vssd1 vccd1 vccd1 _3964_/A sky130_fd_sc_hd__nand2_1
X_3889_ _5089_/Q _3888_/Y _4890_/B _4978_/Q vssd1 vssd1 vccd1 vccd1 _3889_/X sky130_fd_sc_hd__o22a_1
X_2909_ _2916_/B vssd1 vssd1 vccd1 vccd1 _2917_/B sky130_fd_sc_hd__inv_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4930_ _5096_/Q _4930_/B vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__nor2_1
X_4861_ _4873_/A input6/X vssd1 vssd1 vccd1 vccd1 _4862_/A sky130_fd_sc_hd__or2_1
X_3812_ _3826_/A vssd1 vssd1 vccd1 vccd1 _3824_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4792_ _5000_/Q _4987_/Q _4790_/Y _4791_/X _4772_/X vssd1 vssd1 vccd1 vccd1 _5000_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3743_ _5135_/Q _3739_/X _3735_/X _3742_/Y vssd1 vssd1 vccd1 vccd1 _5135_/D sky130_fd_sc_hd__o211a_1
X_3674_ _3676_/A _3674_/B vssd1 vssd1 vccd1 vccd1 _3674_/Y sky130_fd_sc_hd__nand2_1
X_2625_ _5283_/Q _4650_/A vssd1 vssd1 vccd1 vccd1 _2741_/A sky130_fd_sc_hd__nor2_1
X_2556_ _5271_/Q _2544_/X _2547_/X _2555_/Y vssd1 vssd1 vccd1 vccd1 _5271_/D sky130_fd_sc_hd__o211a_1
X_2487_ _3738_/A vssd1 vssd1 vccd1 vccd1 _2557_/A sky130_fd_sc_hd__clkbuf_2
X_5275_ _5278_/CLK _5275_/D vssd1 vssd1 vccd1 vccd1 _5275_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4226_ _5070_/Q _5038_/Q vssd1 vssd1 vccd1 vccd1 _4455_/A sky130_fd_sc_hd__nor2_1
X_4157_ _4069_/A _4162_/C _4261_/A vssd1 vssd1 vccd1 vccd1 _4158_/C sky130_fd_sc_hd__o21ai_1
X_3108_ _3712_/B _5146_/Q vssd1 vssd1 vccd1 vccd1 _3109_/A sky130_fd_sc_hd__nand2_1
X_4088_ _4110_/A _4088_/B vssd1 vssd1 vccd1 vccd1 _4093_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3039_ _3093_/A _3091_/A _3253_/A vssd1 vssd1 vccd1 vccd1 _3240_/A sky130_fd_sc_hd__a21o_1
XFILLER_43_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 phase_in[1] vssd1 vssd1 vccd1 vccd1 _4971_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3390_ _5196_/Q vssd1 vssd1 vccd1 vccd1 _3835_/B sky130_fd_sc_hd__inv_2
X_5060_ _5063_/CLK _5060_/D vssd1 vssd1 vccd1 vccd1 _5060_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4011_ _4011_/A _4015_/B _4022_/B vssd1 vssd1 vccd1 vccd1 _4033_/A sky130_fd_sc_hd__nand3_2
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4913_ _5093_/Q _4913_/B vssd1 vssd1 vccd1 vccd1 _4914_/B sky130_fd_sc_hd__nor2_1
XFILLER_20_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4844_ _4846_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4844_/Y sky130_fd_sc_hd__nor2_1
X_4775_ _4774_/X _4769_/A _4501_/X vssd1 vssd1 vccd1 vccd1 _4775_/X sky130_fd_sc_hd__a21o_1
X_3726_ _3730_/A _3726_/B vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__nand2_1
X_3657_ _3657_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3657_/X sky130_fd_sc_hd__and2_1
X_3588_ _5177_/Q _3580_/X _3584_/X _3586_/Y _3587_/X vssd1 vssd1 vccd1 vccd1 _5177_/D
+ sky130_fd_sc_hd__o221a_1
X_2608_ _4992_/Q _2603_/X _2585_/X _2607_/Y vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__o211a_1
XFILLER_87_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2539_ _5275_/Q _2525_/X _2526_/X _2538_/Y vssd1 vssd1 vccd1 vccd1 _5275_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5258_ _5259_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _5258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4209_ _4212_/B vssd1 vssd1 vccd1 vccd1 _4209_/Y sky130_fd_sc_hd__inv_2
X_5189_ _5193_/CLK _5189_/D vssd1 vssd1 vccd1 vccd1 _5189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2890_ _2890_/A _2890_/B vssd1 vssd1 vccd1 vccd1 _2890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4560_ _4617_/A _4557_/Y _4617_/B vssd1 vssd1 vccd1 vccd1 _4737_/A sky130_fd_sc_hd__o21bai_1
X_4491_ _4486_/A _4490_/Y _4407_/X vssd1 vssd1 vccd1 vccd1 _4491_/X sky130_fd_sc_hd__a21o_1
X_3511_ _5191_/Q _3307_/X _3509_/Y _3510_/X _3315_/X vssd1 vssd1 vccd1 vccd1 _5191_/D
+ sky130_fd_sc_hd__o221a_1
X_3442_ _5208_/Q vssd1 vssd1 vccd1 vccd1 _3803_/B sky130_fd_sc_hd__inv_2
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ _5206_/Q vssd1 vssd1 vccd1 vccd1 _3808_/B sky130_fd_sc_hd__inv_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5112_ _5209_/CLK _5112_/D vssd1 vssd1 vccd1 vccd1 _5112_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5043_ _5045_/CLK _5043_/D vssd1 vssd1 vccd1 vccd1 _5043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_80_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _4993_/Q _4987_/Q _4824_/X _4826_/X _4772_/X vssd1 vssd1 vccd1 vccd1 _4993_/D
+ sky130_fd_sc_hd__o221a_1
X_4758_ _4759_/B _4759_/A vssd1 vssd1 vccd1 vccd1 _4758_/Y sky130_fd_sc_hd__nor2_1
X_4689_ _5020_/Q _4987_/Q _4686_/X _4688_/Y _4511_/X vssd1 vssd1 vccd1 vccd1 _5020_/D
+ sky130_fd_sc_hd__o221a_1
X_3709_ _3716_/A _3709_/B vssd1 vssd1 vccd1 vccd1 _3709_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_74_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3991_ _3986_/A _3986_/B _3986_/C _4012_/B vssd1 vssd1 vccd1 vccd1 _3992_/B sky130_fd_sc_hd__a31oi_4
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2942_ _2942_/A vssd1 vssd1 vccd1 vccd1 _2943_/B sky130_fd_sc_hd__inv_2
XFILLER_30_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2873_ _2603_/X _2870_/X _2609_/X _2872_/Y vssd1 vssd1 vccd1 vccd1 _5246_/D sky130_fd_sc_hd__o211a_1
X_4612_ _4612_/A _4612_/B vssd1 vssd1 vccd1 vccd1 _4613_/B sky130_fd_sc_hd__nor2_1
X_4543_ _4543_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4544_/B sky130_fd_sc_hd__nor2_1
X_4474_ _4474_/A _4474_/B vssd1 vssd1 vccd1 vccd1 _4481_/A sky130_fd_sc_hd__and2_1
X_3425_ _3607_/B _3425_/B vssd1 vssd1 vccd1 vccd1 _3611_/B sky130_fd_sc_hd__nand2_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3356_ _3345_/Y _3350_/X _3354_/Y _3354_/A _3355_/Y vssd1 vssd1 vccd1 vccd1 _3515_/A
+ sky130_fd_sc_hd__a311o_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _3287_/A _3287_/B vssd1 vssd1 vccd1 vccd1 _3288_/B sky130_fd_sc_hd__nand2_1
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _5265_/CLK _5026_/D vssd1 vssd1 vccd1 vccd1 _5026_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4190_ _4188_/Y _4189_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5056_/D sky130_fd_sc_hd__a21oi_1
XFILLER_5_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3210_ _5217_/Q _3528_/B _4144_/B vssd1 vssd1 vccd1 vccd1 _3210_/Y sky130_fd_sc_hd__o21ai_1
X_3141_ _3690_/B _5154_/Q vssd1 vssd1 vccd1 vccd1 _3142_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3072_ _3292_/B _3288_/A vssd1 vssd1 vccd1 vccd1 _3072_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3974_ _3994_/A _3975_/A _3972_/X _3973_/Y vssd1 vssd1 vccd1 vccd1 _4001_/C sky130_fd_sc_hd__o2bb2ai_2
XFILLER_50_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2925_ _2925_/A _2925_/B vssd1 vssd1 vccd1 vccd1 _2926_/B sky130_fd_sc_hd__and2_1
XFILLER_50_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2856_ _2862_/B _2862_/A vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__or2_1
X_2787_ _2755_/B _2755_/A _2797_/B _2797_/C vssd1 vssd1 vccd1 vccd1 _2787_/Y sky130_fd_sc_hd__a22oi_1
X_4526_ _4526_/A _4526_/B vssd1 vssd1 vccd1 vccd1 _4526_/X sky130_fd_sc_hd__and2_1
X_4457_ _4457_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4458_/B sky130_fd_sc_hd__and2_1
X_3408_ _5104_/Q _3824_/B vssd1 vssd1 vccd1 vccd1 _3626_/B sky130_fd_sc_hd__or2_1
X_4388_ _4406_/A _4406_/B _4347_/A vssd1 vssd1 vccd1 vccd1 _4396_/A sky130_fd_sc_hd__o21ai_1
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _5127_/Q _3764_/B vssd1 vssd1 vccd1 vccd1 _3507_/A sky130_fd_sc_hd__nor2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5009_ _5051_/CLK _5009_/D vssd1 vssd1 vccd1 vccd1 _5009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2710_ _2900_/B _2710_/B vssd1 vssd1 vccd1 vccd1 _2711_/A sky130_fd_sc_hd__nand2_1
X_3690_ _3690_/A _3690_/B vssd1 vssd1 vccd1 vccd1 _3690_/Y sky130_fd_sc_hd__nand2_1
X_2641_ _4628_/A _5275_/Q vssd1 vssd1 vccd1 vccd1 _2716_/B sky130_fd_sc_hd__and2_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2572_ _4999_/Q vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__inv_2
X_4311_ _4311_/A _4631_/B vssd1 vssd1 vccd1 vccd1 _4312_/A sky130_fd_sc_hd__nor2_1
X_4242_ _5060_/Q _5028_/Q vssd1 vssd1 vccd1 vccd1 _4258_/B sky130_fd_sc_hd__nor2_1
X_4173_ _4820_/B _5058_/Q vssd1 vssd1 vccd1 vccd1 _4173_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3124_ _3693_/B _5153_/Q vssd1 vssd1 vccd1 vccd1 _3206_/B sky130_fd_sc_hd__and2_1
XFILLER_82_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3055_ _5229_/Q _3048_/Y _3310_/A _3310_/B vssd1 vssd1 vccd1 vccd1 _3304_/A sky130_fd_sc_hd__o22ai_4
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3957_ _3957_/A _3995_/D vssd1 vssd1 vccd1 vccd1 _3958_/A sky130_fd_sc_hd__nand2_1
X_2908_ _2908_/A _2908_/B vssd1 vssd1 vccd1 vccd1 _2916_/B sky130_fd_sc_hd__nand2_1
X_3888_ _4979_/Q vssd1 vssd1 vccd1 vccd1 _3888_/Y sky130_fd_sc_hd__inv_2
X_2839_ _4849_/A vssd1 vssd1 vccd1 vccd1 _2839_/X sky130_fd_sc_hd__buf_6
X_4509_ _4509_/A _4509_/B vssd1 vssd1 vccd1 vccd1 _4509_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5254_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5227_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_17_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4860_ _4860_/A vssd1 vssd1 vccd1 vccd1 _4982_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_17_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3811_ _5109_/Q _3805_/X _3802_/X _3810_/Y vssd1 vssd1 vccd1 vccd1 _5109_/D sky130_fd_sc_hd__o211a_1
X_4791_ _4790_/B _4790_/A _4181_/X vssd1 vssd1 vccd1 vccd1 _4791_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3742_ _3744_/A _3742_/B vssd1 vssd1 vccd1 vccd1 _3742_/Y sky130_fd_sc_hd__nand2_1
X_3673_ _5161_/Q _3671_/X _3644_/X _3672_/Y vssd1 vssd1 vccd1 vccd1 _5161_/D sky130_fd_sc_hd__o211a_1
X_2624_ _2624_/A vssd1 vssd1 vccd1 vccd1 _2745_/A sky130_fd_sc_hd__inv_2
X_2555_ _2555_/A _4612_/A vssd1 vssd1 vccd1 vccd1 _2555_/Y sky130_fd_sc_hd__nand2_1
X_2486_ _2836_/A vssd1 vssd1 vccd1 vccd1 _3738_/A sky130_fd_sc_hd__clkbuf_2
X_5274_ _5278_/CLK _5274_/D vssd1 vssd1 vccd1 vccd1 _5274_/Q sky130_fd_sc_hd__dfxtp_1
X_4225_ _4225_/A vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__inv_2
X_4156_ _4151_/A _4151_/B _4158_/A _4240_/A _4873_/A vssd1 vssd1 vccd1 vccd1 _5062_/D
+ sky130_fd_sc_hd__a221oi_1
X_3107_ _3106_/Y _3100_/A _3101_/A vssd1 vssd1 vccd1 vccd1 _3221_/B sky130_fd_sc_hd__a21oi_1
XFILLER_28_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4087_ _4327_/A _4087_/B vssd1 vssd1 vccd1 vccd1 _4088_/B sky130_fd_sc_hd__nor2_1
XFILLER_70_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3038_ _5143_/Q _3720_/B vssd1 vssd1 vccd1 vccd1 _3253_/A sky130_fd_sc_hd__nor2_1
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4989_ _5137_/CLK _4989_/D vssd1 vssd1 vccd1 vccd1 _4989_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput15 phase_in[2] vssd1 vssd1 vccd1 vccd1 _4969_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4010_ _4020_/B _4018_/A _3992_/A _3992_/B vssd1 vssd1 vccd1 vccd1 _4022_/B sky130_fd_sc_hd__o2bb2ai_4
XFILLER_77_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4912_ _4912_/A _4912_/B vssd1 vssd1 vccd1 vccd1 _4918_/A sky130_fd_sc_hd__nor2_1
X_4843_ _4838_/Y _4839_/X _4847_/B vssd1 vssd1 vccd1 vccd1 _4990_/D sky130_fd_sc_hd__o21a_1
X_4774_ _4774_/A _4774_/B vssd1 vssd1 vccd1 vccd1 _4774_/X sky130_fd_sc_hd__or2_1
X_3725_ _3725_/A vssd1 vssd1 vccd1 vccd1 _3725_/X sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_9_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5045_/CLK sky130_fd_sc_hd__clkbuf_16
X_3656_ _3655_/Y _3663_/B _3657_/A _2809_/A vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__a31o_1
X_3587_ _4183_/A vssd1 vssd1 vccd1 vccd1 _3587_/X sky130_fd_sc_hd__clkbuf_2
X_2607_ _3199_/A _2985_/B vssd1 vssd1 vccd1 vccd1 _2607_/Y sky130_fd_sc_hd__nand2_1
X_2538_ _2555_/A _4628_/A vssd1 vssd1 vccd1 vccd1 _2538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5257_ _5289_/CLK _5257_/D vssd1 vssd1 vccd1 vccd1 _5257_/Q sky130_fd_sc_hd__dfxtp_1
X_4208_ _4208_/A _4543_/B vssd1 vssd1 vccd1 vccd1 _4212_/B sky130_fd_sc_hd__nor2_1
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5188_ _5193_/CLK _5188_/D vssd1 vssd1 vccd1 vccd1 _5188_/Q sky130_fd_sc_hd__dfxtp_1
X_4139_ _5067_/Q _4135_/A _4138_/X vssd1 vssd1 vccd1 vccd1 _5067_/D sky130_fd_sc_hd__o21a_1
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3510_ _3485_/Y _3488_/Y _3508_/Y _2803_/A vssd1 vssd1 vccd1 vccd1 _3510_/X sky130_fd_sc_hd__a31o_1
X_4490_ _4490_/A _4490_/B vssd1 vssd1 vccd1 vccd1 _4490_/Y sky130_fd_sc_hd__nand2_1
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3441_ _3800_/B _5113_/Q vssd1 vssd1 vccd1 vccd1 _3583_/B sky130_fd_sc_hd__and2_1
XFILLER_6_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ _3453_/A _3566_/B _3571_/B _3369_/Y _3371_/Y vssd1 vssd1 vccd1 vccd1 _3372_/Y
+ sky130_fd_sc_hd__o41ai_2
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5111_ _5209_/CLK _5111_/D vssd1 vssd1 vccd1 vccd1 _5111_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _5283_/CLK _5042_/D vssd1 vssd1 vccd1 vccd1 _5042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4826_ _4826_/A _4826_/B _4826_/C vssd1 vssd1 vccd1 vccd1 _4826_/X sky130_fd_sc_hd__and3_1
XFILLER_21_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4619_/A _4763_/B _4557_/Y vssd1 vssd1 vccd1 vccd1 _4759_/A sky130_fd_sc_hd__o21a_1
X_4688_ _4688_/A _4987_/Q vssd1 vssd1 vccd1 vccd1 _4688_/Y sky130_fd_sc_hd__nand2_1
X_3708_ _3735_/A vssd1 vssd1 vccd1 vccd1 _3708_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3639_ _3639_/A _3639_/B vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__nand2_1
XFILLER_88_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4 hold4/A vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_66_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3990_ _4026_/A _4027_/A _4026_/B vssd1 vssd1 vccd1 vccd1 _4192_/B sky130_fd_sc_hd__nand3_2
XFILLER_62_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2941_ _2603_/X _2938_/X _2903_/X _2940_/Y vssd1 vssd1 vccd1 vccd1 _5234_/D sky130_fd_sc_hd__o211a_1
XFILLER_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4611_ _5004_/Q _5036_/Q vssd1 vssd1 vccd1 vccd1 _4613_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2872_ _3199_/A _3701_/B vssd1 vssd1 vccd1 vccd1 _2872_/Y sky130_fd_sc_hd__nand2_1
X_4542_ _5014_/Q _5046_/Q vssd1 vssd1 vccd1 vccd1 _4552_/A sky130_fd_sc_hd__nor2_1
X_4473_ _4987_/Q _5035_/Q _4469_/X _4472_/Y vssd1 vssd1 vccd1 vccd1 _5035_/D sky130_fd_sc_hd__o211a_1
X_3424_ _3813_/B _5108_/Q vssd1 vssd1 vccd1 vccd1 _3425_/B sky130_fd_sc_hd__nand2_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3355_ _3355_/A _3355_/B vssd1 vssd1 vccd1 vccd1 _3355_/Y sky130_fd_sc_hd__nor2_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _3740_/B _5136_/Q _3292_/A vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__a21o_1
X_5025_ _5058_/CLK _5025_/D vssd1 vssd1 vccd1 vccd1 _5025_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4809_ _4810_/A _4810_/C _4810_/B vssd1 vssd1 vccd1 vccd1 _4809_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_79_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140_ _3186_/A _3140_/B vssd1 vssd1 vccd1 vccd1 _3146_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3071_ _3071_/A _3071_/B vssd1 vssd1 vccd1 vccd1 _3288_/A sky130_fd_sc_hd__or2_1
XFILLER_54_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _4968_/Q _3973_/B vssd1 vssd1 vccd1 vccd1 _3973_/Y sky130_fd_sc_hd__nor2_1
XFILLER_50_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2924_ _2925_/A _2926_/A _2925_/B _2898_/X vssd1 vssd1 vccd1 vccd1 _2924_/X sky130_fd_sc_hd__a31o_1
X_2855_ _2731_/Y _2854_/Y _2733_/B vssd1 vssd1 vccd1 vccd1 _2862_/A sky130_fd_sc_hd__o21ai_1
X_4525_ _4526_/B _4526_/A _4987_/Q vssd1 vssd1 vccd1 vccd1 _4525_/Y sky130_fd_sc_hd__o21ai_1
X_2786_ _2804_/A vssd1 vssd1 vccd1 vccd1 _2797_/C sky130_fd_sc_hd__inv_2
X_4456_ _4457_/A _4458_/A _4457_/B _3881_/A vssd1 vssd1 vccd1 vccd1 _4456_/X sky130_fd_sc_hd__a31o_1
X_4387_ _4535_/A vssd1 vssd1 vccd1 vccd1 _4387_/X sky130_fd_sc_hd__clkbuf_4
X_3407_ _5200_/Q vssd1 vssd1 vccd1 vccd1 _3824_/B sky130_fd_sc_hd__inv_2
X_3338_ _5223_/Q vssd1 vssd1 vccd1 vccd1 _3764_/B sky130_fd_sc_hd__inv_2
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3269_ _3268_/B _3268_/A _3244_/X vssd1 vssd1 vccd1 vccd1 _3269_/X sky130_fd_sc_hd__a21o_1
X_5008_ _5278_/CLK _5008_/D vssd1 vssd1 vccd1 vccd1 _5008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2640_ _5274_/Q _4754_/A vssd1 vssd1 vccd1 vccd1 _2889_/B sky130_fd_sc_hd__or2_1
X_2571_ _5267_/Q _2564_/X _2565_/X _2570_/Y vssd1 vssd1 vccd1 vccd1 _5267_/D sky130_fd_sc_hd__o211a_1
X_4310_ _5039_/Q vssd1 vssd1 vccd1 vccd1 _4631_/B sky130_fd_sc_hd__inv_2
X_4241_ _4263_/A _4497_/C _4263_/B vssd1 vssd1 vccd1 vccd1 _4484_/A sky130_fd_sc_hd__o21bai_1
X_4172_ _4701_/A vssd1 vssd1 vccd1 vccd1 _4820_/B sky130_fd_sc_hd__buf_2
X_3123_ _5249_/Q vssd1 vssd1 vccd1 vccd1 _3693_/B sky130_fd_sc_hd__inv_2
X_3054_ _3751_/B _5132_/Q _3318_/A _3326_/B vssd1 vssd1 vccd1 vccd1 _3310_/B sky130_fd_sc_hd__a22oi_4
XFILLER_27_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3956_ _3995_/C _3957_/A _3995_/D vssd1 vssd1 vccd1 vccd1 _3996_/A sky130_fd_sc_hd__nand3b_2
X_2907_ _3230_/B vssd1 vssd1 vccd1 vccd1 _2907_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3887_ _4983_/Q vssd1 vssd1 vccd1 vccd1 _3887_/Y sky130_fd_sc_hd__inv_2
X_2838_ _3815_/A vssd1 vssd1 vccd1 vccd1 _4849_/A sky130_fd_sc_hd__buf_6
X_2769_ _2656_/Y _2953_/A _2768_/X vssd1 vssd1 vccd1 vccd1 _2942_/A sky130_fd_sc_hd__o21bai_1
X_4508_ _5059_/Q _5027_/Q _4507_/X vssd1 vssd1 vccd1 vccd1 _4509_/B sky130_fd_sc_hd__a21o_1
X_4439_ _4987_/Q _5042_/Q _4435_/Y _4437_/X _4438_/X vssd1 vssd1 vccd1 vccd1 _5042_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4790_ _4790_/A _4790_/B vssd1 vssd1 vccd1 vccd1 _4790_/Y sky130_fd_sc_hd__nor2_1
X_3810_ _3810_/A _3810_/B vssd1 vssd1 vccd1 vccd1 _3810_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3741_ _5136_/Q _3739_/X _3735_/X _3740_/Y vssd1 vssd1 vccd1 vccd1 _5136_/D sky130_fd_sc_hd__o211a_1
XFILLER_9_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _3676_/A _3672_/B vssd1 vssd1 vccd1 vccd1 _3672_/Y sky130_fd_sc_hd__nand2_1
X_2623_ _2835_/A _2828_/B vssd1 vssd1 vccd1 vccd1 _2624_/A sky130_fd_sc_hd__nand2_1
X_2554_ _5004_/Q vssd1 vssd1 vccd1 vccd1 _4612_/A sky130_fd_sc_hd__inv_2
X_2485_ _4853_/A vssd1 vssd1 vccd1 vccd1 _2485_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5273_ _5288_/CLK _5273_/D vssd1 vssd1 vccd1 vccd1 _5273_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4224_ _4212_/A _4211_/A _4209_/Y _4223_/Y vssd1 vssd1 vccd1 vccd1 _4225_/A sky130_fd_sc_hd__o211a_1
X_4155_ _4163_/B _5061_/Q vssd1 vssd1 vccd1 vccd1 _4158_/A sky130_fd_sc_hd__nand2_1
X_3106_ _5144_/Q _3716_/B vssd1 vssd1 vccd1 vccd1 _3106_/Y sky130_fd_sc_hd__nor2_1
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4086_ _4086_/A vssd1 vssd1 vccd1 vccd1 _4110_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3037_ _3720_/B _5143_/Q vssd1 vssd1 vccd1 vccd1 _3091_/A sky130_fd_sc_hd__nand2_1
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4988_ _5201_/CLK _4988_/D vssd1 vssd1 vccd1 vccd1 _4988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3939_ _4970_/Q hold5/A vssd1 vssd1 vccd1 vccd1 _4003_/B sky130_fd_sc_hd__xor2_2
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 phase_in[3] vssd1 vssd1 vccd1 vccd1 _4967_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4911_ _4911_/A vssd1 vssd1 vccd1 vccd1 _4911_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_33_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4842_ _4846_/A _4952_/S _4103_/A vssd1 vssd1 vccd1 vccd1 _4847_/B sky130_fd_sc_hd__o21a_1
X_4773_ _5004_/Q _4987_/Q _4770_/Y _4771_/X _4772_/X vssd1 vssd1 vccd1 vccd1 _5004_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3724_ _5142_/Q _3711_/X _3722_/X _3723_/Y vssd1 vssd1 vccd1 vccd1 _5142_/D sky130_fd_sc_hd__o211a_1
X_3655_ _3655_/A _3655_/B vssd1 vssd1 vccd1 vccd1 _3655_/Y sky130_fd_sc_hd__nor2_1
X_2606_ _5259_/Q vssd1 vssd1 vccd1 vccd1 _2985_/B sky130_fd_sc_hd__inv_2
X_3586_ _3586_/A _3586_/B vssd1 vssd1 vccd1 vccd1 _3586_/Y sky130_fd_sc_hd__nor2_1
X_2537_ _5008_/Q vssd1 vssd1 vccd1 vccd1 _4628_/A sky130_fd_sc_hd__inv_2
XFILLER_87_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5256_ _5263_/CLK _5256_/D vssd1 vssd1 vccd1 vccd1 _5256_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4207_ _5046_/Q vssd1 vssd1 vccd1 vccd1 _4543_/B sky130_fd_sc_hd__inv_2
XFILLER_68_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5187_ _5195_/CLK _5187_/D vssd1 vssd1 vccd1 vccd1 _5187_/Q sky130_fd_sc_hd__dfxtp_1
X_4138_ _4283_/A _4144_/A _4849_/A vssd1 vssd1 vccd1 vccd1 _4138_/X sky130_fd_sc_hd__o21a_1
XFILLER_56_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4069_ _4069_/A _4069_/B _4162_/C vssd1 vssd1 vccd1 vccd1 _4086_/A sky130_fd_sc_hd__nor3_2
XFILLER_36_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3440_ _5113_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3583_/A sky130_fd_sc_hd__nor2_1
X_3371_ _3371_/A _3371_/B vssd1 vssd1 vccd1 vccd1 _3371_/Y sky130_fd_sc_hd__nor2_1
XFILLER_88_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5110_ _5209_/CLK _5110_/D vssd1 vssd1 vccd1 vccd1 _5110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5041_ _5051_/CLK _5041_/D vssd1 vssd1 vccd1 vccd1 _5041_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4825_ _4829_/A _4825_/B vssd1 vssd1 vccd1 vccd1 _4826_/A sky130_fd_sc_hd__nand2_1
X_4756_ _4756_/A _4756_/B vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__and2_1
X_4687_ _4687_/A _4687_/B _4690_/B _4687_/D vssd1 vssd1 vccd1 vccd1 _4688_/A sky130_fd_sc_hd__or4_1
X_3707_ _5148_/Q _3698_/X _3695_/X _3706_/Y vssd1 vssd1 vccd1 vccd1 _5148_/D sky130_fd_sc_hd__o211a_1
X_3638_ _3639_/A _3639_/B _3641_/A _2809_/A vssd1 vssd1 vccd1 vccd1 _3638_/X sky130_fd_sc_hd__a31o_1
X_3569_ _3567_/X _3568_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5180_/D sky130_fd_sc_hd__a21oi_1
XFILLER_88_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5239_ _5288_/CLK _5239_/D vssd1 vssd1 vccd1 vccd1 _5239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_83_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2940_ _3199_/A _3733_/B vssd1 vssd1 vccd1 vccd1 _2940_/Y sky130_fd_sc_hd__nand2_1
X_2871_ _5246_/Q vssd1 vssd1 vccd1 vccd1 _3701_/B sky130_fd_sc_hd__inv_2
X_4610_ _4610_/A vssd1 vssd1 vccd1 vccd1 _4774_/A sky130_fd_sc_hd__inv_2
X_4541_ _4541_/A _4551_/A vssd1 vssd1 vccd1 vccd1 _4727_/B sky130_fd_sc_hd__or2_1
X_4472_ _4470_/Y _4471_/X _4987_/Q vssd1 vssd1 vccd1 vccd1 _4472_/Y sky130_fd_sc_hd__o21ai_1
X_3423_ _5108_/Q _3813_/B vssd1 vssd1 vccd1 vccd1 _3607_/B sky130_fd_sc_hd__or2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _3354_/A _3355_/A vssd1 vssd1 vccd1 vccd1 _3354_/Y sky130_fd_sc_hd__nor2_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3285_ _3047_/Y _3295_/A _3064_/Y vssd1 vssd1 vccd1 vccd1 _3292_/A sky130_fd_sc_hd__o21ai_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _5058_/CLK _5024_/D vssd1 vssd1 vccd1 vccd1 _5024_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4808_ _4813_/B _4813_/A vssd1 vssd1 vccd1 vccd1 _4810_/A sky130_fd_sc_hd__nand2_1
XFILLER_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4739_ _4744_/B _4744_/A vssd1 vssd1 vccd1 vccd1 _4739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3070_ _3736_/B _5137_/Q vssd1 vssd1 vccd1 vccd1 _3071_/B sky130_fd_sc_hd__and2_1
XFILLER_54_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3972_ _3973_/B _4968_/Q vssd1 vssd1 vccd1 vccd1 _3972_/X sky130_fd_sc_hd__and2_1
X_2923_ _2929_/B _2929_/A vssd1 vssd1 vccd1 vccd1 _2925_/A sky130_fd_sc_hd__nand2_1
XFILLER_50_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2854_ _2870_/B _2854_/B vssd1 vssd1 vccd1 vccd1 _2854_/Y sky130_fd_sc_hd__nand2_1
X_2785_ _2751_/B _5020_/Q _2816_/A _2784_/Y vssd1 vssd1 vccd1 vccd1 _2797_/B sky130_fd_sc_hd__o22ai_2
X_4524_ _4524_/A _4524_/B vssd1 vssd1 vccd1 vccd1 _4526_/A sky130_fd_sc_hd__and2_1
XFILLER_7_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4455_ _4455_/A _4455_/B vssd1 vssd1 vccd1 vccd1 _4458_/A sky130_fd_sc_hd__nor2_1
X_4386_ _4987_/Q _5051_/Q _4384_/X _4385_/Y _4183_/X vssd1 vssd1 vccd1 vccd1 _5051_/D
+ sky130_fd_sc_hd__o221a_1
X_3406_ _3637_/A vssd1 vssd1 vccd1 vccd1 _3406_/Y sky130_fd_sc_hd__inv_2
X_3337_ _5224_/Q _5128_/Q vssd1 vssd1 vccd1 vccd1 _3502_/A sky130_fd_sc_hd__nor2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _3268_/A _3268_/B vssd1 vssd1 vccd1 vccd1 _3268_/Y sky130_fd_sc_hd__nor2_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3199_ _3199_/A _3777_/B vssd1 vssd1 vccd1 vccd1 _3199_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5007_ _5278_/CLK _5007_/D vssd1 vssd1 vccd1 vccd1 _5007_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_81_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _2573_/A _4598_/A vssd1 vssd1 vccd1 vccd1 _2570_/Y sky130_fd_sc_hd__nand2_1
X_4240_ _4240_/A _4569_/B vssd1 vssd1 vccd1 vccd1 _4263_/B sky130_fd_sc_hd__nor2_1
X_4171_ _4169_/X _4987_/Q _4171_/C vssd1 vssd1 vccd1 vccd1 _4171_/Y sky130_fd_sc_hd__nand3b_1
X_3122_ _3122_/A _3122_/B vssd1 vssd1 vccd1 vccd1 _3202_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3053_ _5131_/Q _5227_/Q vssd1 vssd1 vccd1 vccd1 _3326_/B sky130_fd_sc_hd__or2b_1
XFILLER_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3955_ _3954_/A _3954_/B _3954_/C vssd1 vssd1 vccd1 vccd1 _3995_/D sky130_fd_sc_hd__o21ai_2
X_2906_ _5240_/Q _2847_/X _2903_/X _2905_/X vssd1 vssd1 vccd1 vccd1 _5240_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3886_ _3886_/A vssd1 vssd1 vccd1 vccd1 _3886_/X sky130_fd_sc_hd__clkbuf_4
X_2837_ _2837_/A _3832_/A _2837_/C vssd1 vssd1 vccd1 vccd1 _2837_/X sky130_fd_sc_hd__and3_1
X_2768_ _2768_/A _2955_/B vssd1 vssd1 vccd1 vccd1 _2768_/X sky130_fd_sc_hd__or2_1
X_4507_ _4507_/A _4520_/C _4507_/C vssd1 vssd1 vccd1 vccd1 _4507_/X sky130_fd_sc_hd__and3_1
X_2699_ _4607_/A _5270_/Q vssd1 vssd1 vccd1 vccd1 _2700_/B sky130_fd_sc_hd__nand2_1
X_4438_ _4772_/A vssd1 vssd1 vccd1 vccd1 _4438_/X sky130_fd_sc_hd__buf_2
X_4369_ _4369_/A _4369_/B _4987_/Q vssd1 vssd1 vccd1 vccd1 _4369_/Y sky130_fd_sc_hd__nand3_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_73_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3740_ _3744_/A _3740_/B vssd1 vssd1 vccd1 vccd1 _3740_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3671_ _3725_/A vssd1 vssd1 vccd1 vccd1 _3671_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2622_ _2630_/A _2622_/B vssd1 vssd1 vccd1 vccd1 _2828_/B sky130_fd_sc_hd__nor2_1
X_2553_ _5272_/Q _2544_/X _2547_/X hold14/X vssd1 vssd1 vccd1 vccd1 _5272_/D sky130_fd_sc_hd__o211a_1
X_2484_ _3815_/A vssd1 vssd1 vccd1 vccd1 _4853_/A sky130_fd_sc_hd__clkbuf_2
X_5272_ _5272_/CLK _5272_/D vssd1 vssd1 vccd1 vccd1 _5272_/Q sky130_fd_sc_hd__dfxtp_1
X_4223_ _4324_/A _4223_/B vssd1 vssd1 vccd1 vccd1 _4223_/Y sky130_fd_sc_hd__nand2_1
X_4154_ _4151_/Y _4267_/A _4153_/X vssd1 vssd1 vccd1 vccd1 _5063_/D sky130_fd_sc_hd__a21oi_1
X_4085_ _4873_/A _4085_/B _4085_/C vssd1 vssd1 vccd1 vccd1 _5081_/D sky130_fd_sc_hd__nor3_1
X_3105_ _5240_/Q vssd1 vssd1 vccd1 vccd1 _3716_/B sky130_fd_sc_hd__inv_2
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3036_ _5239_/Q vssd1 vssd1 vccd1 vccd1 _3720_/B sky130_fd_sc_hd__inv_2
XFILLER_55_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4987_ _5201_/CLK _4987_/D vssd1 vssd1 vccd1 vccd1 _4987_/Q sky130_fd_sc_hd__dfxtp_4
X_3938_ _3938_/A hold21/A vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__nand2_1
X_3869_ _5092_/Q vssd1 vssd1 vccd1 vccd1 _3898_/B sky130_fd_sc_hd__inv_2
XFILLER_3_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput17 phase_in[4] vssd1 vssd1 vccd1 vccd1 _4965_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4910_ _4915_/A _4910_/B vssd1 vssd1 vccd1 vccd1 _4911_/A sky130_fd_sc_hd__and2_1
XFILLER_33_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4841_ _4841_/A _4872_/A vssd1 vssd1 vccd1 vccd1 _4952_/S sky130_fd_sc_hd__nor2_1
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4772_ _4772_/A vssd1 vssd1 vccd1 vccd1 _4772_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3723_ _3730_/A _3723_/B vssd1 vssd1 vccd1 vccd1 _3723_/Y sky130_fd_sc_hd__nand2_1
X_3654_ _3835_/B _5100_/Q vssd1 vssd1 vccd1 vccd1 _3655_/B sky130_fd_sc_hd__and2_1
X_2605_ _2809_/A vssd1 vssd1 vccd1 vccd1 _3199_/A sky130_fd_sc_hd__clkbuf_4
X_3585_ _3585_/A _3585_/B vssd1 vssd1 vccd1 vccd1 _3586_/B sky130_fd_sc_hd__and2_1
X_2536_ _2557_/A vssd1 vssd1 vccd1 vccd1 _2555_/A sky130_fd_sc_hd__clkbuf_2
X_5255_ _5259_/CLK _5255_/D vssd1 vssd1 vccd1 vccd1 _5255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4206_ _4415_/B vssd1 vssd1 vccd1 vccd1 _4211_/A sky130_fd_sc_hd__inv_2
XFILLER_68_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5186_ _5195_/CLK _5186_/D vssd1 vssd1 vccd1 vccd1 _5186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4135_/Y _4288_/A _4136_/Y vssd1 vssd1 vccd1 vccd1 _5068_/D sky130_fd_sc_hd__a21oi_1
XFILLER_56_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4068_ _4068_/A vssd1 vssd1 vccd1 vccd1 _4069_/B sky130_fd_sc_hd__inv_2
XFILLER_73_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3019_ hold25/A _5148_/Q vssd1 vssd1 vccd1 vccd1 _3020_/B sky130_fd_sc_hd__nand2_1
XFILLER_24_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3370_ _3370_/A _3370_/B vssd1 vssd1 vccd1 vccd1 _3371_/B sky130_fd_sc_hd__nor2_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _5051_/CLK _5040_/D vssd1 vssd1 vccd1 vccd1 _5040_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4824_ _4822_/Y _4829_/A _4825_/B _3881_/A vssd1 vssd1 vccd1 vccd1 _4824_/X sky130_fd_sc_hd__a31o_1
X_4755_ _3886_/X _4753_/X _4715_/X _4754_/Y vssd1 vssd1 vccd1 vccd1 _5007_/D sky130_fd_sc_hd__o211a_1
X_3706_ _3716_/A hold25/X vssd1 vssd1 vccd1 vccd1 _3706_/Y sky130_fd_sc_hd__nand2_1
X_4686_ _4687_/A _4687_/B _4690_/B _4687_/D vssd1 vssd1 vccd1 vccd1 _4686_/X sky130_fd_sc_hd__o22a_1
X_3637_ _3637_/A _3637_/B vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__nor2_1
X_3568_ _3568_/A _5180_/Q vssd1 vssd1 vccd1 vccd1 _3568_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2519_ _5013_/Q vssd1 vssd1 vccd1 vccd1 _4726_/B sky130_fd_sc_hd__clkinv_2
XFILLER_0_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3499_ _5127_/Q vssd1 vssd1 vccd1 vccd1 _3500_/B sky130_fd_sc_hd__inv_2
X_5238_ _5254_/CLK _5238_/D vssd1 vssd1 vccd1 vccd1 _5238_/Q sky130_fd_sc_hd__dfxtp_1
X_5169_ _5203_/CLK _5169_/D vssd1 vssd1 vccd1 vccd1 _5169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold6 hold6/A vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2870_ _2869_/X _2870_/B vssd1 vssd1 vccd1 vccd1 _2870_/X sky130_fd_sc_hd__and2b_1
XFILLER_90_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_10_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5076_/CLK sky130_fd_sc_hd__clkbuf_16
X_4540_ _4726_/B _4540_/B vssd1 vssd1 vccd1 vccd1 _4551_/A sky130_fd_sc_hd__nor2_1
X_4471_ _4471_/A _4471_/B vssd1 vssd1 vccd1 vccd1 _4471_/X sky130_fd_sc_hd__and2_1
X_3422_ _5204_/Q vssd1 vssd1 vccd1 vccd1 _3813_/B sky130_fd_sc_hd__inv_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _3769_/B _5125_/Q vssd1 vssd1 vccd1 vccd1 _3355_/A sky130_fd_sc_hd__and2_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3284_ _5202_/Q _3261_/X _3247_/X _3283_/X vssd1 vssd1 vccd1 vccd1 _5202_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _5058_/CLK _5023_/D vssd1 vssd1 vccd1 vccd1 _5023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4807_ _4807_/A _4819_/C vssd1 vssd1 vccd1 vccd1 _4813_/B sky130_fd_sc_hd__and2_1
X_2999_ _5158_/Q vssd1 vssd1 vccd1 vccd1 _3174_/B sky130_fd_sc_hd__inv_2
X_4738_ _4634_/B _4753_/B _4636_/Y vssd1 vssd1 vccd1 vccd1 _4744_/B sky130_fd_sc_hd__o21ai_1
X_4669_ _4692_/A _4692_/B _4690_/A vssd1 vssd1 vccd1 vccd1 _4687_/D sky130_fd_sc_hd__a21oi_1
XFILLER_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3971_ _4968_/D vssd1 vssd1 vccd1 vccd1 _3973_/B sky130_fd_sc_hd__inv_2
XFILLER_62_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2922_ _2922_/A _2922_/B vssd1 vssd1 vccd1 vccd1 _2929_/B sky130_fd_sc_hd__nand2_1
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2853_ _2869_/A _2869_/B _2869_/C vssd1 vssd1 vccd1 vccd1 _2870_/B sky130_fd_sc_hd__a21o_1
X_2784_ _5286_/Q hold24/A _2818_/A _2818_/B vssd1 vssd1 vccd1 vccd1 _2784_/Y sky130_fd_sc_hd__a22oi_1
X_4523_ _4529_/B _4523_/B vssd1 vssd1 vccd1 vccd1 _4526_/B sky130_fd_sc_hd__nor2_1
X_4454_ _4460_/B _4460_/A vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__or2_1
X_4385_ _4381_/Y _4383_/X _4382_/Y _4987_/Q vssd1 vssd1 vccd1 vccd1 _4385_/Y sky130_fd_sc_hd__o31ai_1
X_3405_ _5199_/Q _3405_/B vssd1 vssd1 vccd1 vccd1 _3637_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3336_ _5224_/Q _5128_/Q vssd1 vssd1 vccd1 vccd1 _3502_/B sky130_fd_sc_hd__and2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _3267_/A _3267_/B vssd1 vssd1 vccd1 vccd1 _3268_/B sky130_fd_sc_hd__nand2_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _5272_/CLK _5006_/D vssd1 vssd1 vccd1 vccd1 _5006_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3198_ _5218_/Q vssd1 vssd1 vccd1 vccd1 _3777_/B sky130_fd_sc_hd__inv_2
XFILLER_38_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _4179_/A _4169_/D _4169_/A _4169_/B vssd1 vssd1 vccd1 vccd1 _4171_/C sky130_fd_sc_hd__a22o_1
XFILLER_67_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3121_ _3701_/B _5150_/Q vssd1 vssd1 vccd1 vccd1 _3122_/B sky130_fd_sc_hd__nand2_1
XFILLER_67_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3052_ _5131_/Q _3754_/B _5226_/Q _3051_/Y vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3954_ _3954_/A _3954_/B _3954_/C vssd1 vssd1 vccd1 vccd1 _3957_/A sky130_fd_sc_hd__or3_1
XFILLER_16_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3885_ _3867_/X _4951_/X _3868_/X _3884_/Y vssd1 vssd1 vccd1 vccd1 _5088_/D sky130_fd_sc_hd__o211a_1
X_2905_ _2904_/X _2900_/A _2850_/X vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__a21o_1
X_2836_ _2836_/A vssd1 vssd1 vccd1 vccd1 _3832_/A sky130_fd_sc_hd__clkbuf_4
X_2767_ _2767_/A vssd1 vssd1 vccd1 vccd1 _2955_/B sky130_fd_sc_hd__inv_2
X_4506_ _4506_/A _4806_/B vssd1 vssd1 vccd1 vccd1 _4520_/C sky130_fd_sc_hd__nand2_1
X_2698_ _2698_/A _5003_/Q vssd1 vssd1 vccd1 vccd1 _2700_/A sky130_fd_sc_hd__nand2_1
X_4437_ _4435_/B _4435_/A _4436_/X vssd1 vssd1 vccd1 vccd1 _4437_/X sky130_fd_sc_hd__a21o_1
XFILLER_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4368_ _4200_/Y _4368_/B _4368_/C vssd1 vssd1 vccd1 vccd1 _4369_/B sky130_fd_sc_hd__nand3b_1
XFILLER_76_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4299_ _4299_/A _4637_/B vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3319_ _3319_/A vssd1 vssd1 vccd1 vccd1 _3319_/Y sky130_fd_sc_hd__inv_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3670_ _3738_/A vssd1 vssd1 vccd1 vccd1 _3725_/A sky130_fd_sc_hd__clkbuf_2
X_2621_ _2621_/A vssd1 vssd1 vccd1 vccd1 _2835_/A sky130_fd_sc_hd__inv_2
X_2552_ _2555_/A _4764_/A vssd1 vssd1 vccd1 vccd1 hold14/A sky130_fd_sc_hd__nand2_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5271_ _5288_/CLK _5271_/D vssd1 vssd1 vccd1 vccd1 _5271_/Q sky130_fd_sc_hd__dfxtp_1
X_4222_ _4217_/Y _4410_/A _4321_/A vssd1 vssd1 vccd1 vccd1 _4223_/B sky130_fd_sc_hd__a21oi_1
X_2483_ _2791_/A vssd1 vssd1 vccd1 vccd1 _3815_/A sky130_fd_sc_hd__clkbuf_4
X_4153_ _4074_/X _4075_/X _4141_/C _4873_/A vssd1 vssd1 vccd1 vccd1 _4153_/X sky130_fd_sc_hd__a31o_1
XFILLER_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4084_ _4074_/X _4075_/X _4057_/X _4080_/A _5081_/Q vssd1 vssd1 vccd1 vccd1 _4085_/B
+ sky130_fd_sc_hd__a41oi_1
X_3104_ _3240_/A _3240_/B _3103_/Y vssd1 vssd1 vccd1 vccd1 _3221_/A sky130_fd_sc_hd__o21bai_1
X_3035_ _5142_/Q _3723_/B vssd1 vssd1 vccd1 vccd1 _3093_/A sky130_fd_sc_hd__nor2_1
XFILLER_70_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4986_ _5281_/CLK _4986_/D vssd1 vssd1 vccd1 vccd1 _4986_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3937_ _3981_/A vssd1 vssd1 vccd1 vccd1 _3937_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3868_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3868_/X sky130_fd_sc_hd__clkbuf_2
X_3799_ _3826_/A vssd1 vssd1 vccd1 vccd1 _3810_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2819_ _2819_/A _2819_/B vssd1 vssd1 vccd1 vccd1 _2819_/Y sky130_fd_sc_hd__nor2_1
XFILLER_11_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_74_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput18 phase_in[5] vssd1 vssd1 vccd1 vccd1 _4963_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_6_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4840_ _4840_/A _4846_/B _4990_/Q vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__and3_1
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4771_ _4770_/B _4770_/A _4181_/X vssd1 vssd1 vccd1 vccd1 _4771_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3722_ _3735_/A vssd1 vssd1 vccd1 vccd1 _3722_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_9_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3653_ _5165_/Q _3634_/X _3651_/Y _3652_/X _3642_/X vssd1 vssd1 vccd1 vccd1 _5165_/D
+ sky130_fd_sc_hd__o221a_1
X_2604_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2809_/A sky130_fd_sc_hd__buf_2
X_3584_ _3585_/A _3586_/A _3585_/B _2898_/X vssd1 vssd1 vccd1 vccd1 _3584_/X sky130_fd_sc_hd__a31o_1
X_2535_ _5276_/Q _2525_/X _2526_/X _2534_/Y vssd1 vssd1 vccd1 vccd1 _5276_/D sky130_fd_sc_hd__o211a_1
X_5254_ _5254_/CLK _5254_/D vssd1 vssd1 vccd1 vccd1 _5254_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_87_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4205_ _4210_/A _4540_/B vssd1 vssd1 vccd1 vccd1 _4415_/B sky130_fd_sc_hd__nor2_1
X_5185_ _5195_/CLK _5185_/D vssd1 vssd1 vccd1 vccd1 _5185_/Q sky130_fd_sc_hd__dfxtp_1
X_4136_ _4129_/B _4144_/A _4093_/B vssd1 vssd1 vccd1 vccd1 _4136_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_3_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4067_ _5085_/Q _4065_/Y _4066_/Y vssd1 vssd1 vccd1 vccd1 _5085_/D sky130_fd_sc_hd__o21a_1
XFILLER_71_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3018_ _5148_/Q hold25/A vssd1 vssd1 vccd1 vccd1 _3032_/B sky130_fd_sc_hd__or2_1
XFILLER_24_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4969_ _5070_/CLK _4969_/D vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__dfxtp_1
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4823_ _4823_/A vssd1 vssd1 vccd1 vccd1 _4829_/A sky130_fd_sc_hd__inv_2
X_4754_ _4754_/A _4754_/B vssd1 vssd1 vccd1 vccd1 _4754_/Y sky130_fd_sc_hd__nand2_1
X_3705_ _3705_/A vssd1 vssd1 vccd1 vccd1 _3716_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4685_ _5020_/Q _5052_/Q vssd1 vssd1 vccd1 vccd1 _4687_/B sky130_fd_sc_hd__nor2_1
X_3636_ _5103_/Q _3827_/B vssd1 vssd1 vccd1 vccd1 _3637_/B sky130_fd_sc_hd__nor2_1
X_3567_ _3577_/A _3567_/B _3567_/C vssd1 vssd1 vccd1 vccd1 _3567_/X sky130_fd_sc_hd__or3_1
X_2518_ _2557_/A vssd1 vssd1 vccd1 vccd1 _2534_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3498_ _3494_/Y _3496_/Y _3497_/Y vssd1 vssd1 vccd1 vccd1 _5193_/D sky130_fd_sc_hd__a21oi_1
X_5237_ _5259_/CLK _5237_/D vssd1 vssd1 vccd1 vccd1 _5237_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5168_ _5168_/CLK _5168_/D vssd1 vssd1 vccd1 vccd1 _5168_/Q sky130_fd_sc_hd__dfxtp_1
X_4119_ _5073_/Q _4121_/C _4118_/Y vssd1 vssd1 vccd1 vccd1 _5073_/D sky130_fd_sc_hd__o21a_1
X_5099_ _5201_/CLK _5099_/D vssd1 vssd1 vccd1 vccd1 _5099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_35_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4470_ _4471_/B _4471_/A vssd1 vssd1 vccd1 vccd1 _4470_/Y sky130_fd_sc_hd__nor2_1
X_3421_ _3615_/A _3615_/B _3420_/X vssd1 vssd1 vccd1 vccd1 _3605_/B sky130_fd_sc_hd__a21oi_1
X_3352_ _5125_/Q _3769_/B vssd1 vssd1 vccd1 vccd1 _3354_/A sky130_fd_sc_hd__nor2_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _3277_/X _3282_/Y _3272_/X vssd1 vssd1 vccd1 vccd1 _3283_/X sky130_fd_sc_hd__a21o_1
X_5022_ _5070_/CLK _5022_/D vssd1 vssd1 vccd1 vccd1 hold4/A sky130_fd_sc_hd__dfxtp_2
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_80_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ hold7/A _4806_/B vssd1 vssd1 vccd1 vccd1 _4819_/C sky130_fd_sc_hd__nand2_1
X_2998_ _5159_/Q _3676_/B vssd1 vssd1 vccd1 vccd1 _3170_/A sky130_fd_sc_hd__nor2_1
X_4737_ _4737_/A _4737_/B vssd1 vssd1 vccd1 vccd1 _4753_/B sky130_fd_sc_hd__nor2_1
X_4668_ _5019_/Q _5051_/Q vssd1 vssd1 vccd1 vccd1 _4690_/A sky130_fd_sc_hd__nor2_1
X_3619_ _3618_/B _3618_/A _3598_/X vssd1 vssd1 vccd1 vccd1 _3619_/X sky130_fd_sc_hd__a21o_1
X_4599_ _4599_/A _4599_/B vssd1 vssd1 vccd1 vccd1 _4790_/A sky130_fd_sc_hd__or2_1
XFILLER_88_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3970_ _3993_/A _3993_/B _3968_/Y _3969_/X vssd1 vssd1 vccd1 vccd1 _3986_/A sky130_fd_sc_hd__o22ai_4
X_2921_ _5238_/Q _2847_/X _2903_/X _2920_/Y vssd1 vssd1 vccd1 vccd1 _5238_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2852_ _5250_/Q _2847_/X _2609_/X _2851_/X vssd1 vssd1 vccd1 vccd1 _5250_/D sky130_fd_sc_hd__o211a_1
X_2783_ _2783_/A vssd1 vssd1 vccd1 vccd1 _2818_/B sky130_fd_sc_hd__inv_2
X_4522_ _4516_/X _4519_/Y _4520_/X _4424_/X _4521_/Y vssd1 vssd1 vccd1 vccd1 _5026_/D
+ sky130_fd_sc_hd__o311a_1
X_4453_ _4453_/A _4453_/B vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__and2_1
X_3404_ _5103_/Q vssd1 vssd1 vccd1 vccd1 _3405_/B sky130_fd_sc_hd__inv_2
X_4384_ _4381_/Y _4382_/Y _4383_/X vssd1 vssd1 vccd1 vccd1 _4384_/X sky130_fd_sc_hd__o21a_1
X_3335_ _3495_/A vssd1 vssd1 vccd1 vccd1 _3335_/Y sky130_fd_sc_hd__inv_2
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3266_ _3271_/B _3271_/A vssd1 vssd1 vccd1 vccd1 _3267_/A sky130_fd_sc_hd__or2_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _5278_/CLK _5005_/D vssd1 vssd1 vccd1 vccd1 _5005_/Q sky130_fd_sc_hd__dfxtp_1
X_3197_ _3197_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3197_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _5150_/Q _3701_/B vssd1 vssd1 vccd1 vccd1 _3122_/A sky130_fd_sc_hd__or2_1
XFILLER_82_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3051_ _5130_/Q vssd1 vssd1 vccd1 vccd1 _3051_/Y sky130_fd_sc_hd__inv_2
XFILLER_75_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3953_ _4972_/Q _4972_/D vssd1 vssd1 vccd1 vccd1 _3954_/C sky130_fd_sc_hd__xnor2_2
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3884_ _4479_/A _4890_/B vssd1 vssd1 vccd1 vccd1 _3884_/Y sky130_fd_sc_hd__nand2_1
X_2904_ _2904_/A _2904_/B vssd1 vssd1 vccd1 vccd1 _2904_/X sky130_fd_sc_hd__or2_1
X_2835_ _2835_/A _2835_/B _2835_/C vssd1 vssd1 vccd1 vccd1 _2837_/A sky130_fd_sc_hd__or3_1
X_2766_ _2908_/B vssd1 vssd1 vccd1 vccd1 _2766_/Y sky130_fd_sc_hd__inv_2
X_4505_ _5026_/Q vssd1 vssd1 vccd1 vccd1 _4806_/B sky130_fd_sc_hd__inv_2
X_2697_ _2647_/Y _2697_/B vssd1 vssd1 vccd1 vccd1 _2911_/A sky130_fd_sc_hd__and2b_1
X_4436_ _4501_/A vssd1 vssd1 vccd1 vccd1 _4436_/X sky130_fd_sc_hd__buf_2
X_4367_ _4360_/Y _4373_/A _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4368_/B sky130_fd_sc_hd__o2bb2ai_1
XFILLER_86_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3318_ _3318_/A _3326_/B vssd1 vssd1 vccd1 vccd1 _3319_/A sky130_fd_sc_hd__and2_1
XFILLER_86_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4298_ _5041_/Q vssd1 vssd1 vccd1 vccd1 _4637_/B sky130_fd_sc_hd__inv_2
XFILLER_58_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3249_ _3241_/X _3248_/Y _2930_/X vssd1 vssd1 vccd1 vccd1 _3249_/X sky130_fd_sc_hd__a21o_1
XFILLER_39_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _2828_/C _2620_/B vssd1 vssd1 vccd1 vccd1 _2621_/A sky130_fd_sc_hd__nand2_1
X_2551_ _5005_/Q vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__inv_2
X_2482_ _4873_/A vssd1 vssd1 vccd1 vccd1 _2791_/A sky130_fd_sc_hd__inv_2
X_5270_ _5288_/CLK _5270_/D vssd1 vssd1 vccd1 vccd1 _5270_/Q sky130_fd_sc_hd__dfxtp_1
X_4221_ _5076_/Q _5044_/Q vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__nor2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4152_ _5063_/Q vssd1 vssd1 vccd1 vccd1 _4267_/A sky130_fd_sc_hd__inv_2
XFILLER_68_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4083_ _5082_/Q _4085_/C _4082_/Y vssd1 vssd1 vccd1 vccd1 _5082_/D sky130_fd_sc_hd__o21a_1
X_3103_ _3103_/A vssd1 vssd1 vccd1 vccd1 _3103_/Y sky130_fd_sc_hd__inv_2
X_3034_ _5238_/Q vssd1 vssd1 vccd1 vccd1 _3723_/B sky130_fd_sc_hd__inv_2
XFILLER_55_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4985_ _5281_/CLK _4985_/D vssd1 vssd1 vccd1 vccd1 _4985_/Q sky130_fd_sc_hd__dfxtp_1
X_3936_ hold21/A _3938_/A vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3867_ _3886_/A vssd1 vssd1 vccd1 vccd1 _3867_/X sky130_fd_sc_hd__clkbuf_2
X_3798_ _5114_/Q _3792_/X _3789_/X _3797_/Y vssd1 vssd1 vccd1 vccd1 _5114_/D sky130_fd_sc_hd__o211a_1
X_2818_ _2818_/A _2818_/B vssd1 vssd1 vccd1 vccd1 _2819_/B sky130_fd_sc_hd__nand2_1
X_2749_ _2816_/A vssd1 vssd1 vccd1 vccd1 _2806_/B sky130_fd_sc_hd__inv_2
XFILLER_78_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4419_ _4987_/Q _4540_/B _4415_/C _4418_/X vssd1 vssd1 vccd1 vccd1 _4420_/B sky130_fd_sc_hd__o22a_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 phase_in[6] vssd1 vssd1 vccd1 vccd1 _4961_/D sky130_fd_sc_hd__clkbuf_1
XFILLER_77_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4770_ _4770_/A _4770_/B vssd1 vssd1 vccd1 vccd1 _4770_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3721_ _5143_/Q _3711_/X _3708_/X _3720_/Y vssd1 vssd1 vccd1 vccd1 hold12/A sky130_fd_sc_hd__o211a_1
XFILLER_9_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3652_ _3651_/B _3651_/A _3598_/X vssd1 vssd1 vccd1 vccd1 _3652_/X sky130_fd_sc_hd__a21o_1
X_3583_ _3583_/A _3583_/B vssd1 vssd1 vccd1 vccd1 _3586_/A sky130_fd_sc_hd__nor2_1
X_2603_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2603_/X sky130_fd_sc_hd__buf_2
X_2534_ _2534_/A _4637_/A vssd1 vssd1 vccd1 vccd1 _2534_/Y sky130_fd_sc_hd__nand2_1
X_5253_ _5287_/CLK _5253_/D vssd1 vssd1 vccd1 vccd1 _5253_/Q sky130_fd_sc_hd__dfxtp_1
X_4204_ _5045_/Q vssd1 vssd1 vccd1 vccd1 _4540_/B sky130_fd_sc_hd__inv_2
X_5184_ _5195_/CLK _5184_/D vssd1 vssd1 vccd1 vccd1 _5184_/Q sky130_fd_sc_hd__dfxtp_1
X_4135_ _4135_/A _5067_/Q vssd1 vssd1 vccd1 vccd1 _4135_/Y sky130_fd_sc_hd__nand2_1
XFILLER_3_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4066_ _4151_/A _4057_/X _4058_/X _3931_/A _4873_/A vssd1 vssd1 vccd1 vccd1 _4066_/Y
+ sky130_fd_sc_hd__a41oi_1
XFILLER_71_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3017_ _5244_/Q vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__inv_2
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4968_ _5064_/CLK _4968_/D vssd1 vssd1 vccd1 vccd1 _4968_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3919_ _4311_/A vssd1 vssd1 vccd1 vccd1 _4313_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4899_ _4915_/A _4899_/B vssd1 vssd1 vccd1 vccd1 _4900_/A sky130_fd_sc_hd__and2_1
XFILLER_22_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_88_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4822_ _4826_/C _4826_/B vssd1 vssd1 vccd1 vccd1 _4822_/Y sky130_fd_sc_hd__nand2_1
X_4753_ _4753_/A _4753_/B vssd1 vssd1 vccd1 vccd1 _4753_/X sky130_fd_sc_hd__xor2_1
X_3704_ _5149_/Q _3698_/X _3695_/X _3703_/Y vssd1 vssd1 vccd1 vccd1 hold23/A sky130_fd_sc_hd__o211a_1
X_4684_ _4682_/X _4683_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5021_/D sky130_fd_sc_hd__a21oi_1
X_3635_ _3635_/A vssd1 vssd1 vccd1 vccd1 _3639_/A sky130_fd_sc_hd__inv_2
X_3566_ _3566_/A _3566_/B vssd1 vssd1 vccd1 vccd1 _3567_/C sky130_fd_sc_hd__and2_1
X_3497_ _5193_/Q _2979_/B _4115_/B vssd1 vssd1 vccd1 vccd1 _3497_/Y sky130_fd_sc_hd__o21ai_1
X_2517_ _5281_/Q _2506_/X _2507_/X _2516_/Y vssd1 vssd1 vccd1 vccd1 _5281_/D sky130_fd_sc_hd__o211a_1
X_5236_ _5254_/CLK _5236_/D vssd1 vssd1 vccd1 vccd1 _5236_/Q sky130_fd_sc_hd__dfxtp_1
X_5167_ _5168_/CLK _5167_/D vssd1 vssd1 vccd1 vccd1 _5167_/Q sky130_fd_sc_hd__dfxtp_1
X_4118_ _4130_/B _4113_/X _4873_/A vssd1 vssd1 vccd1 vccd1 _4118_/Y sky130_fd_sc_hd__a21oi_1
X_5098_ _5201_/CLK _5098_/D vssd1 vssd1 vccd1 vccd1 _5098_/Q sky130_fd_sc_hd__dfxtp_1
X_4049_ _4126_/A _4049_/B _4151_/B vssd1 vssd1 vccd1 vccd1 _4068_/A sky130_fd_sc_hd__and3_1
XFILLER_56_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold8 hold8/A vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__clkdlybuf4s50_1
XFILLER_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3420_ _3621_/B _3614_/A vssd1 vssd1 vccd1 vccd1 _3420_/X sky130_fd_sc_hd__or2_1
X_3351_ _5221_/Q vssd1 vssd1 vccd1 vccd1 _3769_/B sky130_fd_sc_hd__inv_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _3282_/A _3282_/B vssd1 vssd1 vccd1 vccd1 _3282_/Y sky130_fd_sc_hd__nand2_1
X_5021_ _5070_/CLK _5021_/D vssd1 vssd1 vccd1 vccd1 _5021_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4805_ _4997_/Q _4987_/Q _4784_/X _4804_/X vssd1 vssd1 vccd1 vccd1 _4997_/D sky130_fd_sc_hd__o211a_1
XFILLER_21_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2997_ _5256_/Q _5160_/Q vssd1 vssd1 vccd1 vccd1 _3165_/A sky130_fd_sc_hd__nor2_1
X_4736_ _3886_/X _4734_/Y _4715_/X _4735_/Y vssd1 vssd1 vccd1 vccd1 _5011_/D sky130_fd_sc_hd__o211a_1
X_4667_ _4663_/B _4665_/X _4660_/B _4666_/Y vssd1 vssd1 vccd1 vccd1 _4692_/B sky130_fd_sc_hd__a211oi_1
X_3618_ _3618_/A _3618_/B vssd1 vssd1 vccd1 vccd1 _3618_/Y sky130_fd_sc_hd__nor2_1
X_4598_ _4598_/A _4598_/B vssd1 vssd1 vccd1 vccd1 _4599_/B sky130_fd_sc_hd__nor2_1
X_3549_ _5185_/Q _3528_/B _4849_/A vssd1 vssd1 vccd1 vccd1 _3549_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_0_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5219_ _5219_/CLK _5219_/D vssd1 vssd1 vccd1 vccd1 _5219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2920_ _2916_/Y _2917_/Y _4940_/A vssd1 vssd1 vccd1 vccd1 _2920_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2851_ _2848_/X _2843_/A _2850_/X vssd1 vssd1 vccd1 vccd1 _2851_/X sky130_fd_sc_hd__a21o_1
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2782_ _2765_/Y _2781_/Y _2745_/Y vssd1 vssd1 vccd1 vccd1 _2818_/A sky130_fd_sc_hd__o21bai_1
X_4521_ _4754_/B _4806_/B vssd1 vssd1 vccd1 vccd1 _4521_/Y sky130_fd_sc_hd__nand2_1
X_4452_ _4987_/Q _5039_/Q _3907_/X _4451_/X vssd1 vssd1 vccd1 vccd1 _5039_/D sky130_fd_sc_hd__o211a_1
X_3403_ _3645_/A _3649_/A _3645_/B vssd1 vssd1 vccd1 vccd1 _3635_/A sky130_fd_sc_hd__a21oi_2
X_4383_ _4383_/A _4383_/B vssd1 vssd1 vccd1 vccd1 _4383_/X sky130_fd_sc_hd__or2_1
X_3334_ _5128_/Q _3761_/B vssd1 vssd1 vccd1 vccd1 _3495_/A sky130_fd_sc_hd__nor2_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _3265_/A _3265_/B vssd1 vssd1 vccd1 vccd1 _3271_/A sky130_fd_sc_hd__nor2_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5004_ _5272_/CLK _5004_/D vssd1 vssd1 vccd1 vccd1 _5004_/Q sky130_fd_sc_hd__dfxtp_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _3196_/A _3196_/B _3196_/C vssd1 vssd1 vccd1 vccd1 _3197_/A sky130_fd_sc_hd__and3_1
XFILLER_38_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4719_ _4719_/A _4719_/B vssd1 vssd1 vccd1 vccd1 _4734_/B sky130_fd_sc_hd__and2_1
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3050_ _5132_/Q _3751_/B vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__nor2_2
XFILLER_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3952_ _4974_/Q hold20/A vssd1 vssd1 vccd1 vccd1 _3954_/B sky130_fd_sc_hd__and2_1
XFILLER_16_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2903_ _2903_/A vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_3883_ _3883_/A vssd1 vssd1 vccd1 vccd1 _4890_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2834_ _3686_/B _3228_/B vssd1 vssd1 vccd1 vccd1 _2834_/Y sky130_fd_sc_hd__nor2_1
X_4504_ _4504_/A vssd1 vssd1 vccd1 vccd1 _4509_/A sky130_fd_sc_hd__inv_2
X_2765_ _2824_/B vssd1 vssd1 vccd1 vccd1 _2765_/Y sky130_fd_sc_hd__inv_2
X_2696_ _2692_/B _2925_/B _2695_/Y vssd1 vssd1 vccd1 vccd1 _2908_/B sky130_fd_sc_hd__o21a_1
X_4435_ _4435_/A _4435_/B vssd1 vssd1 vccd1 vccd1 _4435_/Y sky130_fd_sc_hd__nor2_1
X_4366_ _4200_/Y _4364_/Y _4368_/C vssd1 vssd1 vccd1 vccd1 _4369_/A sky130_fd_sc_hd__o21bai_1
XFILLER_86_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3317_ _3751_/B _5132_/Q vssd1 vssd1 vccd1 vccd1 _3317_/X sky130_fd_sc_hd__and2_1
XFILLER_86_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4297_ _4453_/A _4453_/B _4296_/X vssd1 vssd1 vccd1 vccd1 _4431_/B sky130_fd_sc_hd__a21oi_2
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3248_ _3248_/A _3248_/B vssd1 vssd1 vccd1 vccd1 _3248_/Y sky130_fd_sc_hd__nand2_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3179_ _5222_/Q _2972_/X _3177_/X _3178_/Y _2980_/X vssd1 vssd1 vccd1 vccd1 _5222_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_39_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _5273_/Q _2544_/X _2547_/X _2549_/Y vssd1 vssd1 vccd1 vccd1 _5273_/D sky130_fd_sc_hd__o211a_1
X_2481_ _3528_/B vssd1 vssd1 vccd1 vccd1 _2481_/X sky130_fd_sc_hd__clkbuf_2
X_4220_ _4421_/A vssd1 vssd1 vccd1 vccd1 _4410_/A sky130_fd_sc_hd__inv_2
XFILLER_68_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4151_ _4151_/A _4151_/B vssd1 vssd1 vccd1 vccd1 _4151_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4082_ _4130_/B _4058_/X _4873_/A vssd1 vssd1 vccd1 vccd1 _4082_/Y sky130_fd_sc_hd__a21oi_1
X_3102_ _3248_/B _3243_/A vssd1 vssd1 vccd1 vccd1 _3103_/A sky130_fd_sc_hd__and2b_1
X_3033_ _3025_/Y _3031_/X _3023_/A _3032_/Y vssd1 vssd1 vccd1 vccd1 _3201_/A sky130_fd_sc_hd__a211o_1
XFILLER_36_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4984_ _4984_/CLK _4984_/D vssd1 vssd1 vccd1 vccd1 _4984_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_63_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3935_ _4960_/Q vssd1 vssd1 vccd1 vccd1 _3938_/A sky130_fd_sc_hd__inv_2
X_3866_ _3844_/X _4946_/X _3845_/X _3865_/Y vssd1 vssd1 vccd1 vccd1 _5093_/D sky130_fd_sc_hd__o211a_1
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3797_ _3797_/A _3797_/B vssd1 vssd1 vccd1 vccd1 _3797_/Y sky130_fd_sc_hd__nand2_1
X_2817_ _2817_/A vssd1 vssd1 vccd1 vccd1 _2819_/A sky130_fd_sc_hd__inv_2
X_2748_ _5286_/Q hold24/A vssd1 vssd1 vccd1 vccd1 _2816_/A sky130_fd_sc_hd__nor2_1
X_4418_ _4413_/B _4413_/A _4501_/A vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__a21o_1
X_2679_ _2669_/A _4997_/Q _2933_/B _2771_/A vssd1 vssd1 vccd1 vccd1 _2679_/Y sky130_fd_sc_hd__a31oi_1
XFILLER_86_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4349_ _4349_/A vssd1 vssd1 vccd1 vccd1 _4349_/Y sky130_fd_sc_hd__inv_2
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3720_ _3730_/A _3720_/B vssd1 vssd1 vccd1 vccd1 _3720_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_40_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5209_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3651_ _3651_/A _3651_/B vssd1 vssd1 vccd1 vccd1 _3651_/Y sky130_fd_sc_hd__nor2_1
X_3582_ _3590_/B _3590_/A vssd1 vssd1 vccd1 vccd1 _3585_/A sky130_fd_sc_hd__or2_1
X_2602_ _2898_/A vssd1 vssd1 vccd1 vccd1 _2603_/A sky130_fd_sc_hd__clkbuf_4
X_2533_ _5009_/Q vssd1 vssd1 vccd1 vccd1 _4637_/A sky130_fd_sc_hd__inv_2
X_5252_ _5289_/CLK _5252_/D vssd1 vssd1 vccd1 vccd1 _5252_/Q sky130_fd_sc_hd__dfxtp_1
X_4203_ _5078_/Q _5046_/Q vssd1 vssd1 vccd1 vccd1 _4212_/A sky130_fd_sc_hd__nor2_1
X_5183_ _5195_/CLK _5183_/D vssd1 vssd1 vccd1 vccd1 _5183_/Q sky130_fd_sc_hd__dfxtp_1
X_4134_ _4141_/A _4141_/B _4134_/C vssd1 vssd1 vccd1 vccd1 _4135_/A sky130_fd_sc_hd__and3_1
XFILLER_68_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _4087_/B _4065_/B _4065_/C vssd1 vssd1 vccd1 vccd1 _4065_/Y sky130_fd_sc_hd__nor3_1
X_3016_ _3186_/B _3140_/B _3186_/A _3010_/A _3015_/Y vssd1 vssd1 vccd1 vccd1 _3016_/X
+ sky130_fd_sc_hd__a311o_2
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4967_ _5064_/CLK _4967_/D vssd1 vssd1 vccd1 vccd1 _4968_/D sky130_fd_sc_hd__dfxtp_1
X_3918_ _5071_/Q vssd1 vssd1 vccd1 vccd1 _4311_/A sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_31_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5195_/CLK sky130_fd_sc_hd__clkbuf_16
X_4898_ _5090_/Q _4891_/B _4902_/B vssd1 vssd1 vccd1 vccd1 _4899_/B sky130_fd_sc_hd__o21a_1
X_3849_ _3897_/B _4754_/B vssd1 vssd1 vccd1 vccd1 _3849_/Y sky130_fd_sc_hd__nand2_1
XFILLER_0_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _5058_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4821_ _3861_/A _4818_/Y _4819_/X _4760_/X _4820_/Y vssd1 vssd1 vccd1 vccd1 _4994_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_13_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5074_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4752_ _5008_/Q _4987_/Q _4750_/Y _4751_/X _4713_/X vssd1 vssd1 vccd1 vccd1 _5008_/D
+ sky130_fd_sc_hd__o221a_1
X_4683_ _4746_/A _5021_/Q vssd1 vssd1 vccd1 vccd1 _4683_/Y sky130_fd_sc_hd__nand2_1
X_3703_ _3703_/A _3703_/B vssd1 vssd1 vccd1 vccd1 _3703_/Y sky130_fd_sc_hd__nand2_1
X_3634_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3634_/X sky130_fd_sc_hd__clkbuf_2
X_3565_ _3566_/B _3566_/A vssd1 vssd1 vccd1 vccd1 _3567_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3496_ _3504_/B _3495_/Y _3568_/A vssd1 vssd1 vccd1 vccd1 _3496_/Y sky130_fd_sc_hd__a21oi_1
X_2516_ _2516_/A _4543_/A vssd1 vssd1 vccd1 vccd1 _2516_/Y sky130_fd_sc_hd__nand2_1
X_5235_ _5259_/CLK _5235_/D vssd1 vssd1 vccd1 vccd1 _5235_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5166_ _5168_/CLK _5166_/D vssd1 vssd1 vccd1 vccd1 _5166_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4117_ _4309_/A _4313_/A _4117_/C vssd1 vssd1 vccd1 vccd1 _4121_/C sky130_fd_sc_hd__nor3_1
X_5097_ _5281_/CLK _5097_/D vssd1 vssd1 vccd1 vccd1 _5097_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4048_ _4240_/A _4261_/A vssd1 vssd1 vccd1 vccd1 _4151_/B sky130_fd_sc_hd__nor2_1
XFILLER_12_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_74_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3350_ _3531_/A _3533_/A _3531_/B vssd1 vssd1 vccd1 vccd1 _3350_/X sky130_fd_sc_hd__o21ba_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ _5051_/CLK _5020_/D vssd1 vssd1 vccd1 vccd1 _5020_/Q sky130_fd_sc_hd__dfxtp_2
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _5203_/Q _3252_/X _3279_/Y _3280_/X _3259_/X vssd1 vssd1 vccd1 vccd1 _5203_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_2_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5090_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4804_ _4800_/A _4803_/Y _4501_/X vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__a21o_1
X_2996_ _5256_/Q _5160_/Q vssd1 vssd1 vccd1 vccd1 _3165_/B sky130_fd_sc_hd__and2_1
X_4735_ _4735_/A _4754_/B vssd1 vssd1 vccd1 vccd1 _4735_/Y sky130_fd_sc_hd__nand2_1
X_4666_ _4666_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4666_/Y sky130_fd_sc_hd__nor2_1
X_4597_ _5000_/Q _5032_/Q vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__nor2_1
X_3617_ _3820_/B _5106_/Q _3616_/X vssd1 vssd1 vccd1 vccd1 _3618_/B sky130_fd_sc_hd__o21a_1
X_3548_ _3468_/B _3548_/B _3548_/C vssd1 vssd1 vccd1 vccd1 _3548_/Y sky130_fd_sc_hd__nand3b_1
X_3479_ _3533_/A vssd1 vssd1 vccd1 vccd1 _3481_/A sky130_fd_sc_hd__inv_2
X_5218_ _5227_/CLK _5218_/D vssd1 vssd1 vccd1 vccd1 _5218_/Q sky130_fd_sc_hd__dfxtp_1
X_5149_ _5289_/CLK hold23/X vssd1 vssd1 vccd1 vccd1 _5149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2850_ _3598_/A vssd1 vssd1 vccd1 vccd1 _2850_/X sky130_fd_sc_hd__buf_4
X_2781_ _2869_/A _2869_/B _2734_/X vssd1 vssd1 vccd1 vccd1 _2781_/Y sky130_fd_sc_hd__a21oi_1
X_4520_ _4520_/A _4520_/B _4520_/C vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__and3_1
X_4451_ _4447_/A _4450_/Y _4407_/X vssd1 vssd1 vccd1 vccd1 _4451_/X sky130_fd_sc_hd__a21o_1
X_3402_ _3639_/B _3402_/B vssd1 vssd1 vccd1 vccd1 _3645_/B sky130_fd_sc_hd__nand2_1
XFILLER_7_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4382_ _4382_/A vssd1 vssd1 vccd1 vccd1 _4382_/Y sky130_fd_sc_hd__inv_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _5224_/Q vssd1 vssd1 vccd1 vccd1 _3761_/B sky130_fd_sc_hd__inv_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3264_ _5206_/Q _3261_/X _3247_/X _3263_/X vssd1 vssd1 vccd1 vccd1 _5206_/D sky130_fd_sc_hd__o211a_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5003_ _5272_/CLK _5003_/D vssd1 vssd1 vccd1 vccd1 _5003_/Q sky130_fd_sc_hd__dfxtp_1
X_3195_ _5219_/Q _3190_/X _3192_/X _3193_/Y _3194_/X vssd1 vssd1 vccd1 vccd1 _5219_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2979_ _2979_/A _2979_/B vssd1 vssd1 vccd1 vccd1 _2979_/Y sky130_fd_sc_hd__nand2_1
X_4718_ _5015_/Q _4987_/Q _4715_/X _4717_/X vssd1 vssd1 vccd1 vccd1 _5015_/D sky130_fd_sc_hd__o211a_1
X_4649_ _5016_/Q _5048_/Q vssd1 vssd1 vccd1 vccd1 _4651_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _4974_/Q hold20/A vssd1 vssd1 vccd1 vccd1 _3954_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2902_ _5241_/Q _2814_/X _2899_/X _2901_/Y _2822_/X vssd1 vssd1 vccd1 vccd1 _5241_/D
+ sky130_fd_sc_hd__o221a_1
X_3882_ _5088_/Q vssd1 vssd1 vccd1 vccd1 _3883_/A sky130_fd_sc_hd__inv_2
X_2833_ _2978_/A vssd1 vssd1 vccd1 vccd1 _3228_/B sky130_fd_sc_hd__buf_4
X_2764_ _2798_/A _2761_/Y _3568_/A vssd1 vssd1 vccd1 vccd1 _2764_/Y sky130_fd_sc_hd__a21oi_1
X_4503_ _4987_/Q _5029_/Q _4469_/X _4502_/X vssd1 vssd1 vccd1 vccd1 _5029_/D sky130_fd_sc_hd__o211a_1
X_2695_ _2695_/A vssd1 vssd1 vccd1 vccd1 _2695_/Y sky130_fd_sc_hd__inv_2
X_4434_ _4434_/A _4434_/B vssd1 vssd1 vccd1 vccd1 _4435_/B sky130_fd_sc_hd__nand2_1
X_4365_ _5086_/Q _5054_/Q vssd1 vssd1 vccd1 vccd1 _4368_/C sky130_fd_sc_hd__xnor2_1
X_3316_ _5197_/Q _3307_/X _3311_/Y _3313_/X _3315_/X vssd1 vssd1 vccd1 vccd1 _5197_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_86_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4296_ _4455_/B _4455_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _4296_/X sky130_fd_sc_hd__or3_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _3644_/A vssd1 vssd1 vccd1 vccd1 _3247_/X sky130_fd_sc_hd__clkbuf_2
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3178_ _3016_/X _3176_/Y _3147_/Y _2979_/B vssd1 vssd1 vccd1 vccd1 _3178_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_39_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2480_ _2836_/A vssd1 vssd1 vccd1 vccd1 _3528_/B sky130_fd_sc_hd__buf_4
X_4150_ _5064_/Q _4146_/A _4149_/Y vssd1 vssd1 vccd1 vccd1 _5064_/D sky130_fd_sc_hd__o21a_1
XFILLER_68_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3101_ _3101_/A _3101_/B vssd1 vssd1 vccd1 vccd1 _3243_/A sky130_fd_sc_hd__nor2_1
X_4081_ _4339_/A _4081_/B _4117_/C vssd1 vssd1 vccd1 vccd1 _4085_/C sky130_fd_sc_hd__nor3_1
XFILLER_83_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3032_ _3032_/A _3032_/B vssd1 vssd1 vccd1 vccd1 _3032_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4983_ _5045_/CLK _4983_/D vssd1 vssd1 vccd1 vccd1 _4983_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3934_ _4964_/Q _3934_/B vssd1 vssd1 vccd1 vccd1 _3987_/A sky130_fd_sc_hd__nor2_1
X_3865_ _3879_/A _4912_/A vssd1 vssd1 vccd1 vccd1 _3865_/Y sky130_fd_sc_hd__nand2_1
X_2816_ _2816_/A _2816_/B vssd1 vssd1 vccd1 vccd1 _2817_/A sky130_fd_sc_hd__nor2_1
X_3796_ _5115_/Q _3792_/X _3789_/X _3795_/Y vssd1 vssd1 vccd1 vccd1 _5115_/D sky130_fd_sc_hd__o211a_1
XFILLER_11_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2747_ _2815_/B _5019_/Q _2783_/A _2746_/Y vssd1 vssd1 vccd1 vccd1 _2806_/A sky130_fd_sc_hd__o22ai_2
X_2678_ _2678_/A vssd1 vssd1 vccd1 vccd1 _2771_/A sky130_fd_sc_hd__inv_2
X_4417_ _4987_/Q _5046_/Q _4414_/X _4416_/Y _4183_/X vssd1 vssd1 vccd1 vccd1 _5046_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4348_ _4406_/A _4406_/B _4347_/Y vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__o21bai_2
X_4279_ _4279_/A _4478_/C vssd1 vssd1 vccd1 vccd1 _4481_/B sky130_fd_sc_hd__nand2_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3650_ _3655_/A _3650_/B vssd1 vssd1 vccd1 vccd1 _3651_/B sky130_fd_sc_hd__or2_1
X_2601_ _2849_/A vssd1 vssd1 vccd1 vccd1 _2898_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3581_ _3581_/A _3581_/B vssd1 vssd1 vccd1 vccd1 _3590_/A sky130_fd_sc_hd__nor2_1
X_2532_ _5277_/Q _2525_/X _2526_/X _2531_/Y vssd1 vssd1 vccd1 vccd1 _5277_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5251_ _5251_/CLK _5251_/D vssd1 vssd1 vccd1 vccd1 _5251_/Q sky130_fd_sc_hd__dfxtp_1
X_4202_ _4202_/A _4538_/B vssd1 vssd1 vccd1 vccd1 _4383_/B sky130_fd_sc_hd__nor2_1
X_5182_ _5219_/CLK _5182_/D vssd1 vssd1 vccd1 vccd1 _5182_/Q sky130_fd_sc_hd__dfxtp_1
X_4133_ _4873_/A _4133_/B _4133_/C vssd1 vssd1 vccd1 vccd1 _5069_/D sky130_fd_sc_hd__nor3_1
X_4064_ _4064_/A vssd1 vssd1 vccd1 vccd1 _4065_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_68_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3015_ _3015_/A _3015_/B vssd1 vssd1 vccd1 vccd1 _3015_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4966_ _5064_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _4966_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_11_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3917_ _5072_/Q vssd1 vssd1 vccd1 vccd1 _4309_/A sky130_fd_sc_hd__inv_2
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4897_ _4901_/B vssd1 vssd1 vccd1 vccd1 _4902_/B sky130_fd_sc_hd__inv_2
XFILLER_32_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3848_ _4701_/A vssd1 vssd1 vccd1 vccd1 _4754_/B sky130_fd_sc_hd__clkbuf_4
X_3779_ _3792_/A vssd1 vssd1 vccd1 vccd1 _3779_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_78_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4820_ hold7/A _4820_/B vssd1 vssd1 vccd1 vccd1 _4820_/Y sky130_fd_sc_hd__nand2_1
X_4751_ _4750_/B _4750_/A _4711_/X vssd1 vssd1 vccd1 vccd1 _4751_/X sky130_fd_sc_hd__a21o_1
X_4682_ _4745_/A _4682_/B _4682_/C vssd1 vssd1 vccd1 vccd1 _4682_/X sky130_fd_sc_hd__or3_1
X_3702_ _5150_/Q _3698_/X _3695_/X _3701_/Y vssd1 vssd1 vccd1 vccd1 _5150_/D sky130_fd_sc_hd__o211a_1
X_3633_ _5168_/Q _3601_/X _3589_/X _3632_/X vssd1 vssd1 vccd1 vccd1 _5168_/D sky130_fd_sc_hd__o211a_1
X_3564_ _5181_/Q _3512_/X _3562_/Y _3563_/X _3518_/X vssd1 vssd1 vccd1 vccd1 _5181_/D
+ sky130_fd_sc_hd__o221a_1
X_2515_ _5014_/Q vssd1 vssd1 vccd1 vccd1 _4543_/A sky130_fd_sc_hd__inv_2
X_3495_ _3495_/A _3495_/B _3495_/C vssd1 vssd1 vccd1 vccd1 _3495_/Y sky130_fd_sc_hd__nor3_1
X_5234_ _5282_/CLK _5234_/D vssd1 vssd1 vccd1 vccd1 _5234_/Q sky130_fd_sc_hd__dfxtp_1
X_5165_ _5168_/CLK _5165_/D vssd1 vssd1 vccd1 vccd1 _5165_/Q sky130_fd_sc_hd__dfxtp_1
X_4116_ _4116_/A _4116_/B vssd1 vssd1 vccd1 vccd1 _5074_/D sky130_fd_sc_hd__nor2_1
XFILLER_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5096_ _5281_/CLK _5096_/D vssd1 vssd1 vccd1 vccd1 _5096_/Q sky130_fd_sc_hd__dfxtp_1
X_4047_ _5061_/Q vssd1 vssd1 vccd1 vccd1 _4261_/A sky130_fd_sc_hd__inv_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4949_ _4900_/X _4899_/B _4951_/S vssd1 vssd1 vccd1 vccd1 _4949_/X sky130_fd_sc_hd__mux2_1
XFILLER_58_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3280_ _3279_/B _3279_/A _3244_/X vssd1 vssd1 vccd1 vccd1 _3280_/X sky130_fd_sc_hd__a21o_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4803_ _4803_/A _4803_/B vssd1 vssd1 vccd1 vccd1 _4803_/Y sky130_fd_sc_hd__nand2_1
X_2995_ _3158_/A vssd1 vssd1 vccd1 vccd1 _2995_/Y sky130_fd_sc_hd__inv_2
X_4734_ _4734_/A _4734_/B vssd1 vssd1 vccd1 vccd1 _4734_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4665_ _4651_/B _4646_/A _4651_/A vssd1 vssd1 vccd1 vccd1 _4665_/X sky130_fd_sc_hd__o21ba_1
X_3616_ _3621_/B _3621_/A vssd1 vssd1 vccd1 vccd1 _3616_/X sky130_fd_sc_hd__or2_1
X_4596_ _4596_/A _4596_/B vssd1 vssd1 vccd1 vccd1 _4793_/A sky130_fd_sc_hd__nand2_1
X_3547_ _3548_/B _3548_/C _3468_/B vssd1 vssd1 vccd1 vccd1 _3547_/X sky130_fd_sc_hd__a21bo_1
XFILLER_0_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3478_ _3467_/B _3475_/Y _3477_/X _3473_/B vssd1 vssd1 vccd1 vccd1 _3538_/C sky130_fd_sc_hd__o22a_1
XFILLER_69_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5217_ _5230_/CLK _5217_/D vssd1 vssd1 vccd1 vccd1 _5217_/Q sky130_fd_sc_hd__dfxtp_1
X_5148_ _5289_/CLK _5148_/D vssd1 vssd1 vccd1 vccd1 _5148_/Q sky130_fd_sc_hd__dfxtp_1
X_5079_ _5080_/CLK _5079_/D vssd1 vssd1 vccd1 vccd1 _5079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_44_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2780_ _2780_/A vssd1 vssd1 vccd1 vccd1 _2869_/B sky130_fd_sc_hd__inv_2
X_4450_ _4450_/A _4450_/B vssd1 vssd1 vccd1 vccd1 _4450_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4381_/Y sky130_fd_sc_hd__inv_2
X_3401_ _3830_/B _5102_/Q vssd1 vssd1 vccd1 vccd1 _3402_/B sky130_fd_sc_hd__nand2_1
X_3332_ _5194_/Q _3307_/X _3330_/Y _3331_/Y _3315_/X vssd1 vssd1 vccd1 vccd1 _5194_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_85_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3263_ _3255_/X _3262_/Y _2930_/X vssd1 vssd1 vccd1 vccd1 _3263_/X sky130_fd_sc_hd__a21o_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _5272_/CLK _5002_/D vssd1 vssd1 vccd1 vccd1 _5002_/Q sky130_fd_sc_hd__dfxtp_1
X_3194_ _3259_/A vssd1 vssd1 vccd1 vccd1 _3194_/X sky130_fd_sc_hd__clkbuf_2
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2978_ _2978_/A vssd1 vssd1 vccd1 vccd1 _2979_/B sky130_fd_sc_hd__buf_2
X_4717_ _4709_/A _4716_/X _4501_/X vssd1 vssd1 vccd1 vccd1 _4717_/X sky130_fd_sc_hd__a21o_1
X_4648_ _4709_/B _4648_/B vssd1 vssd1 vccd1 vccd1 _4708_/A sky130_fd_sc_hd__nand2_1
X_4579_ _4579_/A _4579_/B vssd1 vssd1 vccd1 vccd1 _4826_/C sky130_fd_sc_hd__nand2_1
XFILLER_1_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3950_ _4954_/Q _4954_/D vssd1 vssd1 vccd1 vccd1 _3995_/C sky130_fd_sc_hd__xor2_2
XFILLER_63_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2901_ _2901_/A _2901_/B vssd1 vssd1 vccd1 vccd1 _2901_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3881_ _3881_/A vssd1 vssd1 vccd1 vccd1 _4479_/A sky130_fd_sc_hd__clkbuf_4
X_2832_ _5252_/Q vssd1 vssd1 vccd1 vccd1 _3686_/B sky130_fd_sc_hd__inv_2
X_2763_ _3577_/A vssd1 vssd1 vccd1 vccd1 _3568_/A sky130_fd_sc_hd__buf_4
X_4502_ _4497_/A _4500_/Y _4501_/X vssd1 vssd1 vccd1 vccd1 _4502_/X sky130_fd_sc_hd__a21o_1
X_2694_ _2654_/Y _2685_/Y _2693_/Y vssd1 vssd1 vccd1 vccd1 _2908_/A sky130_fd_sc_hd__o21bai_1
X_4433_ _4440_/B _4440_/A vssd1 vssd1 vccd1 vccd1 _4434_/A sky130_fd_sc_hd__nand2_1
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4364_ _4373_/A _4360_/Y _4373_/B vssd1 vssd1 vccd1 vccd1 _4364_/Y sky130_fd_sc_hd__a21oi_1
X_4295_ _4457_/B _4295_/B vssd1 vssd1 vccd1 vccd1 _4460_/B sky130_fd_sc_hd__nand2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _4183_/A vssd1 vssd1 vccd1 vccd1 _3315_/X sky130_fd_sc_hd__clkbuf_2
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3246_ _5209_/Q _3190_/X _3243_/Y _3245_/X _3194_/X vssd1 vssd1 vccd1 vccd1 _5209_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3177_ _3016_/X _3147_/Y _3176_/Y vssd1 vssd1 vccd1 vccd1 _3177_/X sky130_fd_sc_hd__o21a_1
XFILLER_39_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_82_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3100_ _3100_/A vssd1 vssd1 vccd1 vccd1 _3101_/B sky130_fd_sc_hd__inv_2
X_4080_ _4080_/A vssd1 vssd1 vccd1 vccd1 _4081_/B sky130_fd_sc_hd__inv_2
XFILLER_83_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3031_ _3111_/A _3110_/A _3111_/B vssd1 vssd1 vccd1 vccd1 _3031_/X sky130_fd_sc_hd__o21ba_1
XFILLER_36_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4982_ _5045_/CLK _4982_/D vssd1 vssd1 vccd1 vccd1 _4982_/Q sky130_fd_sc_hd__dfxtp_1
X_3933_ _3934_/B _4964_/Q vssd1 vssd1 vccd1 vccd1 _3987_/B sky130_fd_sc_hd__and2_1
X_3864_ _5093_/Q vssd1 vssd1 vccd1 vccd1 _4912_/A sky130_fd_sc_hd__inv_2
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2815_ _5019_/Q _2815_/B vssd1 vssd1 vccd1 vccd1 _2816_/B sky130_fd_sc_hd__nor2_1
X_3795_ _3797_/A _3795_/B vssd1 vssd1 vccd1 vccd1 _3795_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2746_ _2824_/A _2824_/B _2745_/Y vssd1 vssd1 vccd1 vccd1 _2746_/Y sky130_fd_sc_hd__a21oi_1
X_2677_ _2656_/Y _2953_/A _2767_/A _2676_/Y vssd1 vssd1 vccd1 vccd1 _2677_/Y sky130_fd_sc_hd__o211ai_1
X_4416_ _4416_/A _4987_/Q vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__nand2_1
X_4347_ _4347_/A _4347_/B vssd1 vssd1 vccd1 vccd1 _4347_/Y sky130_fd_sc_hd__nand2_1
X_4278_ _4278_/A _4603_/B vssd1 vssd1 vccd1 vccd1 _4279_/A sky130_fd_sc_hd__nand2_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _3229_/A _3229_/B vssd1 vssd1 vccd1 vccd1 _3230_/C sky130_fd_sc_hd__nand2_1
XFILLER_36_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3580_ _3634_/A vssd1 vssd1 vccd1 vccd1 _3580_/X sky130_fd_sc_hd__clkbuf_2
X_2600_ _2600_/A vssd1 vssd1 vccd1 vccd1 _2849_/A sky130_fd_sc_hd__inv_2
X_2531_ _2534_/A _4623_/A vssd1 vssd1 vccd1 vccd1 _2531_/Y sky130_fd_sc_hd__nand2_1
X_5250_ _5289_/CLK _5250_/D vssd1 vssd1 vccd1 vccd1 _5250_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4201_ _5051_/Q vssd1 vssd1 vccd1 vccd1 _4538_/B sky130_fd_sc_hd__inv_2
XFILLER_5_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5181_ _5181_/CLK _5181_/D vssd1 vssd1 vccd1 vccd1 _5181_/Q sky130_fd_sc_hd__dfxtp_1
X_4132_ _4125_/A _4074_/X _4075_/X _4134_/C _5069_/Q vssd1 vssd1 vccd1 vccd1 _4133_/B
+ sky130_fd_sc_hd__a41oi_1
XFILLER_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4063_ _4359_/A _4202_/A _4063_/C vssd1 vssd1 vccd1 vccd1 _4065_/B sky130_fd_sc_hd__or3_1
XFILLER_83_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3014_ _3014_/A vssd1 vssd1 vccd1 vccd1 _3186_/A sky130_fd_sc_hd__inv_2
XFILLER_36_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4965_ _5064_/CLK _4965_/D vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__dfxtp_1
X_3916_ _5073_/Q vssd1 vssd1 vccd1 vccd1 _4299_/A sky130_fd_sc_hd__inv_2
X_4896_ _5090_/Q _5089_/Q _5088_/Q vssd1 vssd1 vccd1 vccd1 _4901_/B sky130_fd_sc_hd__and3_1
XFILLER_32_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3847_ _4395_/A vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3778_ _5122_/Q _3766_/X _3776_/X _3777_/Y vssd1 vssd1 vccd1 vccd1 _5122_/D sky130_fd_sc_hd__o211a_1
X_2729_ _2729_/A _2729_/B vssd1 vssd1 vccd1 vccd1 _2862_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4750_ _4750_/A _4750_/B vssd1 vssd1 vccd1 vccd1 _4750_/Y sky130_fd_sc_hd__nor2_1
X_4681_ _4681_/A _4681_/B _4681_/C vssd1 vssd1 vccd1 vccd1 _4682_/C sky130_fd_sc_hd__and3_1
X_3701_ _3703_/A _3701_/B vssd1 vssd1 vccd1 vccd1 _3701_/Y sky130_fd_sc_hd__nand2_1
X_3632_ _3630_/X _3631_/Y _2603_/A vssd1 vssd1 vccd1 vccd1 _3632_/X sky130_fd_sc_hd__a21o_1
X_3563_ _3562_/B _3562_/A _3312_/X vssd1 vssd1 vccd1 vccd1 _3563_/X sky130_fd_sc_hd__a21o_1
X_3494_ _3335_/Y _3504_/B _3495_/B _3495_/C vssd1 vssd1 vccd1 vccd1 _3494_/Y sky130_fd_sc_hd__o2bb2ai_1
X_2514_ _5282_/Q _2506_/X _2507_/X _2513_/Y vssd1 vssd1 vccd1 vccd1 _5282_/D sky130_fd_sc_hd__o211a_1
X_5233_ _5259_/CLK _5233_/D vssd1 vssd1 vccd1 vccd1 _5233_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5164_ _5168_/CLK _5164_/D vssd1 vssd1 vccd1 vccd1 _5164_/Q sky130_fd_sc_hd__dfxtp_1
X_4115_ _4115_/A _4115_/B vssd1 vssd1 vccd1 vccd1 _4116_/B sky130_fd_sc_hd__nand2_1
XFILLER_29_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5095_ _5281_/CLK _5095_/D vssd1 vssd1 vccd1 vccd1 _5095_/Q sky130_fd_sc_hd__dfxtp_1
X_4046_ _5062_/Q vssd1 vssd1 vccd1 vccd1 _4240_/A sky130_fd_sc_hd__inv_2
XFILLER_71_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4948_ _4905_/X _4904_/B _4951_/S vssd1 vssd1 vccd1 vccd1 _4948_/X sky130_fd_sc_hd__mux2_1
X_4879_ _3861_/B _4983_/Q _3883_/A _4977_/Q _4878_/X vssd1 vssd1 vccd1 vccd1 _4880_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_79_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2994_ _5160_/Q _3674_/B vssd1 vssd1 vccd1 vccd1 _3158_/A sky130_fd_sc_hd__nor2_1
X_4802_ _4516_/X _4799_/Y _4800_/X _4760_/X _4801_/Y vssd1 vssd1 vccd1 vccd1 _4998_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4733_ _5012_/Q _4987_/Q _4731_/Y _4732_/X _4713_/X vssd1 vssd1 vccd1 vccd1 _5012_/D
+ sky130_fd_sc_hd__o221a_1
X_4664_ _4716_/A _4716_/B _4663_/Y vssd1 vssd1 vccd1 vccd1 _4692_/A sky130_fd_sc_hd__o21bai_2
X_3615_ _3615_/A _3615_/B vssd1 vssd1 vccd1 vccd1 _3621_/A sky130_fd_sc_hd__and2_1
X_4595_ _4999_/Q _5031_/Q vssd1 vssd1 vccd1 vccd1 _4596_/B sky130_fd_sc_hd__nand2_1
X_3546_ _3551_/B _3551_/A vssd1 vssd1 vccd1 vccd1 _3548_/B sky130_fd_sc_hd__or2_1
X_5216_ _5219_/CLK _5216_/D vssd1 vssd1 vccd1 vccd1 _5216_/Q sky130_fd_sc_hd__dfxtp_1
X_3477_ _3476_/Y _3458_/A _3472_/B vssd1 vssd1 vccd1 vccd1 _3477_/X sky130_fd_sc_hd__a21o_1
XFILLER_69_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5147_ _5254_/CLK _5147_/D vssd1 vssd1 vccd1 vccd1 _5147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5078_ _5080_/CLK _5078_/D vssd1 vssd1 vccd1 vccd1 _5078_/Q sky130_fd_sc_hd__dfxtp_1
X_4029_ _5056_/Q _4025_/X _4192_/B _4177_/A vssd1 vssd1 vccd1 vccd1 _4030_/C sky130_fd_sc_hd__o211ai_1
XFILLER_71_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4380_ _4987_/Q _5052_/Q _4377_/X _4379_/Y _4183_/X vssd1 vssd1 vccd1 vccd1 _5052_/D
+ sky130_fd_sc_hd__o221a_1
X_3400_ _3400_/A vssd1 vssd1 vccd1 vccd1 _3649_/A sky130_fd_sc_hd__inv_2
X_3331_ _3668_/A _3331_/B vssd1 vssd1 vccd1 vccd1 _3331_/Y sky130_fd_sc_hd__nand2_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _3262_/A _3262_/B vssd1 vssd1 vccd1 vccd1 _3262_/Y sky130_fd_sc_hd__nand2_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _3145_/B _3005_/A _3197_/B _2979_/B vssd1 vssd1 vccd1 vccd1 _3193_/Y sky130_fd_sc_hd__o31ai_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _5288_/CLK _5001_/D vssd1 vssd1 vccd1 vccd1 _5001_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_78_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2977_ _2977_/A _2977_/B _2977_/C vssd1 vssd1 vccd1 vccd1 _2979_/A sky130_fd_sc_hd__or3_1
X_4716_ _4716_/A _4716_/B _4708_/A vssd1 vssd1 vccd1 vccd1 _4716_/X sky130_fd_sc_hd__or3b_1
X_4647_ hold15/A _4647_/B vssd1 vssd1 vccd1 vccd1 _4648_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4578_ _5025_/Q vssd1 vssd1 vccd1 vccd1 _4579_/B sky130_fd_sc_hd__inv_2
X_3529_ _3568_/A _5188_/Q vssd1 vssd1 vccd1 vccd1 _3529_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_75_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2900_ _2900_/A _2900_/B vssd1 vssd1 vccd1 vccd1 _2901_/B sky130_fd_sc_hd__and2_1
XFILLER_45_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3880_ _3867_/X _4950_/X _3868_/X _3879_/Y vssd1 vssd1 vccd1 vccd1 _5089_/D sky130_fd_sc_hd__o211a_1
XFILLER_43_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2831_ _2803_/X _2827_/Y _2828_/X _2808_/X _2830_/Y vssd1 vssd1 vccd1 vccd1 _5253_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2762_ _2849_/A vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__clkbuf_2
X_4501_ _4501_/A vssd1 vssd1 vccd1 vccd1 _4501_/X sky130_fd_sc_hd__clkbuf_4
X_4432_ _4316_/B _4450_/A _4318_/Y vssd1 vssd1 vccd1 vccd1 _4440_/B sky130_fd_sc_hd__o21ai_1
XANTENNA_0 _4849_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2693_ _2929_/A _2926_/A vssd1 vssd1 vccd1 vccd1 _2693_/Y sky130_fd_sc_hd__nand2_1
X_4363_ _4363_/A _4363_/B vssd1 vssd1 vccd1 vccd1 _4373_/B sky130_fd_sc_hd__nor2_1
X_4294_ _4294_/A _4556_/B vssd1 vssd1 vccd1 vccd1 _4295_/B sky130_fd_sc_hd__nand2_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _4103_/A vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__clkbuf_8
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _3243_/B _3243_/A _3244_/X vssd1 vssd1 vccd1 vccd1 _3245_/X sky130_fd_sc_hd__a21o_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3176_ _3176_/A vssd1 vssd1 vccd1 vccd1 _3176_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3030_ _3709_/B _5147_/Q vssd1 vssd1 vccd1 vccd1 _3111_/B sky130_fd_sc_hd__and2_1
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _5281_/CLK _4981_/D vssd1 vssd1 vccd1 vccd1 _4981_/Q sky130_fd_sc_hd__dfxtp_1
X_3932_ hold8/A vssd1 vssd1 vccd1 vccd1 _3934_/B sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_43_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5168_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3863_ _3881_/A vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__clkbuf_2
X_2814_ _3230_/B vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__clkbuf_2
X_3794_ _5116_/Q _3792_/X _3789_/X _3793_/Y vssd1 vssd1 vccd1 vccd1 _5116_/D sky130_fd_sc_hd__o211a_1
X_2745_ _2745_/A _2825_/B vssd1 vssd1 vccd1 vccd1 _2745_/Y sky130_fd_sc_hd__nand2_1
X_2676_ _2768_/A _2945_/A vssd1 vssd1 vccd1 vccd1 _2676_/Y sky130_fd_sc_hd__nor2_1
X_4415_ _4415_/A _4415_/B _4415_/C vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__or3_1
X_4346_ _4396_/B _4353_/C vssd1 vssd1 vccd1 vccd1 _4347_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4277_ _5033_/Q vssd1 vssd1 vccd1 vccd1 _4603_/B sky130_fd_sc_hd__inv_2
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3228_ _3793_/B _3228_/B vssd1 vssd1 vccd1 vccd1 _3228_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3159_ _3167_/B _3158_/Y _3568_/A vssd1 vssd1 vccd1 vccd1 _3159_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_34_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5213_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_2_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_25_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _5288_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_9_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2530_ _5010_/Q vssd1 vssd1 vccd1 vccd1 _4623_/A sky130_fd_sc_hd__inv_2
XFILLER_5_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4200_ _4362_/B _4537_/B vssd1 vssd1 vccd1 vccd1 _4200_/Y sky130_fd_sc_hd__nor2_1
XFILLER_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5180_ _5181_/CLK _5180_/D vssd1 vssd1 vccd1 vccd1 _5180_/Q sky130_fd_sc_hd__dfxtp_1
X_4131_ _5070_/Q _4133_/C _4130_/Y vssd1 vssd1 vccd1 vccd1 _5070_/D sky130_fd_sc_hd__o21a_1
XFILLER_3_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4062_ _5083_/Q vssd1 vssd1 vccd1 vccd1 _4202_/A sky130_fd_sc_hd__inv_2
XFILLER_83_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3013_ _3015_/B _3013_/B vssd1 vssd1 vccd1 vccd1 _3014_/A sky130_fd_sc_hd__nand2_1
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4964_ _4964_/CLK hold8/X vssd1 vssd1 vccd1 vccd1 _4964_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_16_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _5272_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_51_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3915_ _5074_/Q vssd1 vssd1 vccd1 vccd1 _4304_/A sky130_fd_sc_hd__inv_2
X_4895_ _4895_/A vssd1 vssd1 vccd1 vccd1 _4895_/X sky130_fd_sc_hd__clkbuf_1
X_3846_ _5097_/Q vssd1 vssd1 vccd1 vccd1 _3897_/B sky130_fd_sc_hd__inv_2
X_3777_ _3784_/A _3777_/B vssd1 vssd1 vccd1 vccd1 _3777_/Y sky130_fd_sc_hd__nand2_1
X_2728_ _4726_/B _5280_/Q vssd1 vssd1 vccd1 vccd1 _2729_/B sky130_fd_sc_hd__nand2_1
X_2659_ _5258_/Q _2990_/B _4992_/Q _2985_/B vssd1 vssd1 vccd1 vccd1 _2975_/A sky130_fd_sc_hd__o2bb2ai_1
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4329_ _4329_/A _4402_/B vssd1 vssd1 vccd1 vccd1 _4335_/A sky130_fd_sc_hd__nand2_1
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3700_ _5151_/Q _3698_/X _3695_/X _3699_/Y vssd1 vssd1 vccd1 vccd1 _5151_/D sky130_fd_sc_hd__o211a_1
XFILLER_53_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4680_ _4873_/A _4680_/B _4680_/C vssd1 vssd1 vccd1 vccd1 _5022_/D sky130_fd_sc_hd__nor3_1
X_3631_ _3631_/A _3631_/B vssd1 vssd1 vccd1 vccd1 _3631_/Y sky130_fd_sc_hd__nand2_1
X_3562_ _3562_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3562_/Y sky130_fd_sc_hd__nor2_1
X_2513_ _2516_/A hold15/X vssd1 vssd1 vccd1 vccd1 _2513_/Y sky130_fd_sc_hd__nand2_1
X_3493_ _3758_/B _5129_/Q vssd1 vssd1 vccd1 vccd1 _3495_/C sky130_fd_sc_hd__and2_1
X_5232_ _5254_/CLK _5232_/D vssd1 vssd1 vccd1 vccd1 _5232_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_5_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5287_/CLK sky130_fd_sc_hd__clkbuf_16
X_5163_ _5168_/CLK _5163_/D vssd1 vssd1 vccd1 vccd1 _5163_/Q sky130_fd_sc_hd__dfxtp_1
X_4114_ _4130_/B _4113_/X _5074_/Q vssd1 vssd1 vccd1 vccd1 _4116_/A sky130_fd_sc_hd__a21oi_1
XFILLER_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5094_ _5282_/CLK _5094_/D vssd1 vssd1 vccd1 vccd1 _5094_/Q sky130_fd_sc_hd__dfxtp_1
X_4045_ _4125_/A _5070_/Q _5069_/Q vssd1 vssd1 vccd1 vccd1 _4049_/B sky130_fd_sc_hd__and3_1
XFILLER_37_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4947_ _4911_/X _4910_/B _4951_/S vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__mux2_1
X_4878_ _5097_/Q _3901_/Y _5095_/Q _3899_/Y vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__o22a_1
X_3829_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3829_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_20_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_90_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_65_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4801_ _4801_/A _4820_/B vssd1 vssd1 vccd1 vccd1 _4801_/Y sky130_fd_sc_hd__nand2_1
X_2993_ _5256_/Q vssd1 vssd1 vccd1 vccd1 _3674_/B sky130_fd_sc_hd__inv_2
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4732_ _4731_/B _4731_/A _4711_/X vssd1 vssd1 vccd1 vccd1 _4732_/X sky130_fd_sc_hd__a21o_1
X_4663_ _4663_/A _4663_/B vssd1 vssd1 vccd1 vccd1 _4663_/Y sky130_fd_sc_hd__nand2_1
X_3614_ _3614_/A vssd1 vssd1 vccd1 vccd1 _3618_/A sky130_fd_sc_hd__inv_2
X_4594_ _4794_/A _4594_/B vssd1 vssd1 vccd1 vccd1 _4596_/A sky130_fd_sc_hd__nand2_1
X_3545_ _3544_/Y _3476_/Y _3458_/A _3472_/B vssd1 vssd1 vccd1 vccd1 _3551_/A sky130_fd_sc_hd__a31o_1
X_3476_ _3476_/A vssd1 vssd1 vccd1 vccd1 _3476_/Y sky130_fd_sc_hd__inv_2
X_5215_ _5215_/CLK _5215_/D vssd1 vssd1 vccd1 vccd1 _5215_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5146_ _5254_/CLK _5146_/D vssd1 vssd1 vccd1 vccd1 _5146_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5077_ _5080_/CLK _5077_/D vssd1 vssd1 vccd1 vccd1 _5077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4028_ _4191_/A _4191_/B _5055_/Q vssd1 vssd1 vccd1 vccd1 _4177_/A sky130_fd_sc_hd__a21boi_1
XFILLER_44_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3330_ _5130_/Q _3756_/B vssd1 vssd1 vccd1 vccd1 _3330_/Y sky130_fd_sc_hd__nor2_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _5265_/CLK _5000_/D vssd1 vssd1 vccd1 vccd1 _5000_/Q sky130_fd_sc_hd__dfxtp_1
X_3261_ _3601_/A vssd1 vssd1 vccd1 vccd1 _3261_/X sky130_fd_sc_hd__clkbuf_2
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3192_ _3005_/A _3197_/B _3145_/B vssd1 vssd1 vccd1 vccd1 _3192_/X sky130_fd_sc_hd__o21a_1
XFILLER_38_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2976_ _2977_/A _2977_/B _2977_/C vssd1 vssd1 vccd1 vccd1 _2976_/X sky130_fd_sc_hd__o21a_1
X_4715_ _4784_/A vssd1 vssd1 vccd1 vccd1 _4715_/X sky130_fd_sc_hd__clkbuf_2
X_4646_ _4646_/A vssd1 vssd1 vccd1 vccd1 _4709_/B sky130_fd_sc_hd__inv_2
X_4577_ _4992_/Q _5024_/Q vssd1 vssd1 vccd1 vccd1 _4823_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3528_ _3528_/A _3528_/B _3528_/C vssd1 vssd1 vccd1 vccd1 _3528_/Y sky130_fd_sc_hd__nand3_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3459_ _5216_/Q vssd1 vssd1 vccd1 vccd1 _3782_/B sky130_fd_sc_hd__inv_2
X_5129_ _5227_/CLK _5129_/D vssd1 vssd1 vccd1 vccd1 _5129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2830_ _3238_/A hold17/A vssd1 vssd1 vccd1 vccd1 _2830_/Y sky130_fd_sc_hd__nand2_1
X_2761_ _2761_/A _2761_/B _2761_/C vssd1 vssd1 vccd1 vccd1 _2761_/Y sky130_fd_sc_hd__nor3_1
X_4500_ _4500_/A _4500_/B vssd1 vssd1 vccd1 vccd1 _4500_/Y sky130_fd_sc_hd__nand2_1
X_2692_ _2695_/A _2692_/B vssd1 vssd1 vccd1 vccd1 _2926_/A sky130_fd_sc_hd__nor2_1
X_4431_ _4431_/A _4431_/B vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__nor2_1
XANTENNA_1 _3861_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4362_ _5053_/Q _4362_/B vssd1 vssd1 vccd1 vccd1 _4363_/B sky130_fd_sc_hd__nor2_1
X_4293_ _4289_/A _4285_/B _4289_/B vssd1 vssd1 vccd1 vccd1 _4453_/B sky130_fd_sc_hd__o21ba_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _3311_/B _3311_/A _3312_/X vssd1 vssd1 vccd1 vccd1 _3313_/X sky130_fd_sc_hd__a21o_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _3598_/A vssd1 vssd1 vccd1 vccd1 _3244_/X sky130_fd_sc_hd__clkbuf_2
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3175_ _3175_/A _3175_/B vssd1 vssd1 vccd1 vccd1 _3176_/A sky130_fd_sc_hd__nor2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2959_ _3238_/A _3742_/B vssd1 vssd1 vccd1 vccd1 _2959_/Y sky130_fd_sc_hd__nand2_1
XFILLER_41_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4629_ _4629_/A _4631_/B vssd1 vssd1 vccd1 vccd1 _4630_/A sky130_fd_sc_hd__nor2_1
XFILLER_1_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _5090_/CLK _4980_/D vssd1 vssd1 vccd1 vccd1 _4980_/Q sky130_fd_sc_hd__dfxtp_1
X_3931_ _3931_/A _5086_/Q vssd1 vssd1 vccd1 vccd1 _4052_/B sky130_fd_sc_hd__nand2_1
X_3862_ _3844_/X _4945_/X _3845_/X _3861_/Y vssd1 vssd1 vccd1 vccd1 _5094_/D sky130_fd_sc_hd__o211a_1
X_2813_ _3718_/A vssd1 vssd1 vccd1 vccd1 _3230_/B sky130_fd_sc_hd__buf_2
X_3793_ _3797_/A _3793_/B vssd1 vssd1 vccd1 vccd1 _3793_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2744_ _2844_/A _2843_/B _2841_/C vssd1 vssd1 vccd1 vccd1 _2825_/B sky130_fd_sc_hd__and3_1
X_2675_ _2678_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _2945_/A sky130_fd_sc_hd__nand2_1
X_4414_ _4415_/B _4415_/C _4415_/A vssd1 vssd1 vccd1 vccd1 _4414_/X sky130_fd_sc_hd__o21a_1
X_4345_ _4345_/A vssd1 vssd1 vccd1 vccd1 _4353_/C sky130_fd_sc_hd__inv_2
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4276_ _4273_/A _4486_/B _4273_/B vssd1 vssd1 vccd1 vccd1 _4474_/B sky130_fd_sc_hd__o21ba_1
X_3227_ _5212_/Q vssd1 vssd1 vccd1 vccd1 _3793_/B sky130_fd_sc_hd__inv_2
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3158_ _3158_/A _3158_/B _3158_/C vssd1 vssd1 vccd1 vccd1 _3158_/Y sky130_fd_sc_hd__nor3_1
XFILLER_82_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3089_ _3265_/A _3265_/B _3088_/X vssd1 vssd1 vccd1 vccd1 _3254_/A sky130_fd_sc_hd__o21bai_1
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_73_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4130_ _4873_/A _4130_/B vssd1 vssd1 vccd1 vccd1 _4130_/Y sky130_fd_sc_hd__nor2_1
X_4061_ _5084_/Q vssd1 vssd1 vccd1 vccd1 _4359_/A sky130_fd_sc_hd__inv_2
XFILLER_68_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3012_ _3686_/B _5156_/Q vssd1 vssd1 vccd1 vccd1 _3013_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4963_ _5064_/CLK _4963_/D vssd1 vssd1 vccd1 vccd1 hold8/A sky130_fd_sc_hd__dfxtp_1
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3914_ _4343_/A _4339_/A _4332_/A _4327_/A vssd1 vssd1 vccd1 vccd1 _4063_/C sky130_fd_sc_hd__or4_1
XFILLER_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4894_ _4915_/A _4894_/B vssd1 vssd1 vccd1 vccd1 _4895_/A sky130_fd_sc_hd__and2_1
XFILLER_32_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3845_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3845_/X sky130_fd_sc_hd__clkbuf_2
X_3776_ _3802_/A vssd1 vssd1 vccd1 vccd1 _3776_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2727_ _5280_/Q _4726_/B vssd1 vssd1 vccd1 vccd1 _2729_/A sky130_fd_sc_hd__or2_1
X_2658_ _5260_/Q _4579_/A vssd1 vssd1 vccd1 vccd1 _2977_/A sky130_fd_sc_hd__nor2_1
X_2589_ _5263_/Q _2584_/X _2585_/X _2588_/Y vssd1 vssd1 vccd1 vccd1 _5263_/D sky130_fd_sc_hd__o211a_1
X_4328_ _5079_/Q _5047_/Q vssd1 vssd1 vccd1 vccd1 _4402_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4259_ _4259_/A _4259_/B vssd1 vssd1 vccd1 vccd1 _4494_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3630_ _3631_/B _3631_/A vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__or2_1
X_3561_ _3566_/B _3566_/A _3370_/B vssd1 vssd1 vccd1 vccd1 _3562_/B sky130_fd_sc_hd__o21a_1
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2512_ _4645_/A vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__clkbuf_2
X_3492_ _5129_/Q _3758_/B vssd1 vssd1 vccd1 vccd1 _3495_/B sky130_fd_sc_hd__nor2_1
X_5231_ _5282_/CLK _5231_/D vssd1 vssd1 vccd1 vccd1 _5231_/Q sky130_fd_sc_hd__dfxtp_1
X_5162_ _5168_/CLK _5162_/D vssd1 vssd1 vccd1 vccd1 _5162_/Q sky130_fd_sc_hd__dfxtp_1
X_4113_ _5073_/Q _5072_/Q _5071_/Q vssd1 vssd1 vccd1 vccd1 _4113_/X sky130_fd_sc_hd__and3_1
X_5093_ _5282_/CLK _5093_/D vssd1 vssd1 vccd1 vccd1 _5093_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_68_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4044_ _4288_/A _4283_/A vssd1 vssd1 vccd1 vccd1 _4125_/A sky130_fd_sc_hd__nor2_1
XFILLER_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4946_ _4916_/X _4915_/B _4951_/S vssd1 vssd1 vccd1 vccd1 _4946_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4877_ _5092_/Q _3902_/Y _5091_/Q _3895_/Y _4876_/X vssd1 vssd1 vccd1 vccd1 _4880_/B
+ sky130_fd_sc_hd__o221a_1
X_3828_ _5103_/Q _3819_/X _3816_/X _3827_/Y vssd1 vssd1 vccd1 vccd1 _5103_/D sky130_fd_sc_hd__o211a_1
X_3759_ _5129_/Q _3753_/X _3750_/X _3758_/Y vssd1 vssd1 vccd1 vccd1 _5129_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4800_ _4800_/A _4800_/B _4800_/C vssd1 vssd1 vccd1 vccd1 _4800_/X sky130_fd_sc_hd__and3_1
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2992_ _5226_/Q _2972_/X _2990_/Y _2991_/Y _2980_/X vssd1 vssd1 vccd1 vccd1 _5226_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_9_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4731_ _4731_/A _4731_/B vssd1 vssd1 vccd1 vccd1 _4731_/Y sky130_fd_sc_hd__nor2_1
X_4662_ _4704_/B _4662_/B vssd1 vssd1 vccd1 vccd1 _4663_/B sky130_fd_sc_hd__nor2_1
X_3613_ _5172_/Q _3601_/X _3589_/X _3612_/X vssd1 vssd1 vccd1 vccd1 _5172_/D sky130_fd_sc_hd__o211a_1
X_4593_ _4797_/A _4797_/B _4592_/Y vssd1 vssd1 vccd1 vccd1 _4788_/B sky130_fd_sc_hd__a21oi_1
X_3544_ _3557_/B _3557_/A vssd1 vssd1 vccd1 vccd1 _3544_/Y sky130_fd_sc_hd__nand2_1
X_3475_ _3475_/A _3475_/B vssd1 vssd1 vccd1 vccd1 _3475_/Y sky130_fd_sc_hd__nor2_1
X_5214_ _5215_/CLK _5214_/D vssd1 vssd1 vccd1 vccd1 _5214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5145_ _5254_/CLK _5145_/D vssd1 vssd1 vccd1 vccd1 _5145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5076_ _5076_/CLK _5076_/D vssd1 vssd1 vccd1 vccd1 _5076_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_84_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4027_ _4027_/A vssd1 vssd1 vccd1 vccd1 _4191_/B sky130_fd_sc_hd__inv_2
XFILLER_52_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4929_ _4929_/A vssd1 vssd1 vccd1 vccd1 _4929_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _5207_/Q _3252_/X _3257_/Y _3258_/X _3259_/X vssd1 vssd1 vccd1 vccd1 _5207_/D
+ sky130_fd_sc_hd__o221a_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3191_ _3196_/B _3191_/B vssd1 vssd1 vccd1 vccd1 _3197_/B sky130_fd_sc_hd__nor2_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4714_ _5016_/Q _4987_/Q _4710_/Y _4712_/X _4713_/X vssd1 vssd1 vccd1 vccd1 _5016_/D
+ sky130_fd_sc_hd__o221a_1
X_2975_ _2975_/A _2986_/B vssd1 vssd1 vccd1 vccd1 _2977_/C sky130_fd_sc_hd__nand2_1
X_4645_ _4645_/A _4647_/B vssd1 vssd1 vccd1 vccd1 _4646_/A sky130_fd_sc_hd__nor2_1
X_4576_ _4576_/A _4810_/C vssd1 vssd1 vccd1 vccd1 _4813_/A sky130_fd_sc_hd__and2_1
X_3527_ _3527_/A _3527_/B vssd1 vssd1 vccd1 vccd1 _3528_/C sky130_fd_sc_hd__nand2_1
X_3458_ _3458_/A _3458_/B vssd1 vssd1 vccd1 vccd1 _3543_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3389_ _5101_/Q vssd1 vssd1 vccd1 vccd1 _3389_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5128_ _5227_/CLK _5128_/D vssd1 vssd1 vccd1 vccd1 _5128_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _5063_/CLK _5059_/D vssd1 vssd1 vccd1 vccd1 _5059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_52_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_71_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2760_ _4940_/B _5289_/Q vssd1 vssd1 vccd1 vccd1 _2761_/C sky130_fd_sc_hd__and2_1
X_2691_ _4782_/A _5269_/Q vssd1 vssd1 vccd1 vccd1 _2692_/B sky130_fd_sc_hd__and2_1
XANTENNA_2 _4760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _4430_/A vssd1 vssd1 vccd1 vccd1 _4435_/A sky130_fd_sc_hd__inv_2
X_4361_ _5085_/Q _4537_/B vssd1 vssd1 vccd1 vccd1 _4363_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4292_ _4463_/A _4463_/B _4291_/Y vssd1 vssd1 vccd1 vccd1 _4453_/A sky130_fd_sc_hd__o21ai_1
X_3312_ _3598_/A vssd1 vssd1 vccd1 vccd1 _3312_/X sky130_fd_sc_hd__buf_2
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _3243_/A _3243_/B vssd1 vssd1 vccd1 vccd1 _3243_/Y sky130_fd_sc_hd__nor2_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3174_ _5254_/Q _3174_/B vssd1 vssd1 vccd1 vccd1 _3175_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2958_ _5231_/Q vssd1 vssd1 vccd1 vccd1 _3742_/B sky130_fd_sc_hd__clkinv_2
X_2889_ _2889_/A _2889_/B vssd1 vssd1 vccd1 vccd1 _2890_/B sky130_fd_sc_hd__nand2_1
X_4628_ _4628_/A _4628_/B vssd1 vssd1 vccd1 vccd1 _4748_/B sky130_fd_sc_hd__nor2_1
XFILLER_1_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4559_ _4761_/A _4559_/B vssd1 vssd1 vccd1 vccd1 _4617_/B sky130_fd_sc_hd__nor2_1
XFILLER_77_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput50 _5166_/Q vssd1 vssd1 vccd1 vccd1 data_out[4] sky130_fd_sc_hd__buf_2
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _5085_/Q _5084_/Q _5083_/Q vssd1 vssd1 vccd1 vccd1 _3931_/A sky130_fd_sc_hd__and3_1
X_3861_ _3861_/A _3861_/B vssd1 vssd1 vccd1 vccd1 _3861_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3792_ _3792_/A vssd1 vssd1 vccd1 vccd1 _3792_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2812_ _2803_/X _2805_/Y _2806_/X _2808_/X _2811_/Y vssd1 vssd1 vccd1 vccd1 _5255_/D
+ sky130_fd_sc_hd__o311a_1
X_2743_ hold15/A _5282_/Q vssd1 vssd1 vccd1 vccd1 _2841_/C sky130_fd_sc_hd__nand2_1
XFILLER_8_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2674_ _4801_/A _5265_/Q vssd1 vssd1 vccd1 vccd1 _2933_/B sky130_fd_sc_hd__nand2_1
X_4413_ _4413_/A _4413_/B vssd1 vssd1 vccd1 vccd1 _4415_/C sky130_fd_sc_hd__nor2_1
X_4344_ _4344_/A _4349_/A vssd1 vssd1 vccd1 vccd1 _4345_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4275_ _4484_/A _4484_/B _4274_/Y vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__o21ai_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _5213_/Q _3190_/X _3224_/Y _3225_/X _3194_/X vssd1 vssd1 vccd1 vccd1 _5213_/D
+ sky130_fd_sc_hd__o221a_1
X_3157_ _2995_/Y _3167_/B _3158_/B _3158_/C vssd1 vssd1 vccd1 vccd1 _3157_/Y sky130_fd_sc_hd__o2bb2ai_1
X_3088_ _3271_/B _3268_/A vssd1 vssd1 vccd1 vccd1 _3088_/X sky130_fd_sc_hd__or2_1
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4060_ _4873_/A _4060_/B _4060_/C vssd1 vssd1 vccd1 vccd1 _5086_/D sky130_fd_sc_hd__nor3_1
X_3011_ _5156_/Q _3686_/B vssd1 vssd1 vccd1 vccd1 _3015_/B sky130_fd_sc_hd__or2_1
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4962_ _5064_/CLK hold19/X vssd1 vssd1 vccd1 vccd1 _4962_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_17_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3913_ _5079_/Q vssd1 vssd1 vccd1 vccd1 _4327_/A sky130_fd_sc_hd__inv_2
X_4893_ _4936_/B vssd1 vssd1 vccd1 vccd1 _4915_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3844_ _3886_/A vssd1 vssd1 vccd1 vccd1 _3844_/X sky130_fd_sc_hd__clkbuf_2
X_3775_ _5123_/Q _3766_/X _3763_/X _3774_/Y vssd1 vssd1 vccd1 vccd1 _5123_/D sky130_fd_sc_hd__o211a_1
X_2726_ _5281_/Q _4543_/A vssd1 vssd1 vccd1 vccd1 _2857_/A sky130_fd_sc_hd__nor2_1
X_2657_ _5261_/Q vssd1 vssd1 vccd1 vccd1 _2966_/B sky130_fd_sc_hd__inv_2
X_2588_ _2594_/A _4811_/A vssd1 vssd1 vccd1 vccd1 _2588_/Y sky130_fd_sc_hd__nand2_1
X_4327_ _4327_/A _4647_/B vssd1 vssd1 vccd1 vccd1 _4329_/A sky130_fd_sc_hd__nand2_1
X_4258_ _4258_/A _4258_/B vssd1 vssd1 vccd1 vccd1 _4259_/B sky130_fd_sc_hd__nor2_1
XFILLER_86_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3209_ _4089_/A vssd1 vssd1 vccd1 vccd1 _4144_/B sky130_fd_sc_hd__buf_4
X_4189_ _4820_/B _5056_/Q vssd1 vssd1 vccd1 vccd1 _4189_/Y sky130_fd_sc_hd__nand2_1
XFILLER_27_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3560_ _3571_/B _3369_/Y _3453_/C _3576_/A vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__o22a_1
X_2511_ _5015_/Q vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__inv_2
X_5230_ _5230_/CLK _5230_/D vssd1 vssd1 vccd1 vccd1 _5230_/Q sky130_fd_sc_hd__dfxtp_1
X_3491_ _5225_/Q vssd1 vssd1 vccd1 vccd1 _3758_/B sky130_fd_sc_hd__inv_2
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5161_ _5228_/CLK _5161_/D vssd1 vssd1 vccd1 vccd1 _5161_/Q sky130_fd_sc_hd__dfxtp_1
X_4112_ _4322_/A _4115_/A _4111_/Y vssd1 vssd1 vccd1 vccd1 _5075_/D sky130_fd_sc_hd__a21oi_1
X_5092_ _5137_/CLK _5092_/D vssd1 vssd1 vccd1 vccd1 _5092_/Q sky130_fd_sc_hd__dfxtp_1
X_4043_ _5067_/Q vssd1 vssd1 vccd1 vccd1 _4283_/A sky130_fd_sc_hd__inv_2
XFILLER_68_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4945_ _4922_/X _4920_/X _4951_/S vssd1 vssd1 vccd1 vccd1 _4945_/X sky130_fd_sc_hd__mux2_1
XFILLER_52_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4876_ _4981_/Q _3898_/B _3897_/B _4986_/Q vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__o22a_1
X_3827_ _3837_/A _3827_/B vssd1 vssd1 vccd1 vccd1 _3827_/Y sky130_fd_sc_hd__nand2_1
X_3758_ _3758_/A _3758_/B vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__nand2_1
X_2709_ _4764_/A _5272_/Q vssd1 vssd1 vccd1 vccd1 _2710_/B sky130_fd_sc_hd__nand2_1
X_3689_ _5155_/Q _3685_/X _3682_/X _3688_/Y vssd1 vssd1 vccd1 vccd1 _5155_/D sky130_fd_sc_hd__o211a_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_87_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2991_ _3668_/A _2991_/B vssd1 vssd1 vccd1 vccd1 _2991_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4730_ _4641_/A _4734_/B _4641_/B vssd1 vssd1 vccd1 vccd1 _4731_/B sky130_fd_sc_hd__o21ba_1
X_4661_ _4661_/A vssd1 vssd1 vccd1 vccd1 _4662_/B sky130_fd_sc_hd__inv_2
X_3612_ _3607_/A _3611_/Y _3577_/X vssd1 vssd1 vccd1 vccd1 _3612_/X sky130_fd_sc_hd__a21o_1
X_4592_ _4796_/A _4800_/B vssd1 vssd1 vccd1 vccd1 _4592_/Y sky130_fd_sc_hd__nand2_1
X_3543_ _3543_/A vssd1 vssd1 vccd1 vccd1 _3557_/A sky130_fd_sc_hd__inv_2
X_3474_ _3372_/Y _3454_/Y _3473_/X vssd1 vssd1 vccd1 vccd1 _3538_/A sky130_fd_sc_hd__o21bai_2
X_5213_ _5213_/CLK _5213_/D vssd1 vssd1 vccd1 vccd1 _5213_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5144_ _5254_/CLK _5144_/D vssd1 vssd1 vccd1 vccd1 _5144_/Q sky130_fd_sc_hd__dfxtp_1
X_5075_ _5076_/CLK _5075_/D vssd1 vssd1 vccd1 vccd1 _5075_/Q sky130_fd_sc_hd__dfxtp_1
X_4026_ _4026_/A _4026_/B vssd1 vssd1 vccd1 vccd1 _4191_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _4936_/B _4931_/B _4928_/C vssd1 vssd1 vccd1 vccd1 _4929_/A sky130_fd_sc_hd__and3_1
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4859_ _4873_/A input7/X vssd1 vssd1 vccd1 vccd1 _4860_/A sky130_fd_sc_hd__or2_1
XFILLER_87_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3190_ _3230_/B vssd1 vssd1 vccd1 vccd1 _3190_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_66_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2974_ _2974_/A vssd1 vssd1 vccd1 vccd1 _2977_/B sky130_fd_sc_hd__inv_2
X_4713_ _4772_/A vssd1 vssd1 vccd1 vccd1 _4713_/X sky130_fd_sc_hd__clkbuf_2
X_4644_ _4719_/A _4719_/B _4643_/X vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__a21oi_1
X_4575_ _4995_/Q _5027_/Q vssd1 vssd1 vccd1 vccd1 _4810_/C sky130_fd_sc_hd__nand2_1
XFILLER_89_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3526_ _3523_/X _3524_/Y _3525_/Y vssd1 vssd1 vccd1 vccd1 _5189_/D sky130_fd_sc_hd__a21oi_1
XFILLER_1_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3457_ _3787_/B _5118_/Q vssd1 vssd1 vccd1 vccd1 _3458_/B sky130_fd_sc_hd__nand2_1
X_3388_ _3827_/B _5103_/Q _3639_/B vssd1 vssd1 vccd1 vccd1 _3388_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5127_ _5193_/CLK _5127_/D vssd1 vssd1 vccd1 vccd1 _5127_/Q sky130_fd_sc_hd__dfxtp_1
X_5058_ _5058_/CLK _5058_/D vssd1 vssd1 vccd1 vccd1 _5058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4009_ _4020_/B _4009_/B _4009_/C vssd1 vssd1 vccd1 vccd1 _4015_/B sky130_fd_sc_hd__nand3_1
XFILLER_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2690_ _5269_/Q _4782_/A vssd1 vssd1 vccd1 vccd1 _2695_/A sky130_fd_sc_hd__nor2_1
XANTENNA_3 _4973_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _4378_/A vssd1 vssd1 vccd1 vccd1 _4360_/Y sky130_fd_sc_hd__inv_2
X_3311_ _3311_/A _3311_/B vssd1 vssd1 vccd1 vccd1 _3311_/Y sky130_fd_sc_hd__nor2_1
X_4291_ _4471_/B _4466_/A vssd1 vssd1 vccd1 vccd1 _4291_/Y sky130_fd_sc_hd__nor2_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _3716_/B _5144_/Q _3241_/X vssd1 vssd1 vccd1 vccd1 _3243_/B sky130_fd_sc_hd__o21a_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _5223_/Q _2972_/X _3171_/Y _3172_/X _2980_/X vssd1 vssd1 vccd1 vccd1 _5223_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_81_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _2957_/A _2957_/B _2957_/C vssd1 vssd1 vccd1 vccd1 _2957_/X sky130_fd_sc_hd__and3_1
XFILLER_41_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2888_ _2893_/B _2893_/A vssd1 vssd1 vccd1 vccd1 _2889_/A sky130_fd_sc_hd__or2_1
X_4627_ _5008_/Q _5040_/Q vssd1 vssd1 vccd1 vccd1 _4748_/A sky130_fd_sc_hd__nor2_1
X_4558_ _5038_/Q vssd1 vssd1 vccd1 vccd1 _4559_/B sky130_fd_sc_hd__inv_2
XFILLER_89_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4489_ _4987_/Q _5032_/Q _4487_/Y _4488_/X _4438_/X vssd1 vssd1 vccd1 vccd1 _5032_/D
+ sky130_fd_sc_hd__o221a_1
X_3509_ _3485_/Y _3488_/Y _3508_/Y vssd1 vssd1 vccd1 vccd1 _3509_/Y sky130_fd_sc_hd__a21oi_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5289_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput51 _5167_/Q vssd1 vssd1 vccd1 vccd1 data_out[5] sky130_fd_sc_hd__buf_2
Xoutput40 _5186_/Q vssd1 vssd1 vccd1 vccd1 data_out[24] sky130_fd_sc_hd__buf_2
XFILLER_0_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5228_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_63_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3860_ _5094_/Q vssd1 vssd1 vccd1 vccd1 _3861_/B sky130_fd_sc_hd__inv_2
X_3791_ _5117_/Q _3779_/X _3789_/X _3790_/Y vssd1 vssd1 vccd1 vccd1 _5117_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2811_ _3238_/A _3676_/B vssd1 vssd1 vccd1 vccd1 _2811_/Y sky130_fd_sc_hd__nand2_1
XFILLER_75_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2742_ _5282_/Q hold15/A vssd1 vssd1 vccd1 vccd1 _2843_/B sky130_fd_sc_hd__or2_1
X_4412_ _4421_/B _4423_/B _4223_/B vssd1 vssd1 vccd1 vccd1 _4413_/B sky130_fd_sc_hd__a21oi_1
XFILLER_8_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2673_ _2673_/A _4998_/Q vssd1 vssd1 vccd1 vccd1 _2678_/A sky130_fd_sc_hd__nand2_1
X_4343_ _4343_/A _4659_/B vssd1 vssd1 vccd1 vccd1 _4349_/A sky130_fd_sc_hd__nor2_1
X_4274_ _4490_/B _4487_/A vssd1 vssd1 vccd1 vccd1 _4274_/Y sky130_fd_sc_hd__nor2_1
X_3225_ _3230_/A _3024_/A _3032_/B _2803_/A vssd1 vssd1 vccd1 vccd1 _3225_/X sky130_fd_sc_hd__a31o_1
XFILLER_67_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ _3672_/B _5161_/Q vssd1 vssd1 vccd1 vccd1 _3158_/C sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_19_clk clkbuf_2_3_0_clk/X vssd1 vssd1 vccd1 vccd1 _5064_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_82_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3087_ _3087_/A vssd1 vssd1 vccd1 vccd1 _3268_/A sky130_fd_sc_hd__inv_2
XFILLER_39_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _4020_/C _4019_/A _4012_/B vssd1 vssd1 vccd1 vccd1 _4026_/B sky130_fd_sc_hd__nand3_1
XFILLER_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3010_ _3010_/A _3015_/A vssd1 vssd1 vccd1 vccd1 _3140_/B sky130_fd_sc_hd__nor2_1
XFILLER_36_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4961_ _5064_/CLK _4961_/D vssd1 vssd1 vccd1 vccd1 hold19/A sky130_fd_sc_hd__dfxtp_1
XFILLER_17_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3912_ _5080_/Q vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__inv_2
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4892_ _4892_/A vssd1 vssd1 vccd1 vccd1 _4936_/B sky130_fd_sc_hd__inv_2
X_3843_ _4501_/A vssd1 vssd1 vccd1 vccd1 _3886_/A sky130_fd_sc_hd__buf_4
X_3774_ _3784_/A _3774_/B vssd1 vssd1 vccd1 vccd1 _3774_/Y sky130_fd_sc_hd__nand2_1
X_2725_ _4543_/A _5281_/Q vssd1 vssd1 vccd1 vccd1 _2857_/B sky130_fd_sc_hd__and2_1
X_2656_ _5263_/Q _4811_/A _2957_/B vssd1 vssd1 vccd1 vccd1 _2656_/Y sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_8_clk _4984_/CLK vssd1 vssd1 vccd1 vccd1 _5281_/CLK sky130_fd_sc_hd__clkbuf_16
X_2587_ _2667_/A vssd1 vssd1 vccd1 vccd1 _4811_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_4326_ _5047_/Q vssd1 vssd1 vccd1 vccd1 _4647_/B sky130_fd_sc_hd__inv_2
X_4257_ _5058_/Q _5026_/Q _4504_/A _4507_/C _4507_/A vssd1 vssd1 vccd1 vccd1 _4494_/A
+ sky130_fd_sc_hd__o2111ai_2
X_4188_ _4178_/B _4185_/Y _4187_/Y vssd1 vssd1 vccd1 vccd1 _4188_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3208_ _3208_/A _3208_/B _3208_/C vssd1 vssd1 vccd1 vccd1 _3208_/Y sky130_fd_sc_hd__nand3_1
X_3139_ _3206_/B _3135_/Y _3138_/Y _3132_/C vssd1 vssd1 vccd1 vccd1 _3196_/C sky130_fd_sc_hd__o22a_1
XFILLER_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3490_ _3502_/B _3502_/A _3507_/A _3489_/Y vssd1 vssd1 vccd1 vccd1 _3504_/B sky130_fd_sc_hd__o22ai_2
X_2510_ _5283_/Q _2506_/X _2507_/X _2509_/Y vssd1 vssd1 vccd1 vccd1 _5283_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5160_ _5228_/CLK _5160_/D vssd1 vssd1 vccd1 vccd1 _5160_/Q sky130_fd_sc_hd__dfxtp_1
X_4111_ _4111_/A _4144_/B vssd1 vssd1 vccd1 vccd1 _4111_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5091_ _5137_/CLK _5091_/D vssd1 vssd1 vccd1 vccd1 _5091_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4042_ _5068_/Q vssd1 vssd1 vccd1 vccd1 _4288_/A sky130_fd_sc_hd__inv_2
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4944_ _4929_/X _4927_/X _4951_/S vssd1 vssd1 vccd1 vccd1 _4944_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4875_ _4925_/B _4984_/Q _4902_/A _4980_/Q _4874_/X vssd1 vssd1 vccd1 vccd1 _4880_/A
+ sky130_fd_sc_hd__o221a_1
X_3826_ _3826_/A vssd1 vssd1 vccd1 vccd1 _3837_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3757_ _5130_/Q _3753_/X _3750_/X _3756_/Y vssd1 vssd1 vccd1 vccd1 _5130_/D sky130_fd_sc_hd__o211a_1
X_2708_ _2708_/A _5005_/Q vssd1 vssd1 vccd1 vccd1 _2900_/B sky130_fd_sc_hd__nand2_1
X_3688_ _3690_/A _3688_/B vssd1 vssd1 vccd1 vccd1 _3688_/Y sky130_fd_sc_hd__nand2_1
X_2639_ _2716_/A vssd1 vssd1 vccd1 vccd1 _2639_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4309_ _4309_/A _4628_/B vssd1 vssd1 vccd1 vccd1 _4445_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5289_ _5289_/CLK _5289_/D vssd1 vssd1 vccd1 vccd1 _5289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_74_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2990_ _5258_/Q _2990_/B vssd1 vssd1 vccd1 vccd1 _2990_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4666_/A _4660_/B vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__nor2_1
XFILLER_14_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3611_ _3611_/A _3611_/B vssd1 vssd1 vccd1 vccd1 _3611_/Y sky130_fd_sc_hd__nand2_1
X_4591_ _4591_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _4800_/B sky130_fd_sc_hd__nor2_1
XFILLER_6_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3542_ _3453_/X _3576_/A _3372_/Y vssd1 vssd1 vccd1 vccd1 _3557_/B sky130_fd_sc_hd__o21bai_1
X_3473_ _3543_/A _3473_/B _3472_/Y vssd1 vssd1 vccd1 vccd1 _3473_/X sky130_fd_sc_hd__or3b_1
XFILLER_69_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5212_ _5215_/CLK _5212_/D vssd1 vssd1 vccd1 vccd1 _5212_/Q sky130_fd_sc_hd__dfxtp_1
X_5143_ _5254_/CLK hold12/X vssd1 vssd1 vccd1 vccd1 _5143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _5074_/CLK _5074_/D vssd1 vssd1 vccd1 vccd1 _5074_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4025_ _4021_/A _4021_/B _4022_/B vssd1 vssd1 vccd1 vccd1 _4025_/X sky130_fd_sc_hd__o21a_1
XFILLER_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4927_ _4927_/A vssd1 vssd1 vccd1 vccd1 _4927_/X sky130_fd_sc_hd__clkbuf_1
X_4858_ _4858_/A vssd1 vssd1 vccd1 vccd1 _4983_/D sky130_fd_sc_hd__clkbuf_1
X_3809_ _5110_/Q _3805_/X _3802_/X _3808_/Y vssd1 vssd1 vccd1 vccd1 _5110_/D sky130_fd_sc_hd__o211a_1
X_4789_ _4793_/B _4596_/A _4596_/B vssd1 vssd1 vccd1 vccd1 _4790_/B sky130_fd_sc_hd__a21bo_1
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_53_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2973_ _4579_/A _5260_/Q vssd1 vssd1 vccd1 vccd1 _2974_/A sky130_fd_sc_hd__nand2_1
X_4712_ _4710_/B _4710_/A _4711_/X vssd1 vssd1 vccd1 vccd1 _4712_/X sky130_fd_sc_hd__a21o_1
X_4643_ _4727_/B _4643_/B _4723_/A vssd1 vssd1 vccd1 vccd1 _4643_/X sky130_fd_sc_hd__or3_1
X_4574_ _4574_/A _4574_/B vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__nand2_1
X_3525_ _5189_/Q _2979_/B _4115_/B vssd1 vssd1 vccd1 vccd1 _3525_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3456_ _5118_/Q _3787_/B vssd1 vssd1 vccd1 vccd1 _3458_/A sky130_fd_sc_hd__or2_1
X_3387_ _5102_/Q _3830_/B vssd1 vssd1 vccd1 vccd1 _3639_/B sky130_fd_sc_hd__or2_1
XFILLER_69_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5126_ _5193_/CLK _5126_/D vssd1 vssd1 vccd1 vccd1 _5126_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5057_ _5058_/CLK _5057_/D vssd1 vssd1 vccd1 vccd1 _5057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4008_ _4192_/B _4022_/A vssd1 vssd1 vccd1 vccd1 _4011_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_4 _4760_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3310_ _3310_/A _3310_/B vssd1 vssd1 vccd1 vccd1 _3311_/B sky130_fd_sc_hd__or2_1
X_4290_ _4290_/A vssd1 vssd1 vccd1 vccd1 _4466_/A sky130_fd_sc_hd__inv_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _3248_/B _3248_/A vssd1 vssd1 vccd1 vccd1 _3241_/X sky130_fd_sc_hd__or2_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3172_ _3148_/Y _3151_/Y _3170_/Y _2866_/X vssd1 vssd1 vccd1 vccd1 _3172_/X sky130_fd_sc_hd__a31o_1
XFILLER_66_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _2957_/A _2957_/B _2957_/C vssd1 vssd1 vccd1 vccd1 _2956_/Y sky130_fd_sc_hd__a21oi_2
X_2887_ _2885_/X _2886_/Y _4873_/A vssd1 vssd1 vccd1 vccd1 _5244_/D sky130_fd_sc_hd__a21oi_1
X_4626_ _4741_/A _4744_/A vssd1 vssd1 vccd1 vccd1 _4634_/A sky130_fd_sc_hd__nand2_1
X_4557_ _4619_/B vssd1 vssd1 vccd1 vccd1 _4557_/Y sky130_fd_sc_hd__inv_2
X_4488_ _4487_/B _4487_/A _4436_/X vssd1 vssd1 vccd1 vccd1 _4488_/X sky130_fd_sc_hd__a21o_1
X_3508_ _3508_/A vssd1 vssd1 vccd1 vccd1 _3508_/Y sky130_fd_sc_hd__inv_2
XFILLER_89_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3439_ _5209_/Q vssd1 vssd1 vccd1 vccd1 _3800_/B sky130_fd_sc_hd__inv_2
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_66_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5109_ _5206_/CLK _5109_/D vssd1 vssd1 vccd1 vccd1 _5109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput52 _5168_/Q vssd1 vssd1 vccd1 vccd1 data_out[6] sky130_fd_sc_hd__buf_2
Xoutput30 _5177_/Q vssd1 vssd1 vccd1 vccd1 data_out[15] sky130_fd_sc_hd__buf_2
Xoutput41 _5187_/Q vssd1 vssd1 vccd1 vccd1 data_out[25] sky130_fd_sc_hd__buf_2
XFILLER_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3790_ _3797_/A _3790_/B vssd1 vssd1 vccd1 vccd1 _3790_/Y sky130_fd_sc_hd__nand2_1
X_2810_ _5255_/Q vssd1 vssd1 vccd1 vccd1 _3676_/B sky130_fd_sc_hd__clkinv_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2741_ _2741_/A _2741_/B vssd1 vssd1 vccd1 vccd1 _2844_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4411_ _4427_/A _4427_/B _4427_/C vssd1 vssd1 vccd1 vccd1 _4421_/B sky130_fd_sc_hd__a21oi_1
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2672_ _5265_/Q vssd1 vssd1 vccd1 vccd1 _2673_/A sky130_fd_sc_hd__inv_2
X_4342_ _5050_/Q vssd1 vssd1 vccd1 vccd1 _4659_/B sky130_fd_sc_hd__inv_2
X_4273_ _4273_/A _4273_/B vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__or2_1
X_3224_ _3230_/A _3032_/B _3024_/A vssd1 vssd1 vccd1 vccd1 _3224_/Y sky130_fd_sc_hd__a21oi_1
.ends

