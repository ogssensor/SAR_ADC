magic
tech sky130A
magscale 1 2
timestamp 1623547275
<< obsli1 >>
rect 1104 1445 178848 117521
<< obsm1 >>
rect 474 756 179570 117552
<< metal2 >>
rect 478 119200 534 120000
rect 1398 119200 1454 120000
rect 2410 119200 2466 120000
rect 3422 119200 3478 120000
rect 4434 119200 4490 120000
rect 5354 119200 5410 120000
rect 6366 119200 6422 120000
rect 7378 119200 7434 120000
rect 8390 119200 8446 120000
rect 9310 119200 9366 120000
rect 10322 119200 10378 120000
rect 11334 119200 11390 120000
rect 12346 119200 12402 120000
rect 13266 119200 13322 120000
rect 14278 119200 14334 120000
rect 15290 119200 15346 120000
rect 16302 119200 16358 120000
rect 17222 119200 17278 120000
rect 18234 119200 18290 120000
rect 19246 119200 19302 120000
rect 20258 119200 20314 120000
rect 21178 119200 21234 120000
rect 22190 119200 22246 120000
rect 23202 119200 23258 120000
rect 24214 119200 24270 120000
rect 25134 119200 25190 120000
rect 26146 119200 26202 120000
rect 27158 119200 27214 120000
rect 28170 119200 28226 120000
rect 29090 119200 29146 120000
rect 30102 119200 30158 120000
rect 31114 119200 31170 120000
rect 32126 119200 32182 120000
rect 33046 119200 33102 120000
rect 34058 119200 34114 120000
rect 35070 119200 35126 120000
rect 36082 119200 36138 120000
rect 37002 119200 37058 120000
rect 38014 119200 38070 120000
rect 39026 119200 39082 120000
rect 40038 119200 40094 120000
rect 40958 119200 41014 120000
rect 41970 119200 42026 120000
rect 42982 119200 43038 120000
rect 43994 119200 44050 120000
rect 44914 119200 44970 120000
rect 45926 119200 45982 120000
rect 46938 119200 46994 120000
rect 47950 119200 48006 120000
rect 48870 119200 48926 120000
rect 49882 119200 49938 120000
rect 50894 119200 50950 120000
rect 51906 119200 51962 120000
rect 52826 119200 52882 120000
rect 53838 119200 53894 120000
rect 54850 119200 54906 120000
rect 55862 119200 55918 120000
rect 56782 119200 56838 120000
rect 57794 119200 57850 120000
rect 58806 119200 58862 120000
rect 59818 119200 59874 120000
rect 60738 119200 60794 120000
rect 61750 119200 61806 120000
rect 62762 119200 62818 120000
rect 63774 119200 63830 120000
rect 64694 119200 64750 120000
rect 65706 119200 65762 120000
rect 66718 119200 66774 120000
rect 67730 119200 67786 120000
rect 68650 119200 68706 120000
rect 69662 119200 69718 120000
rect 70674 119200 70730 120000
rect 71686 119200 71742 120000
rect 72606 119200 72662 120000
rect 73618 119200 73674 120000
rect 74630 119200 74686 120000
rect 75642 119200 75698 120000
rect 76562 119200 76618 120000
rect 77574 119200 77630 120000
rect 78586 119200 78642 120000
rect 79598 119200 79654 120000
rect 80518 119200 80574 120000
rect 81530 119200 81586 120000
rect 82542 119200 82598 120000
rect 83554 119200 83610 120000
rect 84474 119200 84530 120000
rect 85486 119200 85542 120000
rect 86498 119200 86554 120000
rect 87510 119200 87566 120000
rect 88430 119200 88486 120000
rect 89442 119200 89498 120000
rect 90454 119200 90510 120000
rect 91466 119200 91522 120000
rect 92478 119200 92534 120000
rect 93398 119200 93454 120000
rect 94410 119200 94466 120000
rect 95422 119200 95478 120000
rect 96434 119200 96490 120000
rect 97354 119200 97410 120000
rect 98366 119200 98422 120000
rect 99378 119200 99434 120000
rect 100390 119200 100446 120000
rect 101310 119200 101366 120000
rect 102322 119200 102378 120000
rect 103334 119200 103390 120000
rect 104346 119200 104402 120000
rect 105266 119200 105322 120000
rect 106278 119200 106334 120000
rect 107290 119200 107346 120000
rect 108302 119200 108358 120000
rect 109222 119200 109278 120000
rect 110234 119200 110290 120000
rect 111246 119200 111302 120000
rect 112258 119200 112314 120000
rect 113178 119200 113234 120000
rect 114190 119200 114246 120000
rect 115202 119200 115258 120000
rect 116214 119200 116270 120000
rect 117134 119200 117190 120000
rect 118146 119200 118202 120000
rect 119158 119200 119214 120000
rect 120170 119200 120226 120000
rect 121090 119200 121146 120000
rect 122102 119200 122158 120000
rect 123114 119200 123170 120000
rect 124126 119200 124182 120000
rect 125046 119200 125102 120000
rect 126058 119200 126114 120000
rect 127070 119200 127126 120000
rect 128082 119200 128138 120000
rect 129002 119200 129058 120000
rect 130014 119200 130070 120000
rect 131026 119200 131082 120000
rect 132038 119200 132094 120000
rect 132958 119200 133014 120000
rect 133970 119200 134026 120000
rect 134982 119200 135038 120000
rect 135994 119200 136050 120000
rect 136914 119200 136970 120000
rect 137926 119200 137982 120000
rect 138938 119200 138994 120000
rect 139950 119200 140006 120000
rect 140870 119200 140926 120000
rect 141882 119200 141938 120000
rect 142894 119200 142950 120000
rect 143906 119200 143962 120000
rect 144826 119200 144882 120000
rect 145838 119200 145894 120000
rect 146850 119200 146906 120000
rect 147862 119200 147918 120000
rect 148782 119200 148838 120000
rect 149794 119200 149850 120000
rect 150806 119200 150862 120000
rect 151818 119200 151874 120000
rect 152738 119200 152794 120000
rect 153750 119200 153806 120000
rect 154762 119200 154818 120000
rect 155774 119200 155830 120000
rect 156694 119200 156750 120000
rect 157706 119200 157762 120000
rect 158718 119200 158774 120000
rect 159730 119200 159786 120000
rect 160650 119200 160706 120000
rect 161662 119200 161718 120000
rect 162674 119200 162730 120000
rect 163686 119200 163742 120000
rect 164606 119200 164662 120000
rect 165618 119200 165674 120000
rect 166630 119200 166686 120000
rect 167642 119200 167698 120000
rect 168562 119200 168618 120000
rect 169574 119200 169630 120000
rect 170586 119200 170642 120000
rect 171598 119200 171654 120000
rect 172518 119200 172574 120000
rect 173530 119200 173586 120000
rect 174542 119200 174598 120000
rect 175554 119200 175610 120000
rect 176474 119200 176530 120000
rect 177486 119200 177542 120000
rect 178498 119200 178554 120000
rect 179510 119200 179566 120000
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 4526 0 4582 800
rect 5906 0 5962 800
rect 7194 0 7250 800
rect 8482 0 8538 800
rect 9770 0 9826 800
rect 11150 0 11206 800
rect 12438 0 12494 800
rect 13726 0 13782 800
rect 15106 0 15162 800
rect 16394 0 16450 800
rect 17682 0 17738 800
rect 18970 0 19026 800
rect 20350 0 20406 800
rect 21638 0 21694 800
rect 22926 0 22982 800
rect 24306 0 24362 800
rect 25594 0 25650 800
rect 26882 0 26938 800
rect 28170 0 28226 800
rect 29550 0 29606 800
rect 30838 0 30894 800
rect 32126 0 32182 800
rect 33506 0 33562 800
rect 34794 0 34850 800
rect 36082 0 36138 800
rect 37370 0 37426 800
rect 38750 0 38806 800
rect 40038 0 40094 800
rect 41326 0 41382 800
rect 42706 0 42762 800
rect 43994 0 44050 800
rect 45282 0 45338 800
rect 46570 0 46626 800
rect 47950 0 48006 800
rect 49238 0 49294 800
rect 50526 0 50582 800
rect 51906 0 51962 800
rect 53194 0 53250 800
rect 54482 0 54538 800
rect 55770 0 55826 800
rect 57150 0 57206 800
rect 58438 0 58494 800
rect 59726 0 59782 800
rect 61106 0 61162 800
rect 62394 0 62450 800
rect 63682 0 63738 800
rect 64970 0 65026 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68926 0 68982 800
rect 70306 0 70362 800
rect 71594 0 71650 800
rect 72882 0 72938 800
rect 74170 0 74226 800
rect 75550 0 75606 800
rect 76838 0 76894 800
rect 78126 0 78182 800
rect 79506 0 79562 800
rect 80794 0 80850 800
rect 82082 0 82138 800
rect 83370 0 83426 800
rect 84750 0 84806 800
rect 86038 0 86094 800
rect 87326 0 87382 800
rect 88706 0 88762 800
rect 89994 0 90050 800
rect 91282 0 91338 800
rect 92570 0 92626 800
rect 93950 0 94006 800
rect 95238 0 95294 800
rect 96526 0 96582 800
rect 97906 0 97962 800
rect 99194 0 99250 800
rect 100482 0 100538 800
rect 101770 0 101826 800
rect 103150 0 103206 800
rect 104438 0 104494 800
rect 105726 0 105782 800
rect 107106 0 107162 800
rect 108394 0 108450 800
rect 109682 0 109738 800
rect 110970 0 111026 800
rect 112350 0 112406 800
rect 113638 0 113694 800
rect 114926 0 114982 800
rect 116306 0 116362 800
rect 117594 0 117650 800
rect 118882 0 118938 800
rect 120170 0 120226 800
rect 121550 0 121606 800
rect 122838 0 122894 800
rect 124126 0 124182 800
rect 125506 0 125562 800
rect 126794 0 126850 800
rect 128082 0 128138 800
rect 129370 0 129426 800
rect 130750 0 130806 800
rect 132038 0 132094 800
rect 133326 0 133382 800
rect 134706 0 134762 800
rect 135994 0 136050 800
rect 137282 0 137338 800
rect 138570 0 138626 800
rect 139950 0 140006 800
rect 141238 0 141294 800
rect 142526 0 142582 800
rect 143906 0 143962 800
rect 145194 0 145250 800
rect 146482 0 146538 800
rect 147770 0 147826 800
rect 149150 0 149206 800
rect 150438 0 150494 800
rect 151726 0 151782 800
rect 153106 0 153162 800
rect 154394 0 154450 800
rect 155682 0 155738 800
rect 156970 0 157026 800
rect 158350 0 158406 800
rect 159638 0 159694 800
rect 160926 0 160982 800
rect 162306 0 162362 800
rect 163594 0 163650 800
rect 164882 0 164938 800
rect 166170 0 166226 800
rect 167550 0 167606 800
rect 168838 0 168894 800
rect 170126 0 170182 800
rect 171506 0 171562 800
rect 172794 0 172850 800
rect 174082 0 174138 800
rect 175370 0 175426 800
rect 176750 0 176806 800
rect 178038 0 178094 800
rect 179326 0 179382 800
<< obsm2 >>
rect 590 119144 1342 119785
rect 1510 119144 2354 119785
rect 2522 119144 3366 119785
rect 3534 119144 4378 119785
rect 4546 119144 5298 119785
rect 5466 119144 6310 119785
rect 6478 119144 7322 119785
rect 7490 119144 8334 119785
rect 8502 119144 9254 119785
rect 9422 119144 10266 119785
rect 10434 119144 11278 119785
rect 11446 119144 12290 119785
rect 12458 119144 13210 119785
rect 13378 119144 14222 119785
rect 14390 119144 15234 119785
rect 15402 119144 16246 119785
rect 16414 119144 17166 119785
rect 17334 119144 18178 119785
rect 18346 119144 19190 119785
rect 19358 119144 20202 119785
rect 20370 119144 21122 119785
rect 21290 119144 22134 119785
rect 22302 119144 23146 119785
rect 23314 119144 24158 119785
rect 24326 119144 25078 119785
rect 25246 119144 26090 119785
rect 26258 119144 27102 119785
rect 27270 119144 28114 119785
rect 28282 119144 29034 119785
rect 29202 119144 30046 119785
rect 30214 119144 31058 119785
rect 31226 119144 32070 119785
rect 32238 119144 32990 119785
rect 33158 119144 34002 119785
rect 34170 119144 35014 119785
rect 35182 119144 36026 119785
rect 36194 119144 36946 119785
rect 37114 119144 37958 119785
rect 38126 119144 38970 119785
rect 39138 119144 39982 119785
rect 40150 119144 40902 119785
rect 41070 119144 41914 119785
rect 42082 119144 42926 119785
rect 43094 119144 43938 119785
rect 44106 119144 44858 119785
rect 45026 119144 45870 119785
rect 46038 119144 46882 119785
rect 47050 119144 47894 119785
rect 48062 119144 48814 119785
rect 48982 119144 49826 119785
rect 49994 119144 50838 119785
rect 51006 119144 51850 119785
rect 52018 119144 52770 119785
rect 52938 119144 53782 119785
rect 53950 119144 54794 119785
rect 54962 119144 55806 119785
rect 55974 119144 56726 119785
rect 56894 119144 57738 119785
rect 57906 119144 58750 119785
rect 58918 119144 59762 119785
rect 59930 119144 60682 119785
rect 60850 119144 61694 119785
rect 61862 119144 62706 119785
rect 62874 119144 63718 119785
rect 63886 119144 64638 119785
rect 64806 119144 65650 119785
rect 65818 119144 66662 119785
rect 66830 119144 67674 119785
rect 67842 119144 68594 119785
rect 68762 119144 69606 119785
rect 69774 119144 70618 119785
rect 70786 119144 71630 119785
rect 71798 119144 72550 119785
rect 72718 119144 73562 119785
rect 73730 119144 74574 119785
rect 74742 119144 75586 119785
rect 75754 119144 76506 119785
rect 76674 119144 77518 119785
rect 77686 119144 78530 119785
rect 78698 119144 79542 119785
rect 79710 119144 80462 119785
rect 80630 119144 81474 119785
rect 81642 119144 82486 119785
rect 82654 119144 83498 119785
rect 83666 119144 84418 119785
rect 84586 119144 85430 119785
rect 85598 119144 86442 119785
rect 86610 119144 87454 119785
rect 87622 119144 88374 119785
rect 88542 119144 89386 119785
rect 89554 119144 90398 119785
rect 90566 119144 91410 119785
rect 91578 119144 92422 119785
rect 92590 119144 93342 119785
rect 93510 119144 94354 119785
rect 94522 119144 95366 119785
rect 95534 119144 96378 119785
rect 96546 119144 97298 119785
rect 97466 119144 98310 119785
rect 98478 119144 99322 119785
rect 99490 119144 100334 119785
rect 100502 119144 101254 119785
rect 101422 119144 102266 119785
rect 102434 119144 103278 119785
rect 103446 119144 104290 119785
rect 104458 119144 105210 119785
rect 105378 119144 106222 119785
rect 106390 119144 107234 119785
rect 107402 119144 108246 119785
rect 108414 119144 109166 119785
rect 109334 119144 110178 119785
rect 110346 119144 111190 119785
rect 111358 119144 112202 119785
rect 112370 119144 113122 119785
rect 113290 119144 114134 119785
rect 114302 119144 115146 119785
rect 115314 119144 116158 119785
rect 116326 119144 117078 119785
rect 117246 119144 118090 119785
rect 118258 119144 119102 119785
rect 119270 119144 120114 119785
rect 120282 119144 121034 119785
rect 121202 119144 122046 119785
rect 122214 119144 123058 119785
rect 123226 119144 124070 119785
rect 124238 119144 124990 119785
rect 125158 119144 126002 119785
rect 126170 119144 127014 119785
rect 127182 119144 128026 119785
rect 128194 119144 128946 119785
rect 129114 119144 129958 119785
rect 130126 119144 130970 119785
rect 131138 119144 131982 119785
rect 132150 119144 132902 119785
rect 133070 119144 133914 119785
rect 134082 119144 134926 119785
rect 135094 119144 135938 119785
rect 136106 119144 136858 119785
rect 137026 119144 137870 119785
rect 138038 119144 138882 119785
rect 139050 119144 139894 119785
rect 140062 119144 140814 119785
rect 140982 119144 141826 119785
rect 141994 119144 142838 119785
rect 143006 119144 143850 119785
rect 144018 119144 144770 119785
rect 144938 119144 145782 119785
rect 145950 119144 146794 119785
rect 146962 119144 147806 119785
rect 147974 119144 148726 119785
rect 148894 119144 149738 119785
rect 149906 119144 150750 119785
rect 150918 119144 151762 119785
rect 151930 119144 152682 119785
rect 152850 119144 153694 119785
rect 153862 119144 154706 119785
rect 154874 119144 155718 119785
rect 155886 119144 156638 119785
rect 156806 119144 157650 119785
rect 157818 119144 158662 119785
rect 158830 119144 159674 119785
rect 159842 119144 160594 119785
rect 160762 119144 161606 119785
rect 161774 119144 162618 119785
rect 162786 119144 163630 119785
rect 163798 119144 164550 119785
rect 164718 119144 165562 119785
rect 165730 119144 166574 119785
rect 166742 119144 167586 119785
rect 167754 119144 168506 119785
rect 168674 119144 169518 119785
rect 169686 119144 170530 119785
rect 170698 119144 171542 119785
rect 171710 119144 172462 119785
rect 172630 119144 173474 119785
rect 173642 119144 174486 119785
rect 174654 119144 175498 119785
rect 175666 119144 176418 119785
rect 176586 119144 177430 119785
rect 177598 119144 178442 119785
rect 178610 119144 179454 119785
rect 480 856 179564 119144
rect 480 167 606 856
rect 774 167 1894 856
rect 2062 167 3182 856
rect 3350 167 4470 856
rect 4638 167 5850 856
rect 6018 167 7138 856
rect 7306 167 8426 856
rect 8594 167 9714 856
rect 9882 167 11094 856
rect 11262 167 12382 856
rect 12550 167 13670 856
rect 13838 167 15050 856
rect 15218 167 16338 856
rect 16506 167 17626 856
rect 17794 167 18914 856
rect 19082 167 20294 856
rect 20462 167 21582 856
rect 21750 167 22870 856
rect 23038 167 24250 856
rect 24418 167 25538 856
rect 25706 167 26826 856
rect 26994 167 28114 856
rect 28282 167 29494 856
rect 29662 167 30782 856
rect 30950 167 32070 856
rect 32238 167 33450 856
rect 33618 167 34738 856
rect 34906 167 36026 856
rect 36194 167 37314 856
rect 37482 167 38694 856
rect 38862 167 39982 856
rect 40150 167 41270 856
rect 41438 167 42650 856
rect 42818 167 43938 856
rect 44106 167 45226 856
rect 45394 167 46514 856
rect 46682 167 47894 856
rect 48062 167 49182 856
rect 49350 167 50470 856
rect 50638 167 51850 856
rect 52018 167 53138 856
rect 53306 167 54426 856
rect 54594 167 55714 856
rect 55882 167 57094 856
rect 57262 167 58382 856
rect 58550 167 59670 856
rect 59838 167 61050 856
rect 61218 167 62338 856
rect 62506 167 63626 856
rect 63794 167 64914 856
rect 65082 167 66294 856
rect 66462 167 67582 856
rect 67750 167 68870 856
rect 69038 167 70250 856
rect 70418 167 71538 856
rect 71706 167 72826 856
rect 72994 167 74114 856
rect 74282 167 75494 856
rect 75662 167 76782 856
rect 76950 167 78070 856
rect 78238 167 79450 856
rect 79618 167 80738 856
rect 80906 167 82026 856
rect 82194 167 83314 856
rect 83482 167 84694 856
rect 84862 167 85982 856
rect 86150 167 87270 856
rect 87438 167 88650 856
rect 88818 167 89938 856
rect 90106 167 91226 856
rect 91394 167 92514 856
rect 92682 167 93894 856
rect 94062 167 95182 856
rect 95350 167 96470 856
rect 96638 167 97850 856
rect 98018 167 99138 856
rect 99306 167 100426 856
rect 100594 167 101714 856
rect 101882 167 103094 856
rect 103262 167 104382 856
rect 104550 167 105670 856
rect 105838 167 107050 856
rect 107218 167 108338 856
rect 108506 167 109626 856
rect 109794 167 110914 856
rect 111082 167 112294 856
rect 112462 167 113582 856
rect 113750 167 114870 856
rect 115038 167 116250 856
rect 116418 167 117538 856
rect 117706 167 118826 856
rect 118994 167 120114 856
rect 120282 167 121494 856
rect 121662 167 122782 856
rect 122950 167 124070 856
rect 124238 167 125450 856
rect 125618 167 126738 856
rect 126906 167 128026 856
rect 128194 167 129314 856
rect 129482 167 130694 856
rect 130862 167 131982 856
rect 132150 167 133270 856
rect 133438 167 134650 856
rect 134818 167 135938 856
rect 136106 167 137226 856
rect 137394 167 138514 856
rect 138682 167 139894 856
rect 140062 167 141182 856
rect 141350 167 142470 856
rect 142638 167 143850 856
rect 144018 167 145138 856
rect 145306 167 146426 856
rect 146594 167 147714 856
rect 147882 167 149094 856
rect 149262 167 150382 856
rect 150550 167 151670 856
rect 151838 167 153050 856
rect 153218 167 154338 856
rect 154506 167 155626 856
rect 155794 167 156914 856
rect 157082 167 158294 856
rect 158462 167 159582 856
rect 159750 167 160870 856
rect 161038 167 162250 856
rect 162418 167 163538 856
rect 163706 167 164826 856
rect 164994 167 166114 856
rect 166282 167 167494 856
rect 167662 167 168782 856
rect 168950 167 170070 856
rect 170238 167 171450 856
rect 171618 167 172738 856
rect 172906 167 174026 856
rect 174194 167 175314 856
rect 175482 167 176694 856
rect 176862 167 177982 856
rect 178150 167 179270 856
rect 179438 167 179564 856
<< metal3 >>
rect 0 119688 800 119808
rect 0 119416 800 119536
rect 0 119144 800 119264
rect 0 118872 800 118992
rect 0 118600 800 118720
rect 0 118328 800 118448
rect 179200 118192 180000 118312
rect 0 117920 800 118040
rect 0 117648 800 117768
rect 0 117376 800 117496
rect 0 117104 800 117224
rect 0 116832 800 116952
rect 0 116560 800 116680
rect 0 116152 800 116272
rect 0 115880 800 116000
rect 0 115608 800 115728
rect 0 115336 800 115456
rect 0 115064 800 115184
rect 0 114792 800 114912
rect 179200 114928 180000 115048
rect 0 114520 800 114640
rect 0 114112 800 114232
rect 0 113840 800 113960
rect 0 113568 800 113688
rect 0 113296 800 113416
rect 0 113024 800 113144
rect 0 112752 800 112872
rect 0 112344 800 112464
rect 0 112072 800 112192
rect 0 111800 800 111920
rect 0 111528 800 111648
rect 179200 111664 180000 111784
rect 0 111256 800 111376
rect 0 110984 800 111104
rect 0 110576 800 110696
rect 0 110304 800 110424
rect 0 110032 800 110152
rect 0 109760 800 109880
rect 0 109488 800 109608
rect 0 109216 800 109336
rect 0 108944 800 109064
rect 0 108536 800 108656
rect 0 108264 800 108384
rect 179200 108400 180000 108520
rect 0 107992 800 108112
rect 0 107720 800 107840
rect 0 107448 800 107568
rect 0 107176 800 107296
rect 0 106768 800 106888
rect 0 106496 800 106616
rect 0 106224 800 106344
rect 0 105952 800 106072
rect 0 105680 800 105800
rect 0 105408 800 105528
rect 0 105136 800 105256
rect 179200 105136 180000 105256
rect 0 104728 800 104848
rect 0 104456 800 104576
rect 0 104184 800 104304
rect 0 103912 800 104032
rect 0 103640 800 103760
rect 0 103368 800 103488
rect 0 102960 800 103080
rect 0 102688 800 102808
rect 0 102416 800 102536
rect 0 102144 800 102264
rect 0 101872 800 101992
rect 179200 101872 180000 101992
rect 0 101600 800 101720
rect 0 101192 800 101312
rect 0 100920 800 101040
rect 0 100648 800 100768
rect 0 100376 800 100496
rect 0 100104 800 100224
rect 0 99832 800 99952
rect 0 99560 800 99680
rect 0 99152 800 99272
rect 0 98880 800 99000
rect 0 98608 800 98728
rect 179200 98744 180000 98864
rect 0 98336 800 98456
rect 0 98064 800 98184
rect 0 97792 800 97912
rect 0 97384 800 97504
rect 0 97112 800 97232
rect 0 96840 800 96960
rect 0 96568 800 96688
rect 0 96296 800 96416
rect 0 96024 800 96144
rect 0 95752 800 95872
rect 0 95344 800 95464
rect 179200 95480 180000 95600
rect 0 95072 800 95192
rect 0 94800 800 94920
rect 0 94528 800 94648
rect 0 94256 800 94376
rect 0 93984 800 94104
rect 0 93576 800 93696
rect 0 93304 800 93424
rect 0 93032 800 93152
rect 0 92760 800 92880
rect 0 92488 800 92608
rect 0 92216 800 92336
rect 179200 92216 180000 92336
rect 0 91808 800 91928
rect 0 91536 800 91656
rect 0 91264 800 91384
rect 0 90992 800 91112
rect 0 90720 800 90840
rect 0 90448 800 90568
rect 0 90176 800 90296
rect 0 89768 800 89888
rect 0 89496 800 89616
rect 0 89224 800 89344
rect 0 88952 800 89072
rect 179200 88952 180000 89072
rect 0 88680 800 88800
rect 0 88408 800 88528
rect 0 88000 800 88120
rect 0 87728 800 87848
rect 0 87456 800 87576
rect 0 87184 800 87304
rect 0 86912 800 87032
rect 0 86640 800 86760
rect 0 86368 800 86488
rect 0 85960 800 86080
rect 0 85688 800 85808
rect 179200 85688 180000 85808
rect 0 85416 800 85536
rect 0 85144 800 85264
rect 0 84872 800 84992
rect 0 84600 800 84720
rect 0 84192 800 84312
rect 0 83920 800 84040
rect 0 83648 800 83768
rect 0 83376 800 83496
rect 0 83104 800 83224
rect 0 82832 800 82952
rect 0 82424 800 82544
rect 179200 82424 180000 82544
rect 0 82152 800 82272
rect 0 81880 800 82000
rect 0 81608 800 81728
rect 0 81336 800 81456
rect 0 81064 800 81184
rect 0 80792 800 80912
rect 0 80384 800 80504
rect 0 80112 800 80232
rect 0 79840 800 79960
rect 0 79568 800 79688
rect 0 79296 800 79416
rect 179200 79296 180000 79416
rect 0 79024 800 79144
rect 0 78616 800 78736
rect 0 78344 800 78464
rect 0 78072 800 78192
rect 0 77800 800 77920
rect 0 77528 800 77648
rect 0 77256 800 77376
rect 0 76848 800 76968
rect 0 76576 800 76696
rect 0 76304 800 76424
rect 0 76032 800 76152
rect 179200 76032 180000 76152
rect 0 75760 800 75880
rect 0 75488 800 75608
rect 0 75216 800 75336
rect 0 74808 800 74928
rect 0 74536 800 74656
rect 0 74264 800 74384
rect 0 73992 800 74112
rect 0 73720 800 73840
rect 0 73448 800 73568
rect 0 73040 800 73160
rect 0 72768 800 72888
rect 179200 72768 180000 72888
rect 0 72496 800 72616
rect 0 72224 800 72344
rect 0 71952 800 72072
rect 0 71680 800 71800
rect 0 71408 800 71528
rect 0 71000 800 71120
rect 0 70728 800 70848
rect 0 70456 800 70576
rect 0 70184 800 70304
rect 0 69912 800 70032
rect 0 69640 800 69760
rect 179200 69504 180000 69624
rect 0 69232 800 69352
rect 0 68960 800 69080
rect 0 68688 800 68808
rect 0 68416 800 68536
rect 0 68144 800 68264
rect 0 67872 800 67992
rect 0 67464 800 67584
rect 0 67192 800 67312
rect 0 66920 800 67040
rect 0 66648 800 66768
rect 0 66376 800 66496
rect 0 66104 800 66224
rect 179200 66240 180000 66360
rect 0 65832 800 65952
rect 0 65424 800 65544
rect 0 65152 800 65272
rect 0 64880 800 65000
rect 0 64608 800 64728
rect 0 64336 800 64456
rect 0 64064 800 64184
rect 0 63656 800 63776
rect 0 63384 800 63504
rect 0 63112 800 63232
rect 0 62840 800 62960
rect 179200 62976 180000 63096
rect 0 62568 800 62688
rect 0 62296 800 62416
rect 0 62024 800 62144
rect 0 61616 800 61736
rect 0 61344 800 61464
rect 0 61072 800 61192
rect 0 60800 800 60920
rect 0 60528 800 60648
rect 0 60256 800 60376
rect 0 59848 800 59968
rect 179200 59848 180000 59968
rect 0 59576 800 59696
rect 0 59304 800 59424
rect 0 59032 800 59152
rect 0 58760 800 58880
rect 0 58488 800 58608
rect 0 58080 800 58200
rect 0 57808 800 57928
rect 0 57536 800 57656
rect 0 57264 800 57384
rect 0 56992 800 57112
rect 0 56720 800 56840
rect 0 56448 800 56568
rect 179200 56584 180000 56704
rect 0 56040 800 56160
rect 0 55768 800 55888
rect 0 55496 800 55616
rect 0 55224 800 55344
rect 0 54952 800 55072
rect 0 54680 800 54800
rect 0 54272 800 54392
rect 0 54000 800 54120
rect 0 53728 800 53848
rect 0 53456 800 53576
rect 0 53184 800 53304
rect 179200 53320 180000 53440
rect 0 52912 800 53032
rect 0 52640 800 52760
rect 0 52232 800 52352
rect 0 51960 800 52080
rect 0 51688 800 51808
rect 0 51416 800 51536
rect 0 51144 800 51264
rect 0 50872 800 50992
rect 0 50464 800 50584
rect 0 50192 800 50312
rect 0 49920 800 50040
rect 179200 50056 180000 50176
rect 0 49648 800 49768
rect 0 49376 800 49496
rect 0 49104 800 49224
rect 0 48696 800 48816
rect 0 48424 800 48544
rect 0 48152 800 48272
rect 0 47880 800 48000
rect 0 47608 800 47728
rect 0 47336 800 47456
rect 0 47064 800 47184
rect 0 46656 800 46776
rect 179200 46792 180000 46912
rect 0 46384 800 46504
rect 0 46112 800 46232
rect 0 45840 800 45960
rect 0 45568 800 45688
rect 0 45296 800 45416
rect 0 44888 800 45008
rect 0 44616 800 44736
rect 0 44344 800 44464
rect 0 44072 800 44192
rect 0 43800 800 43920
rect 0 43528 800 43648
rect 179200 43528 180000 43648
rect 0 43256 800 43376
rect 0 42848 800 42968
rect 0 42576 800 42696
rect 0 42304 800 42424
rect 0 42032 800 42152
rect 0 41760 800 41880
rect 0 41488 800 41608
rect 0 41080 800 41200
rect 0 40808 800 40928
rect 0 40536 800 40656
rect 0 40264 800 40384
rect 179200 40400 180000 40520
rect 0 39992 800 40112
rect 0 39720 800 39840
rect 0 39312 800 39432
rect 0 39040 800 39160
rect 0 38768 800 38888
rect 0 38496 800 38616
rect 0 38224 800 38344
rect 0 37952 800 38072
rect 0 37680 800 37800
rect 0 37272 800 37392
rect 0 37000 800 37120
rect 179200 37136 180000 37256
rect 0 36728 800 36848
rect 0 36456 800 36576
rect 0 36184 800 36304
rect 0 35912 800 36032
rect 0 35504 800 35624
rect 0 35232 800 35352
rect 0 34960 800 35080
rect 0 34688 800 34808
rect 0 34416 800 34536
rect 0 34144 800 34264
rect 0 33736 800 33856
rect 179200 33872 180000 33992
rect 0 33464 800 33584
rect 0 33192 800 33312
rect 0 32920 800 33040
rect 0 32648 800 32768
rect 0 32376 800 32496
rect 0 32104 800 32224
rect 0 31696 800 31816
rect 0 31424 800 31544
rect 0 31152 800 31272
rect 0 30880 800 31000
rect 0 30608 800 30728
rect 179200 30608 180000 30728
rect 0 30336 800 30456
rect 0 29928 800 30048
rect 0 29656 800 29776
rect 0 29384 800 29504
rect 0 29112 800 29232
rect 0 28840 800 28960
rect 0 28568 800 28688
rect 0 28296 800 28416
rect 0 27888 800 28008
rect 0 27616 800 27736
rect 0 27344 800 27464
rect 179200 27344 180000 27464
rect 0 27072 800 27192
rect 0 26800 800 26920
rect 0 26528 800 26648
rect 0 26120 800 26240
rect 0 25848 800 25968
rect 0 25576 800 25696
rect 0 25304 800 25424
rect 0 25032 800 25152
rect 0 24760 800 24880
rect 0 24352 800 24472
rect 0 24080 800 24200
rect 179200 24080 180000 24200
rect 0 23808 800 23928
rect 0 23536 800 23656
rect 0 23264 800 23384
rect 0 22992 800 23112
rect 0 22720 800 22840
rect 0 22312 800 22432
rect 0 22040 800 22160
rect 0 21768 800 21888
rect 0 21496 800 21616
rect 0 21224 800 21344
rect 0 20952 800 21072
rect 179200 20952 180000 21072
rect 0 20544 800 20664
rect 0 20272 800 20392
rect 0 20000 800 20120
rect 0 19728 800 19848
rect 0 19456 800 19576
rect 0 19184 800 19304
rect 0 18912 800 19032
rect 0 18504 800 18624
rect 0 18232 800 18352
rect 0 17960 800 18080
rect 0 17688 800 17808
rect 179200 17688 180000 17808
rect 0 17416 800 17536
rect 0 17144 800 17264
rect 0 16736 800 16856
rect 0 16464 800 16584
rect 0 16192 800 16312
rect 0 15920 800 16040
rect 0 15648 800 15768
rect 0 15376 800 15496
rect 0 14968 800 15088
rect 0 14696 800 14816
rect 0 14424 800 14544
rect 179200 14424 180000 14544
rect 0 14152 800 14272
rect 0 13880 800 14000
rect 0 13608 800 13728
rect 0 13336 800 13456
rect 0 12928 800 13048
rect 0 12656 800 12776
rect 0 12384 800 12504
rect 0 12112 800 12232
rect 0 11840 800 11960
rect 0 11568 800 11688
rect 0 11160 800 11280
rect 179200 11160 180000 11280
rect 0 10888 800 11008
rect 0 10616 800 10736
rect 0 10344 800 10464
rect 0 10072 800 10192
rect 0 9800 800 9920
rect 0 9528 800 9648
rect 0 9120 800 9240
rect 0 8848 800 8968
rect 0 8576 800 8696
rect 0 8304 800 8424
rect 0 8032 800 8152
rect 0 7760 800 7880
rect 179200 7896 180000 8016
rect 0 7352 800 7472
rect 0 7080 800 7200
rect 0 6808 800 6928
rect 0 6536 800 6656
rect 0 6264 800 6384
rect 0 5992 800 6112
rect 0 5584 800 5704
rect 0 5312 800 5432
rect 0 5040 800 5160
rect 0 4768 800 4888
rect 0 4496 800 4616
rect 179200 4632 180000 4752
rect 0 4224 800 4344
rect 0 3952 800 4072
rect 0 3544 800 3664
rect 0 3272 800 3392
rect 0 3000 800 3120
rect 0 2728 800 2848
rect 0 2456 800 2576
rect 0 2184 800 2304
rect 0 1776 800 1896
rect 0 1504 800 1624
rect 179200 1504 180000 1624
rect 0 1232 800 1352
rect 0 960 800 1080
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
<< obsm3 >>
rect 880 118392 179200 119781
rect 880 118248 179120 118392
rect 800 118120 179120 118248
rect 880 118112 179120 118120
rect 880 116480 179200 118112
rect 800 116352 179200 116480
rect 880 115128 179200 116352
rect 880 114848 179120 115128
rect 880 114440 179200 114848
rect 800 114312 179200 114440
rect 880 112672 179200 114312
rect 800 112544 179200 112672
rect 880 111864 179200 112544
rect 880 111584 179120 111864
rect 880 110904 179200 111584
rect 800 110776 179200 110904
rect 880 108864 179200 110776
rect 800 108736 179200 108864
rect 880 108600 179200 108736
rect 880 108320 179120 108600
rect 880 107096 179200 108320
rect 800 106968 179200 107096
rect 880 105336 179200 106968
rect 880 105056 179120 105336
rect 800 104928 179200 105056
rect 880 103288 179200 104928
rect 800 103160 179200 103288
rect 880 102072 179200 103160
rect 880 101792 179120 102072
rect 880 101520 179200 101792
rect 800 101392 179200 101520
rect 880 99480 179200 101392
rect 800 99352 179200 99480
rect 880 98944 179200 99352
rect 880 98664 179120 98944
rect 880 97712 179200 98664
rect 800 97584 179200 97712
rect 880 95680 179200 97584
rect 880 95672 179120 95680
rect 800 95544 179120 95672
rect 880 95400 179120 95544
rect 880 93904 179200 95400
rect 800 93776 179200 93904
rect 880 92416 179200 93776
rect 880 92136 179120 92416
rect 800 92008 179200 92136
rect 880 90096 179200 92008
rect 800 89968 179200 90096
rect 880 89152 179200 89968
rect 880 88872 179120 89152
rect 880 88328 179200 88872
rect 800 88200 179200 88328
rect 880 86288 179200 88200
rect 800 86160 179200 86288
rect 880 85888 179200 86160
rect 880 85608 179120 85888
rect 880 84520 179200 85608
rect 800 84392 179200 84520
rect 880 82752 179200 84392
rect 800 82624 179200 82752
rect 880 82344 179120 82624
rect 880 80712 179200 82344
rect 800 80584 179200 80712
rect 880 79496 179200 80584
rect 880 79216 179120 79496
rect 880 78944 179200 79216
rect 800 78816 179200 78944
rect 880 77176 179200 78816
rect 800 77048 179200 77176
rect 880 76232 179200 77048
rect 880 75952 179120 76232
rect 880 75136 179200 75952
rect 800 75008 179200 75136
rect 880 73368 179200 75008
rect 800 73240 179200 73368
rect 880 72968 179200 73240
rect 880 72688 179120 72968
rect 880 71328 179200 72688
rect 800 71200 179200 71328
rect 880 69704 179200 71200
rect 880 69560 179120 69704
rect 800 69432 179120 69560
rect 880 69424 179120 69432
rect 880 67792 179200 69424
rect 800 67664 179200 67792
rect 880 66440 179200 67664
rect 880 66160 179120 66440
rect 880 65752 179200 66160
rect 800 65624 179200 65752
rect 880 63984 179200 65624
rect 800 63856 179200 63984
rect 880 63176 179200 63856
rect 880 62896 179120 63176
rect 880 61944 179200 62896
rect 800 61816 179200 61944
rect 880 60176 179200 61816
rect 800 60048 179200 60176
rect 880 59768 179120 60048
rect 880 58408 179200 59768
rect 800 58280 179200 58408
rect 880 56784 179200 58280
rect 880 56504 179120 56784
rect 880 56368 179200 56504
rect 800 56240 179200 56368
rect 880 54600 179200 56240
rect 800 54472 179200 54600
rect 880 53520 179200 54472
rect 880 53240 179120 53520
rect 880 52560 179200 53240
rect 800 52432 179200 52560
rect 880 50792 179200 52432
rect 800 50664 179200 50792
rect 880 50256 179200 50664
rect 880 49976 179120 50256
rect 880 49024 179200 49976
rect 800 48896 179200 49024
rect 880 46992 179200 48896
rect 880 46984 179120 46992
rect 800 46856 179120 46984
rect 880 46712 179120 46856
rect 880 45216 179200 46712
rect 800 45088 179200 45216
rect 880 43728 179200 45088
rect 880 43448 179120 43728
rect 880 43176 179200 43448
rect 800 43048 179200 43176
rect 880 41408 179200 43048
rect 800 41280 179200 41408
rect 880 40600 179200 41280
rect 880 40320 179120 40600
rect 880 39640 179200 40320
rect 800 39512 179200 39640
rect 880 37600 179200 39512
rect 800 37472 179200 37600
rect 880 37336 179200 37472
rect 880 37056 179120 37336
rect 880 35832 179200 37056
rect 800 35704 179200 35832
rect 880 34072 179200 35704
rect 880 34064 179120 34072
rect 800 33936 179120 34064
rect 880 33792 179120 33936
rect 880 32024 179200 33792
rect 800 31896 179200 32024
rect 880 30808 179200 31896
rect 880 30528 179120 30808
rect 880 30256 179200 30528
rect 800 30128 179200 30256
rect 880 28216 179200 30128
rect 800 28088 179200 28216
rect 880 27544 179200 28088
rect 880 27264 179120 27544
rect 880 26448 179200 27264
rect 800 26320 179200 26448
rect 880 24680 179200 26320
rect 800 24552 179200 24680
rect 880 24280 179200 24552
rect 880 24000 179120 24280
rect 880 22640 179200 24000
rect 800 22512 179200 22640
rect 880 21152 179200 22512
rect 880 20872 179120 21152
rect 800 20744 179200 20872
rect 880 18832 179200 20744
rect 800 18704 179200 18832
rect 880 17888 179200 18704
rect 880 17608 179120 17888
rect 880 17064 179200 17608
rect 800 16936 179200 17064
rect 880 15296 179200 16936
rect 800 15168 179200 15296
rect 880 14624 179200 15168
rect 880 14344 179120 14624
rect 880 13256 179200 14344
rect 800 13128 179200 13256
rect 880 11488 179200 13128
rect 800 11360 179200 11488
rect 880 11080 179120 11360
rect 880 9448 179200 11080
rect 800 9320 179200 9448
rect 880 8096 179200 9320
rect 880 7816 179120 8096
rect 880 7680 179200 7816
rect 800 7552 179200 7680
rect 880 5912 179200 7552
rect 800 5784 179200 5912
rect 880 4832 179200 5784
rect 880 4552 179120 4832
rect 880 3872 179200 4552
rect 800 3744 179200 3872
rect 880 2104 179200 3744
rect 800 1976 179200 2104
rect 880 1704 179200 1976
rect 880 1424 179120 1704
rect 880 171 179200 1424
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< labels >>
rlabel metal2 s 478 119200 534 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 30102 119200 30158 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 33046 119200 33102 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 36082 119200 36138 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 39026 119200 39082 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 41970 119200 42026 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 44914 119200 44970 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 47950 119200 48006 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 50894 119200 50950 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 53838 119200 53894 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 56782 119200 56838 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3422 119200 3478 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 59818 119200 59874 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 62762 119200 62818 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 65706 119200 65762 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 68650 119200 68706 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 71686 119200 71742 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 74630 119200 74686 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 77574 119200 77630 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 80518 119200 80574 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 83554 119200 83610 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 86498 119200 86554 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6366 119200 6422 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 89442 119200 89498 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 92478 119200 92534 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 95422 119200 95478 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 98366 119200 98422 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 101310 119200 101366 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 104346 119200 104402 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 107290 119200 107346 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 110234 119200 110290 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9310 119200 9366 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 12346 119200 12402 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 15290 119200 15346 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 18234 119200 18290 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 21178 119200 21234 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 24214 119200 24270 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 27158 119200 27214 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1398 119200 1454 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 31114 119200 31170 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 34058 119200 34114 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 37002 119200 37058 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 40038 119200 40094 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 42982 119200 43038 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 45926 119200 45982 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 48870 119200 48926 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 51906 119200 51962 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 54850 119200 54906 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 57794 119200 57850 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4434 119200 4490 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 60738 119200 60794 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 63774 119200 63830 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 66718 119200 66774 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 69662 119200 69718 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 72606 119200 72662 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 75642 119200 75698 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 78586 119200 78642 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 81530 119200 81586 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 84474 119200 84530 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 87510 119200 87566 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7378 119200 7434 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 90454 119200 90510 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 93398 119200 93454 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 96434 119200 96490 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 99378 119200 99434 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 102322 119200 102378 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 105266 119200 105322 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 108302 119200 108358 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 111246 119200 111302 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10322 119200 10378 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 13266 119200 13322 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 16302 119200 16358 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 19246 119200 19302 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 22190 119200 22246 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 25134 119200 25190 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 28170 119200 28226 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2410 119200 2466 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 32126 119200 32182 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 35070 119200 35126 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 38014 119200 38070 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 40958 119200 41014 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 43994 119200 44050 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 46938 119200 46994 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 49882 119200 49938 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 52826 119200 52882 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 55862 119200 55918 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 58806 119200 58862 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5354 119200 5410 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 61750 119200 61806 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 64694 119200 64750 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 67730 119200 67786 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 70674 119200 70730 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 73618 119200 73674 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 76562 119200 76618 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 79598 119200 79654 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 82542 119200 82598 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 85486 119200 85542 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 88430 119200 88486 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8390 119200 8446 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 91466 119200 91522 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 94410 119200 94466 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 97354 119200 97410 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 100390 119200 100446 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 103334 119200 103390 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 106278 119200 106334 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 109222 119200 109278 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 112258 119200 112314 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11334 119200 11390 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 14278 119200 14334 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 17222 119200 17278 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 20258 119200 20314 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 23202 119200 23258 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 26146 119200 26202 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 29090 119200 29146 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 179200 4632 180000 4752 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 179200 17688 180000 17808 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 145194 0 145250 800 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 0 144 800 264 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 la_data_in[100]
port 119 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 la_data_in[101]
port 120 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 la_data_in[106]
port 125 nsew signal input
rlabel metal3 s 0 94256 800 94376 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 0 95072 800 95192 6 la_data_in[108]
port 127 nsew signal input
rlabel metal3 s 0 96024 800 96144 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 la_data_in[10]
port 129 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 la_data_in[113]
port 133 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 la_data_in[114]
port 134 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 la_data_in[115]
port 135 nsew signal input
rlabel metal3 s 0 102144 800 102264 6 la_data_in[116]
port 136 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 la_data_in[117]
port 137 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 la_data_in[11]
port 140 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal3 s 0 106496 800 106616 6 la_data_in[121]
port 142 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 la_data_in[122]
port 143 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 la_data_in[123]
port 144 nsew signal input
rlabel metal3 s 0 109216 800 109336 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 110032 800 110152 6 la_data_in[125]
port 146 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 10616 800 10736 6 la_data_in[12]
port 149 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 0 12384 800 12504 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 0 15920 800 16040 6 la_data_in[18]
port 155 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 la_data_in[19]
port 156 nsew signal input
rlabel metal3 s 0 960 800 1080 6 la_data_in[1]
port 157 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 la_data_in[21]
port 159 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 0 22992 800 23112 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 la_data_in[28]
port 166 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 la_data_in[29]
port 167 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 la_data_in[2]
port 168 nsew signal input
rlabel metal3 s 0 26528 800 26648 6 la_data_in[30]
port 169 nsew signal input
rlabel metal3 s 0 27344 800 27464 6 la_data_in[31]
port 170 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 la_data_in[32]
port 171 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 la_data_in[33]
port 172 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 la_data_in[35]
port 174 nsew signal input
rlabel metal3 s 0 31696 800 31816 6 la_data_in[36]
port 175 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 la_data_in[38]
port 177 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_data_in[3]
port 179 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 la_data_in[40]
port 180 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 0 37952 800 38072 6 la_data_in[43]
port 183 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 40536 800 40656 6 la_data_in[46]
port 186 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 la_data_in[47]
port 187 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 la_data_in[48]
port 188 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 la_data_in[49]
port 189 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 la_data_in[50]
port 191 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 la_data_in[51]
port 192 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 la_data_in[53]
port 194 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 la_data_in[54]
port 195 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 la_data_in[55]
port 196 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 la_data_in[56]
port 197 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 la_data_in[57]
port 198 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 la_data_in[58]
port 199 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 la_data_in[5]
port 201 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 la_data_in[60]
port 202 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 la_data_in[64]
port 206 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 0 58080 800 58200 6 la_data_in[66]
port 208 nsew signal input
rlabel metal3 s 0 59032 800 59152 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 0 60800 800 60920 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_data_in[71]
port 214 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 la_data_in[72]
port 215 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 la_data_in[73]
port 216 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 la_data_in[74]
port 217 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 la_data_in[75]
port 218 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 0 67872 800 67992 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 0 68688 800 68808 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 la_data_in[7]
port 223 nsew signal input
rlabel metal3 s 0 70456 800 70576 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 la_data_in[82]
port 226 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 la_data_in[84]
port 228 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 la_data_in[88]
port 232 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 la_data_in[89]
port 233 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 la_data_in[8]
port 234 nsew signal input
rlabel metal3 s 0 79296 800 79416 6 la_data_in[90]
port 235 nsew signal input
rlabel metal3 s 0 80112 800 80232 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 la_data_in[92]
port 237 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 la_data_in[93]
port 238 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 la_data_in[99]
port 244 nsew signal input
rlabel metal3 s 0 8032 800 8152 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 416 800 536 6 la_data_out[0]
port 246 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 90176 800 90296 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 0 90992 800 91112 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 92760 800 92880 6 la_data_out[105]
port 252 nsew signal output
rlabel metal3 s 0 93576 800 93696 6 la_data_out[106]
port 253 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 la_data_out[108]
port 255 nsew signal output
rlabel metal3 s 0 96296 800 96416 6 la_data_out[109]
port 256 nsew signal output
rlabel metal3 s 0 9120 800 9240 6 la_data_out[10]
port 257 nsew signal output
rlabel metal3 s 0 97112 800 97232 6 la_data_out[110]
port 258 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 la_data_out[111]
port 259 nsew signal output
rlabel metal3 s 0 98880 800 99000 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 la_data_out[113]
port 261 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 0 102416 800 102536 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 la_data_out[117]
port 265 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 105136 800 105256 6 la_data_out[119]
port 267 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 0 105952 800 106072 6 la_data_out[120]
port 269 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 la_data_out[121]
port 270 nsew signal output
rlabel metal3 s 0 107720 800 107840 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 la_data_out[124]
port 273 nsew signal output
rlabel metal3 s 0 110304 800 110424 6 la_data_out[125]
port 274 nsew signal output
rlabel metal3 s 0 111256 800 111376 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 112072 800 112192 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 0 11840 800 11960 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 la_data_out[15]
port 280 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 la_data_out[16]
port 281 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 0 16192 800 16312 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 la_data_out[19]
port 284 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 0 17960 800 18080 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 la_data_out[21]
port 287 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 0 20544 800 20664 6 la_data_out[23]
port 289 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 la_data_out[24]
port 290 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 0 24080 800 24200 6 la_data_out[27]
port 293 nsew signal output
rlabel metal3 s 0 25032 800 25152 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 la_data_out[2]
port 296 nsew signal output
rlabel metal3 s 0 26800 800 26920 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 la_data_out[31]
port 298 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 la_data_out[32]
port 299 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 la_data_out[33]
port 300 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 la_data_out[34]
port 301 nsew signal output
rlabel metal3 s 0 31152 800 31272 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 32104 800 32224 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 la_data_out[37]
port 304 nsew signal output
rlabel metal3 s 0 33736 800 33856 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 la_data_out[39]
port 306 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 35504 800 35624 6 la_data_out[40]
port 308 nsew signal output
rlabel metal3 s 0 36456 800 36576 6 la_data_out[41]
port 309 nsew signal output
rlabel metal3 s 0 37272 800 37392 6 la_data_out[42]
port 310 nsew signal output
rlabel metal3 s 0 38224 800 38344 6 la_data_out[43]
port 311 nsew signal output
rlabel metal3 s 0 39040 800 39160 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 la_data_out[45]
port 313 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 la_data_out[46]
port 314 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 la_data_out[48]
port 316 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 3952 800 4072 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 la_data_out[50]
port 319 nsew signal output
rlabel metal3 s 0 45296 800 45416 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 46112 800 46232 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 la_data_out[56]
port 325 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 la_data_out[57]
port 326 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 la_data_out[58]
port 327 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 la_data_out[59]
port 328 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 la_data_out[5]
port 329 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 la_data_out[60]
port 330 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 0 56720 800 56840 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 la_data_out[65]
port 335 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 la_data_out[66]
port 336 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 la_data_out[67]
port 337 nsew signal output
rlabel metal3 s 0 60256 800 60376 6 la_data_out[68]
port 338 nsew signal output
rlabel metal3 s 0 61072 800 61192 6 la_data_out[69]
port 339 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 la_data_out[6]
port 340 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 la_data_out[71]
port 342 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 la_data_out[72]
port 343 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 la_data_out[73]
port 344 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 la_data_out[75]
port 346 nsew signal output
rlabel metal3 s 0 67192 800 67312 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 0 68960 800 69080 6 la_data_out[78]
port 349 nsew signal output
rlabel metal3 s 0 69912 800 70032 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 0 6536 800 6656 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 la_data_out[80]
port 352 nsew signal output
rlabel metal3 s 0 71680 800 71800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal3 s 0 72496 800 72616 6 la_data_out[82]
port 354 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 74264 800 74384 6 la_data_out[84]
port 356 nsew signal output
rlabel metal3 s 0 75216 800 75336 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 0 76032 800 76152 6 la_data_out[86]
port 358 nsew signal output
rlabel metal3 s 0 76848 800 76968 6 la_data_out[87]
port 359 nsew signal output
rlabel metal3 s 0 77800 800 77920 6 la_data_out[88]
port 360 nsew signal output
rlabel metal3 s 0 78616 800 78736 6 la_data_out[89]
port 361 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 la_data_out[8]
port 362 nsew signal output
rlabel metal3 s 0 79568 800 79688 6 la_data_out[90]
port 363 nsew signal output
rlabel metal3 s 0 80384 800 80504 6 la_data_out[91]
port 364 nsew signal output
rlabel metal3 s 0 81336 800 81456 6 la_data_out[92]
port 365 nsew signal output
rlabel metal3 s 0 82152 800 82272 6 la_data_out[93]
port 366 nsew signal output
rlabel metal3 s 0 83104 800 83224 6 la_data_out[94]
port 367 nsew signal output
rlabel metal3 s 0 83920 800 84040 6 la_data_out[95]
port 368 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 la_data_out[97]
port 370 nsew signal output
rlabel metal3 s 0 86640 800 86760 6 la_data_out[98]
port 371 nsew signal output
rlabel metal3 s 0 87456 800 87576 6 la_data_out[99]
port 372 nsew signal output
rlabel metal3 s 0 8304 800 8424 6 la_data_out[9]
port 373 nsew signal output
rlabel metal3 s 0 688 800 808 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 0 88680 800 88800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 la_oenb[101]
port 376 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 la_oenb[102]
port 377 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 la_oenb[104]
port 379 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 la_oenb[105]
port 380 nsew signal input
rlabel metal3 s 0 93984 800 94104 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 la_oenb[107]
port 382 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 la_oenb[108]
port 383 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 la_oenb[109]
port 384 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 la_oenb[110]
port 386 nsew signal input
rlabel metal3 s 0 98336 800 98456 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 la_oenb[112]
port 388 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 la_oenb[113]
port 389 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 la_oenb[114]
port 390 nsew signal input
rlabel metal3 s 0 101872 800 101992 6 la_oenb[115]
port 391 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 la_oenb[11]
port 396 nsew signal input
rlabel metal3 s 0 106224 800 106344 6 la_oenb[120]
port 397 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 0 108944 800 109064 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 la_oenb[125]
port 402 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 12112 800 12232 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_oenb[14]
port 407 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 la_oenb[15]
port 408 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_oenb[17]
port 410 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 la_oenb[18]
port 411 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 la_oenb[21]
port 415 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 la_oenb[23]
port 417 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 la_oenb[24]
port 418 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 la_oenb[25]
port 419 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 la_oenb[27]
port 421 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 la_oenb[28]
port 422 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 2456 800 2576 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 la_oenb[30]
port 425 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 la_oenb[31]
port 426 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 la_oenb[32]
port 427 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 0 31424 800 31544 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 la_oenb[36]
port 431 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 0 34144 800 34264 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 34960 800 35080 6 la_oenb[39]
port 434 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 la_oenb[40]
port 436 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 la_oenb[41]
port 437 nsew signal input
rlabel metal3 s 0 37680 800 37800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 la_oenb[44]
port 440 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 la_oenb[45]
port 441 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 la_oenb[46]
port 442 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 la_oenb[4]
port 446 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 la_oenb[50]
port 447 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 46384 800 46504 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 48152 800 48272 6 la_oenb[54]
port 451 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 la_oenb[57]
port 454 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 0 52640 800 52760 6 la_oenb[59]
port 456 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 la_oenb[5]
port 457 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 la_oenb[60]
port 458 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 la_oenb[61]
port 459 nsew signal input
rlabel metal3 s 0 55224 800 55344 6 la_oenb[62]
port 460 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 la_oenb[63]
port 461 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 la_oenb[64]
port 462 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 la_oenb[65]
port 463 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 59576 800 59696 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 64880 800 65000 6 la_oenb[73]
port 472 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 la_oenb[74]
port 473 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 la_oenb[75]
port 474 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 la_oenb[82]
port 482 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 la_oenb[84]
port 484 nsew signal input
rlabel metal3 s 0 75488 800 75608 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 76304 800 76424 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 la_oenb[87]
port 487 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 0 7760 800 7880 6 la_oenb[8]
port 490 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 la_oenb[91]
port 492 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 la_oenb[93]
port 494 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 la_oenb[95]
port 496 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 la_oenb[96]
port 497 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 la_oenb[99]
port 500 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 146850 119200 146906 120000 6 mem_data2_i[0]
port 502 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 mem_data2_i[10]
port 503 nsew signal input
rlabel metal2 s 166630 119200 166686 120000 6 mem_data2_i[11]
port 504 nsew signal input
rlabel metal2 s 167642 119200 167698 120000 6 mem_data2_i[12]
port 505 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 mem_data2_i[13]
port 506 nsew signal input
rlabel metal2 s 169574 119200 169630 120000 6 mem_data2_i[14]
port 507 nsew signal input
rlabel metal3 s 179200 72768 180000 72888 6 mem_data2_i[15]
port 508 nsew signal input
rlabel metal3 s 0 115608 800 115728 6 mem_data2_i[16]
port 509 nsew signal input
rlabel metal3 s 0 115880 800 116000 6 mem_data2_i[17]
port 510 nsew signal input
rlabel metal2 s 172518 119200 172574 120000 6 mem_data2_i[18]
port 511 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 mem_data2_i[19]
port 512 nsew signal input
rlabel metal2 s 148782 119200 148838 120000 6 mem_data2_i[1]
port 513 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 mem_data2_i[20]
port 514 nsew signal input
rlabel metal3 s 179200 82424 180000 82544 6 mem_data2_i[21]
port 515 nsew signal input
rlabel metal2 s 171506 0 171562 800 6 mem_data2_i[22]
port 516 nsew signal input
rlabel metal3 s 179200 88952 180000 89072 6 mem_data2_i[23]
port 517 nsew signal input
rlabel metal2 s 172794 0 172850 800 6 mem_data2_i[24]
port 518 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 mem_data2_i[25]
port 519 nsew signal input
rlabel metal2 s 174082 0 174138 800 6 mem_data2_i[26]
port 520 nsew signal input
rlabel metal2 s 176474 119200 176530 120000 6 mem_data2_i[27]
port 521 nsew signal input
rlabel metal3 s 179200 105136 180000 105256 6 mem_data2_i[28]
port 522 nsew signal input
rlabel metal2 s 176750 0 176806 800 6 mem_data2_i[29]
port 523 nsew signal input
rlabel metal3 s 179200 24080 180000 24200 6 mem_data2_i[2]
port 524 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 mem_data2_i[30]
port 525 nsew signal input
rlabel metal2 s 178498 119200 178554 120000 6 mem_data2_i[31]
port 526 nsew signal input
rlabel metal3 s 179200 30608 180000 30728 6 mem_data2_i[3]
port 527 nsew signal input
rlabel metal3 s 179200 43528 180000 43648 6 mem_data2_i[4]
port 528 nsew signal input
rlabel metal2 s 150438 0 150494 800 6 mem_data2_i[5]
port 529 nsew signal input
rlabel metal2 s 160650 119200 160706 120000 6 mem_data2_i[6]
port 530 nsew signal input
rlabel metal3 s 179200 50056 180000 50176 6 mem_data2_i[7]
port 531 nsew signal input
rlabel metal3 s 0 113840 800 113960 6 mem_data2_i[8]
port 532 nsew signal input
rlabel metal2 s 159638 0 159694 800 6 mem_data2_i[9]
port 533 nsew signal input
rlabel metal3 s 179200 7896 180000 8016 6 mem_data_i[0]
port 534 nsew signal input
rlabel metal2 s 165618 119200 165674 120000 6 mem_data_i[10]
port 535 nsew signal input
rlabel metal3 s 179200 59848 180000 59968 6 mem_data_i[11]
port 536 nsew signal input
rlabel metal2 s 168562 119200 168618 120000 6 mem_data_i[12]
port 537 nsew signal input
rlabel metal3 s 179200 66240 180000 66360 6 mem_data_i[13]
port 538 nsew signal input
rlabel metal2 s 170586 119200 170642 120000 6 mem_data_i[14]
port 539 nsew signal input
rlabel metal2 s 164882 0 164938 800 6 mem_data_i[15]
port 540 nsew signal input
rlabel metal2 s 171598 119200 171654 120000 6 mem_data_i[16]
port 541 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 mem_data_i[17]
port 542 nsew signal input
rlabel metal3 s 179200 79296 180000 79416 6 mem_data_i[18]
port 543 nsew signal input
rlabel metal2 s 174542 119200 174598 120000 6 mem_data_i[19]
port 544 nsew signal input
rlabel metal2 s 149794 119200 149850 120000 6 mem_data_i[1]
port 545 nsew signal input
rlabel metal2 s 175554 119200 175610 120000 6 mem_data_i[20]
port 546 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 mem_data_i[21]
port 547 nsew signal input
rlabel metal3 s 179200 85688 180000 85808 6 mem_data_i[22]
port 548 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 mem_data_i[23]
port 549 nsew signal input
rlabel metal3 s 179200 92216 180000 92336 6 mem_data_i[24]
port 550 nsew signal input
rlabel metal3 s 179200 95480 180000 95600 6 mem_data_i[25]
port 551 nsew signal input
rlabel metal3 s 179200 101872 180000 101992 6 mem_data_i[26]
port 552 nsew signal input
rlabel metal2 s 177486 119200 177542 120000 6 mem_data_i[27]
port 553 nsew signal input
rlabel metal3 s 179200 108400 180000 108520 6 mem_data_i[28]
port 554 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 mem_data_i[29]
port 555 nsew signal input
rlabel metal3 s 0 113024 800 113144 6 mem_data_i[2]
port 556 nsew signal input
rlabel metal3 s 179200 114928 180000 115048 6 mem_data_i[30]
port 557 nsew signal input
rlabel metal2 s 179510 119200 179566 120000 6 mem_data_i[31]
port 558 nsew signal input
rlabel metal2 s 154762 119200 154818 120000 6 mem_data_i[3]
port 559 nsew signal input
rlabel metal3 s 179200 46792 180000 46912 6 mem_data_i[4]
port 560 nsew signal input
rlabel metal2 s 156694 119200 156750 120000 6 mem_data_i[5]
port 561 nsew signal input
rlabel metal2 s 151726 0 151782 800 6 mem_data_i[6]
port 562 nsew signal input
rlabel metal2 s 155682 0 155738 800 6 mem_data_i[7]
port 563 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 mem_data_i[8]
port 564 nsew signal input
rlabel metal2 s 164606 119200 164662 120000 6 mem_data_i[9]
port 565 nsew signal input
rlabel metal2 s 139950 0 140006 800 6 mem_data_o[0]
port 566 nsew signal output
rlabel metal2 s 162306 0 162362 800 6 mem_data_o[10]
port 567 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 mem_data_o[11]
port 568 nsew signal output
rlabel metal3 s 179200 62976 180000 63096 6 mem_data_o[12]
port 569 nsew signal output
rlabel metal3 s 0 115336 800 115456 6 mem_data_o[13]
port 570 nsew signal output
rlabel metal3 s 179200 69504 180000 69624 6 mem_data_o[14]
port 571 nsew signal output
rlabel metal2 s 166170 0 166226 800 6 mem_data_o[15]
port 572 nsew signal output
rlabel metal2 s 167550 0 167606 800 6 mem_data_o[16]
port 573 nsew signal output
rlabel metal3 s 179200 76032 180000 76152 6 mem_data_o[17]
port 574 nsew signal output
rlabel metal2 s 173530 119200 173586 120000 6 mem_data_o[18]
port 575 nsew signal output
rlabel metal3 s 0 116832 800 116952 6 mem_data_o[19]
port 576 nsew signal output
rlabel metal2 s 150806 119200 150862 120000 6 mem_data_o[1]
port 577 nsew signal output
rlabel metal3 s 0 117376 800 117496 6 mem_data_o[20]
port 578 nsew signal output
rlabel metal2 s 170126 0 170182 800 6 mem_data_o[21]
port 579 nsew signal output
rlabel metal3 s 0 117648 800 117768 6 mem_data_o[22]
port 580 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 mem_data_o[23]
port 581 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 mem_data_o[24]
port 582 nsew signal output
rlabel metal3 s 179200 98744 180000 98864 6 mem_data_o[25]
port 583 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 mem_data_o[26]
port 584 nsew signal output
rlabel metal2 s 175370 0 175426 800 6 mem_data_o[27]
port 585 nsew signal output
rlabel metal3 s 179200 111664 180000 111784 6 mem_data_o[28]
port 586 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 mem_data_o[29]
port 587 nsew signal output
rlabel metal2 s 151818 119200 151874 120000 6 mem_data_o[2]
port 588 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 mem_data_o[30]
port 589 nsew signal output
rlabel metal3 s 179200 118192 180000 118312 6 mem_data_o[31]
port 590 nsew signal output
rlabel metal3 s 179200 33872 180000 33992 6 mem_data_o[3]
port 591 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 mem_data_o[4]
port 592 nsew signal output
rlabel metal2 s 157706 119200 157762 120000 6 mem_data_o[5]
port 593 nsew signal output
rlabel metal2 s 153106 0 153162 800 6 mem_data_o[6]
port 594 nsew signal output
rlabel metal2 s 161662 119200 161718 120000 6 mem_data_o[7]
port 595 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 mem_data_o[8]
port 596 nsew signal output
rlabel metal3 s 179200 56584 180000 56704 6 mem_data_o[9]
port 597 nsew signal output
rlabel metal2 s 147862 119200 147918 120000 6 mem_raddr_o[0]
port 598 nsew signal output
rlabel metal2 s 141238 0 141294 800 6 mem_raddr_o[1]
port 599 nsew signal output
rlabel metal3 s 0 113296 800 113416 6 mem_raddr_o[2]
port 600 nsew signal output
rlabel metal3 s 179200 37136 180000 37256 6 mem_raddr_o[3]
port 601 nsew signal output
rlabel metal2 s 155774 119200 155830 120000 6 mem_raddr_o[4]
port 602 nsew signal output
rlabel metal2 s 158718 119200 158774 120000 6 mem_raddr_o[5]
port 603 nsew signal output
rlabel metal3 s 0 113568 800 113688 6 mem_raddr_o[6]
port 604 nsew signal output
rlabel metal2 s 162674 119200 162730 120000 6 mem_raddr_o[7]
port 605 nsew signal output
rlabel metal3 s 179200 53320 180000 53440 6 mem_raddr_o[8]
port 606 nsew signal output
rlabel metal3 s 0 114520 800 114640 6 mem_raddr_o[9]
port 607 nsew signal output
rlabel metal3 s 179200 1504 180000 1624 6 mem_renb_o
port 608 nsew signal output
rlabel metal3 s 179200 11160 180000 11280 6 mem_waddr_o[0]
port 609 nsew signal output
rlabel metal2 s 142526 0 142582 800 6 mem_waddr_o[1]
port 610 nsew signal output
rlabel metal2 s 152738 119200 152794 120000 6 mem_waddr_o[2]
port 611 nsew signal output
rlabel metal2 s 146482 0 146538 800 6 mem_waddr_o[3]
port 612 nsew signal output
rlabel metal2 s 149150 0 149206 800 6 mem_waddr_o[4]
port 613 nsew signal output
rlabel metal2 s 159730 119200 159786 120000 6 mem_waddr_o[5]
port 614 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 mem_waddr_o[6]
port 615 nsew signal output
rlabel metal2 s 163686 119200 163742 120000 6 mem_waddr_o[7]
port 616 nsew signal output
rlabel metal2 s 158350 0 158406 800 6 mem_waddr_o[8]
port 617 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 mem_waddr_o[9]
port 618 nsew signal output
rlabel metal2 s 145838 119200 145894 120000 6 mem_wenb_o
port 619 nsew signal output
rlabel metal2 s 113178 119200 113234 120000 6 phase0_in[0]
port 620 nsew signal input
rlabel metal2 s 142894 119200 142950 120000 6 phase0_in[10]
port 621 nsew signal input
rlabel metal2 s 116214 119200 116270 120000 6 phase0_in[1]
port 622 nsew signal input
rlabel metal2 s 119158 119200 119214 120000 6 phase0_in[2]
port 623 nsew signal input
rlabel metal2 s 122102 119200 122158 120000 6 phase0_in[3]
port 624 nsew signal input
rlabel metal2 s 125046 119200 125102 120000 6 phase0_in[4]
port 625 nsew signal input
rlabel metal2 s 128082 119200 128138 120000 6 phase0_in[5]
port 626 nsew signal input
rlabel metal2 s 131026 119200 131082 120000 6 phase0_in[6]
port 627 nsew signal input
rlabel metal2 s 133970 119200 134026 120000 6 phase0_in[7]
port 628 nsew signal input
rlabel metal2 s 136914 119200 136970 120000 6 phase0_in[8]
port 629 nsew signal input
rlabel metal2 s 139950 119200 140006 120000 6 phase0_in[9]
port 630 nsew signal input
rlabel metal2 s 114190 119200 114246 120000 6 phase1_in[0]
port 631 nsew signal input
rlabel metal2 s 143906 119200 143962 120000 6 phase1_in[10]
port 632 nsew signal input
rlabel metal2 s 117134 119200 117190 120000 6 phase1_in[1]
port 633 nsew signal input
rlabel metal2 s 120170 119200 120226 120000 6 phase1_in[2]
port 634 nsew signal input
rlabel metal2 s 123114 119200 123170 120000 6 phase1_in[3]
port 635 nsew signal input
rlabel metal2 s 126058 119200 126114 120000 6 phase1_in[4]
port 636 nsew signal input
rlabel metal2 s 129002 119200 129058 120000 6 phase1_in[5]
port 637 nsew signal input
rlabel metal2 s 132038 119200 132094 120000 6 phase1_in[6]
port 638 nsew signal input
rlabel metal2 s 134982 119200 135038 120000 6 phase1_in[7]
port 639 nsew signal input
rlabel metal2 s 137926 119200 137982 120000 6 phase1_in[8]
port 640 nsew signal input
rlabel metal2 s 140870 119200 140926 120000 6 phase1_in[9]
port 641 nsew signal input
rlabel metal2 s 115202 119200 115258 120000 6 phase2_in[0]
port 642 nsew signal input
rlabel metal2 s 144826 119200 144882 120000 6 phase2_in[10]
port 643 nsew signal input
rlabel metal2 s 118146 119200 118202 120000 6 phase2_in[1]
port 644 nsew signal input
rlabel metal2 s 121090 119200 121146 120000 6 phase2_in[2]
port 645 nsew signal input
rlabel metal2 s 124126 119200 124182 120000 6 phase2_in[3]
port 646 nsew signal input
rlabel metal2 s 127070 119200 127126 120000 6 phase2_in[4]
port 647 nsew signal input
rlabel metal2 s 130014 119200 130070 120000 6 phase2_in[5]
port 648 nsew signal input
rlabel metal2 s 132958 119200 133014 120000 6 phase2_in[6]
port 649 nsew signal input
rlabel metal2 s 135994 119200 136050 120000 6 phase2_in[7]
port 650 nsew signal input
rlabel metal2 s 138938 119200 138994 120000 6 phase2_in[8]
port 651 nsew signal input
rlabel metal2 s 141882 119200 141938 120000 6 phase2_in[9]
port 652 nsew signal input
rlabel metal3 s 179200 14424 180000 14544 6 vco_enb_o[0]
port 653 nsew signal output
rlabel metal2 s 143906 0 143962 800 6 vco_enb_o[1]
port 654 nsew signal output
rlabel metal2 s 153750 119200 153806 120000 6 vco_enb_o[2]
port 655 nsew signal output
rlabel metal2 s 662 0 718 800 6 wb_clk_i
port 656 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wb_rst_i
port 657 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_ack_o
port 658 nsew signal output
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[0]
port 659 nsew signal input
rlabel metal2 s 53194 0 53250 800 6 wbs_adr_i[10]
port 660 nsew signal input
rlabel metal2 s 57150 0 57206 800 6 wbs_adr_i[11]
port 661 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 wbs_adr_i[12]
port 662 nsew signal input
rlabel metal2 s 64970 0 65026 800 6 wbs_adr_i[13]
port 663 nsew signal input
rlabel metal2 s 68926 0 68982 800 6 wbs_adr_i[14]
port 664 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 wbs_adr_i[15]
port 665 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 wbs_adr_i[16]
port 666 nsew signal input
rlabel metal2 s 80794 0 80850 800 6 wbs_adr_i[17]
port 667 nsew signal input
rlabel metal2 s 84750 0 84806 800 6 wbs_adr_i[18]
port 668 nsew signal input
rlabel metal2 s 88706 0 88762 800 6 wbs_adr_i[19]
port 669 nsew signal input
rlabel metal2 s 13726 0 13782 800 6 wbs_adr_i[1]
port 670 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 wbs_adr_i[20]
port 671 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 wbs_adr_i[21]
port 672 nsew signal input
rlabel metal2 s 100482 0 100538 800 6 wbs_adr_i[22]
port 673 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_adr_i[23]
port 674 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 wbs_adr_i[24]
port 675 nsew signal input
rlabel metal2 s 112350 0 112406 800 6 wbs_adr_i[25]
port 676 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 wbs_adr_i[26]
port 677 nsew signal input
rlabel metal2 s 120170 0 120226 800 6 wbs_adr_i[27]
port 678 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 wbs_adr_i[28]
port 679 nsew signal input
rlabel metal2 s 128082 0 128138 800 6 wbs_adr_i[29]
port 680 nsew signal input
rlabel metal2 s 18970 0 19026 800 6 wbs_adr_i[2]
port 681 nsew signal input
rlabel metal2 s 132038 0 132094 800 6 wbs_adr_i[30]
port 682 nsew signal input
rlabel metal2 s 135994 0 136050 800 6 wbs_adr_i[31]
port 683 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_adr_i[3]
port 684 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[4]
port 685 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 wbs_adr_i[5]
port 686 nsew signal input
rlabel metal2 s 37370 0 37426 800 6 wbs_adr_i[6]
port 687 nsew signal input
rlabel metal2 s 41326 0 41382 800 6 wbs_adr_i[7]
port 688 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 wbs_adr_i[8]
port 689 nsew signal input
rlabel metal2 s 49238 0 49294 800 6 wbs_adr_i[9]
port 690 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_cyc_i
port 691 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 wbs_dat_i[0]
port 692 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 wbs_dat_i[10]
port 693 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 wbs_dat_i[11]
port 694 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 wbs_dat_i[12]
port 695 nsew signal input
rlabel metal2 s 66350 0 66406 800 6 wbs_dat_i[13]
port 696 nsew signal input
rlabel metal2 s 70306 0 70362 800 6 wbs_dat_i[14]
port 697 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 wbs_dat_i[15]
port 698 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 wbs_dat_i[16]
port 699 nsew signal input
rlabel metal2 s 82082 0 82138 800 6 wbs_dat_i[17]
port 700 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 wbs_dat_i[18]
port 701 nsew signal input
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_i[19]
port 702 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[1]
port 703 nsew signal input
rlabel metal2 s 93950 0 94006 800 6 wbs_dat_i[20]
port 704 nsew signal input
rlabel metal2 s 97906 0 97962 800 6 wbs_dat_i[21]
port 705 nsew signal input
rlabel metal2 s 101770 0 101826 800 6 wbs_dat_i[22]
port 706 nsew signal input
rlabel metal2 s 105726 0 105782 800 6 wbs_dat_i[23]
port 707 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 wbs_dat_i[24]
port 708 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 wbs_dat_i[25]
port 709 nsew signal input
rlabel metal2 s 117594 0 117650 800 6 wbs_dat_i[26]
port 710 nsew signal input
rlabel metal2 s 121550 0 121606 800 6 wbs_dat_i[27]
port 711 nsew signal input
rlabel metal2 s 125506 0 125562 800 6 wbs_dat_i[28]
port 712 nsew signal input
rlabel metal2 s 129370 0 129426 800 6 wbs_dat_i[29]
port 713 nsew signal input
rlabel metal2 s 20350 0 20406 800 6 wbs_dat_i[2]
port 714 nsew signal input
rlabel metal2 s 133326 0 133382 800 6 wbs_dat_i[30]
port 715 nsew signal input
rlabel metal2 s 137282 0 137338 800 6 wbs_dat_i[31]
port 716 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 wbs_dat_i[3]
port 717 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_dat_i[4]
port 718 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_i[5]
port 719 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 wbs_dat_i[6]
port 720 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 wbs_dat_i[7]
port 721 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 wbs_dat_i[8]
port 722 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_dat_i[9]
port 723 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[0]
port 724 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 wbs_dat_o[10]
port 725 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_o[11]
port 726 nsew signal output
rlabel metal2 s 63682 0 63738 800 6 wbs_dat_o[12]
port 727 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_o[13]
port 728 nsew signal output
rlabel metal2 s 71594 0 71650 800 6 wbs_dat_o[14]
port 729 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_o[15]
port 730 nsew signal output
rlabel metal2 s 79506 0 79562 800 6 wbs_dat_o[16]
port 731 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 wbs_dat_o[17]
port 732 nsew signal output
rlabel metal2 s 87326 0 87382 800 6 wbs_dat_o[18]
port 733 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 wbs_dat_o[19]
port 734 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 wbs_dat_o[1]
port 735 nsew signal output
rlabel metal2 s 95238 0 95294 800 6 wbs_dat_o[20]
port 736 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 wbs_dat_o[21]
port 737 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 wbs_dat_o[22]
port 738 nsew signal output
rlabel metal2 s 107106 0 107162 800 6 wbs_dat_o[23]
port 739 nsew signal output
rlabel metal2 s 110970 0 111026 800 6 wbs_dat_o[24]
port 740 nsew signal output
rlabel metal2 s 114926 0 114982 800 6 wbs_dat_o[25]
port 741 nsew signal output
rlabel metal2 s 118882 0 118938 800 6 wbs_dat_o[26]
port 742 nsew signal output
rlabel metal2 s 122838 0 122894 800 6 wbs_dat_o[27]
port 743 nsew signal output
rlabel metal2 s 126794 0 126850 800 6 wbs_dat_o[28]
port 744 nsew signal output
rlabel metal2 s 130750 0 130806 800 6 wbs_dat_o[29]
port 745 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[2]
port 746 nsew signal output
rlabel metal2 s 134706 0 134762 800 6 wbs_dat_o[30]
port 747 nsew signal output
rlabel metal2 s 138570 0 138626 800 6 wbs_dat_o[31]
port 748 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 wbs_dat_o[3]
port 749 nsew signal output
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_o[4]
port 750 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_o[5]
port 751 nsew signal output
rlabel metal2 s 40038 0 40094 800 6 wbs_dat_o[6]
port 752 nsew signal output
rlabel metal2 s 43994 0 44050 800 6 wbs_dat_o[7]
port 753 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 wbs_dat_o[8]
port 754 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 wbs_dat_o[9]
port 755 nsew signal output
rlabel metal2 s 12438 0 12494 800 6 wbs_sel_i[0]
port 756 nsew signal input
rlabel metal2 s 17682 0 17738 800 6 wbs_sel_i[1]
port 757 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_sel_i[2]
port 758 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 wbs_sel_i[3]
port 759 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_stb_i
port 760 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_we_i
port 761 nsew signal input
rlabel metal3 s 0 112752 800 112872 6 wmask_o[0]
port 762 nsew signal output
rlabel metal3 s 179200 20952 180000 21072 6 wmask_o[1]
port 763 nsew signal output
rlabel metal3 s 179200 27344 180000 27464 6 wmask_o[2]
port 764 nsew signal output
rlabel metal3 s 179200 40400 180000 40520 6 wmask_o[3]
port 765 nsew signal output
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 766 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 767 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 768 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 770 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 771 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 772 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 773 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 775 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 776 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 777 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 778 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 779 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 780 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 781 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 782 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 783 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 784 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 785 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 786 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 787 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 788 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 789 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 790 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 791 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 792 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 793 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 794 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 795 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 796 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 797 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 798 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 799 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 800 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 801 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 802 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 803 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 804 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 805 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 806 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 807 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 808 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 809 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 810 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 811 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 812 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 813 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 14604816
string GDS_START 978752
<< end >>

