magic
tech sky130A
magscale 1 2
timestamp 1624086562
<< obsli1 >>
rect 1104 1377 178848 117521
<< obsm1 >>
rect 566 892 179386 117552
<< metal2 >>
rect 570 119200 626 120000
rect 1766 119200 1822 120000
rect 2962 119200 3018 120000
rect 4250 119200 4306 120000
rect 5446 119200 5502 120000
rect 6734 119200 6790 120000
rect 7930 119200 7986 120000
rect 9126 119200 9182 120000
rect 10414 119200 10470 120000
rect 11610 119200 11666 120000
rect 12898 119200 12954 120000
rect 14094 119200 14150 120000
rect 15290 119200 15346 120000
rect 16578 119200 16634 120000
rect 17774 119200 17830 120000
rect 19062 119200 19118 120000
rect 20258 119200 20314 120000
rect 21454 119200 21510 120000
rect 22742 119200 22798 120000
rect 23938 119200 23994 120000
rect 25226 119200 25282 120000
rect 26422 119200 26478 120000
rect 27618 119200 27674 120000
rect 28906 119200 28962 120000
rect 30102 119200 30158 120000
rect 31390 119200 31446 120000
rect 32586 119200 32642 120000
rect 33782 119200 33838 120000
rect 35070 119200 35126 120000
rect 36266 119200 36322 120000
rect 37554 119200 37610 120000
rect 38750 119200 38806 120000
rect 39946 119200 40002 120000
rect 41234 119200 41290 120000
rect 42430 119200 42486 120000
rect 43718 119200 43774 120000
rect 44914 119200 44970 120000
rect 46110 119200 46166 120000
rect 47398 119200 47454 120000
rect 48594 119200 48650 120000
rect 49882 119200 49938 120000
rect 51078 119200 51134 120000
rect 52274 119200 52330 120000
rect 53562 119200 53618 120000
rect 54758 119200 54814 120000
rect 56046 119200 56102 120000
rect 57242 119200 57298 120000
rect 58438 119200 58494 120000
rect 59726 119200 59782 120000
rect 60922 119200 60978 120000
rect 62210 119200 62266 120000
rect 63406 119200 63462 120000
rect 64694 119200 64750 120000
rect 65890 119200 65946 120000
rect 67086 119200 67142 120000
rect 68374 119200 68430 120000
rect 69570 119200 69626 120000
rect 70858 119200 70914 120000
rect 72054 119200 72110 120000
rect 73250 119200 73306 120000
rect 74538 119200 74594 120000
rect 75734 119200 75790 120000
rect 77022 119200 77078 120000
rect 78218 119200 78274 120000
rect 79414 119200 79470 120000
rect 80702 119200 80758 120000
rect 81898 119200 81954 120000
rect 83186 119200 83242 120000
rect 84382 119200 84438 120000
rect 85578 119200 85634 120000
rect 86866 119200 86922 120000
rect 88062 119200 88118 120000
rect 89350 119200 89406 120000
rect 90546 119200 90602 120000
rect 91742 119200 91798 120000
rect 93030 119200 93086 120000
rect 94226 119200 94282 120000
rect 95514 119200 95570 120000
rect 96710 119200 96766 120000
rect 97906 119200 97962 120000
rect 99194 119200 99250 120000
rect 100390 119200 100446 120000
rect 101678 119200 101734 120000
rect 102874 119200 102930 120000
rect 104070 119200 104126 120000
rect 105358 119200 105414 120000
rect 106554 119200 106610 120000
rect 107842 119200 107898 120000
rect 109038 119200 109094 120000
rect 110234 119200 110290 120000
rect 111522 119200 111578 120000
rect 112718 119200 112774 120000
rect 114006 119200 114062 120000
rect 115202 119200 115258 120000
rect 116398 119200 116454 120000
rect 117686 119200 117742 120000
rect 118882 119200 118938 120000
rect 120170 119200 120226 120000
rect 121366 119200 121422 120000
rect 122654 119200 122710 120000
rect 123850 119200 123906 120000
rect 125046 119200 125102 120000
rect 126334 119200 126390 120000
rect 127530 119200 127586 120000
rect 128818 119200 128874 120000
rect 130014 119200 130070 120000
rect 131210 119200 131266 120000
rect 132498 119200 132554 120000
rect 133694 119200 133750 120000
rect 134982 119200 135038 120000
rect 136178 119200 136234 120000
rect 137374 119200 137430 120000
rect 138662 119200 138718 120000
rect 139858 119200 139914 120000
rect 141146 119200 141202 120000
rect 142342 119200 142398 120000
rect 143538 119200 143594 120000
rect 144826 119200 144882 120000
rect 146022 119200 146078 120000
rect 147310 119200 147366 120000
rect 148506 119200 148562 120000
rect 149702 119200 149758 120000
rect 150990 119200 151046 120000
rect 152186 119200 152242 120000
rect 153474 119200 153530 120000
rect 154670 119200 154726 120000
rect 155866 119200 155922 120000
rect 157154 119200 157210 120000
rect 158350 119200 158406 120000
rect 159638 119200 159694 120000
rect 160834 119200 160890 120000
rect 162030 119200 162086 120000
rect 163318 119200 163374 120000
rect 164514 119200 164570 120000
rect 165802 119200 165858 120000
rect 166998 119200 167054 120000
rect 168194 119200 168250 120000
rect 169482 119200 169538 120000
rect 170678 119200 170734 120000
rect 171966 119200 172022 120000
rect 173162 119200 173218 120000
rect 174358 119200 174414 120000
rect 175646 119200 175702 120000
rect 176842 119200 176898 120000
rect 178130 119200 178186 120000
rect 179326 119200 179382 120000
rect 754 0 810 800
rect 2226 0 2282 800
rect 3698 0 3754 800
rect 5170 0 5226 800
rect 6642 0 6698 800
rect 8114 0 8170 800
rect 9678 0 9734 800
rect 11150 0 11206 800
rect 12622 0 12678 800
rect 14094 0 14150 800
rect 15566 0 15622 800
rect 17038 0 17094 800
rect 18602 0 18658 800
rect 20074 0 20130 800
rect 21546 0 21602 800
rect 23018 0 23074 800
rect 24490 0 24546 800
rect 25962 0 26018 800
rect 27526 0 27582 800
rect 28998 0 29054 800
rect 30470 0 30526 800
rect 31942 0 31998 800
rect 33414 0 33470 800
rect 34886 0 34942 800
rect 36450 0 36506 800
rect 37922 0 37978 800
rect 39394 0 39450 800
rect 40866 0 40922 800
rect 42338 0 42394 800
rect 43902 0 43958 800
rect 45374 0 45430 800
rect 46846 0 46902 800
rect 48318 0 48374 800
rect 49790 0 49846 800
rect 51262 0 51318 800
rect 52826 0 52882 800
rect 54298 0 54354 800
rect 55770 0 55826 800
rect 57242 0 57298 800
rect 58714 0 58770 800
rect 60186 0 60242 800
rect 61750 0 61806 800
rect 63222 0 63278 800
rect 64694 0 64750 800
rect 66166 0 66222 800
rect 67638 0 67694 800
rect 69110 0 69166 800
rect 70674 0 70730 800
rect 72146 0 72202 800
rect 73618 0 73674 800
rect 75090 0 75146 800
rect 76562 0 76618 800
rect 78126 0 78182 800
rect 79598 0 79654 800
rect 81070 0 81126 800
rect 82542 0 82598 800
rect 84014 0 84070 800
rect 85486 0 85542 800
rect 87050 0 87106 800
rect 88522 0 88578 800
rect 89994 0 90050 800
rect 91466 0 91522 800
rect 92938 0 92994 800
rect 94410 0 94466 800
rect 95974 0 96030 800
rect 97446 0 97502 800
rect 98918 0 98974 800
rect 100390 0 100446 800
rect 101862 0 101918 800
rect 103334 0 103390 800
rect 104898 0 104954 800
rect 106370 0 106426 800
rect 107842 0 107898 800
rect 109314 0 109370 800
rect 110786 0 110842 800
rect 112350 0 112406 800
rect 113822 0 113878 800
rect 115294 0 115350 800
rect 116766 0 116822 800
rect 118238 0 118294 800
rect 119710 0 119766 800
rect 121274 0 121330 800
rect 122746 0 122802 800
rect 124218 0 124274 800
rect 125690 0 125746 800
rect 127162 0 127218 800
rect 128634 0 128690 800
rect 130198 0 130254 800
rect 131670 0 131726 800
rect 133142 0 133198 800
rect 134614 0 134670 800
rect 136086 0 136142 800
rect 137558 0 137614 800
rect 139122 0 139178 800
rect 140594 0 140650 800
rect 142066 0 142122 800
rect 143538 0 143594 800
rect 145010 0 145066 800
rect 146574 0 146630 800
rect 148046 0 148102 800
rect 149518 0 149574 800
rect 150990 0 151046 800
rect 152462 0 152518 800
rect 153934 0 153990 800
rect 155498 0 155554 800
rect 156970 0 157026 800
rect 158442 0 158498 800
rect 159914 0 159970 800
rect 161386 0 161442 800
rect 162858 0 162914 800
rect 164422 0 164478 800
rect 165894 0 165950 800
rect 167366 0 167422 800
rect 168838 0 168894 800
rect 170310 0 170366 800
rect 171782 0 171838 800
rect 173346 0 173402 800
rect 174818 0 174874 800
rect 176290 0 176346 800
rect 177762 0 177818 800
rect 179234 0 179290 800
<< obsm2 >>
rect 682 119144 1710 119513
rect 1878 119144 2906 119513
rect 3074 119144 4194 119513
rect 4362 119144 5390 119513
rect 5558 119144 6678 119513
rect 6846 119144 7874 119513
rect 8042 119144 9070 119513
rect 9238 119144 10358 119513
rect 10526 119144 11554 119513
rect 11722 119144 12842 119513
rect 13010 119144 14038 119513
rect 14206 119144 15234 119513
rect 15402 119144 16522 119513
rect 16690 119144 17718 119513
rect 17886 119144 19006 119513
rect 19174 119144 20202 119513
rect 20370 119144 21398 119513
rect 21566 119144 22686 119513
rect 22854 119144 23882 119513
rect 24050 119144 25170 119513
rect 25338 119144 26366 119513
rect 26534 119144 27562 119513
rect 27730 119144 28850 119513
rect 29018 119144 30046 119513
rect 30214 119144 31334 119513
rect 31502 119144 32530 119513
rect 32698 119144 33726 119513
rect 33894 119144 35014 119513
rect 35182 119144 36210 119513
rect 36378 119144 37498 119513
rect 37666 119144 38694 119513
rect 38862 119144 39890 119513
rect 40058 119144 41178 119513
rect 41346 119144 42374 119513
rect 42542 119144 43662 119513
rect 43830 119144 44858 119513
rect 45026 119144 46054 119513
rect 46222 119144 47342 119513
rect 47510 119144 48538 119513
rect 48706 119144 49826 119513
rect 49994 119144 51022 119513
rect 51190 119144 52218 119513
rect 52386 119144 53506 119513
rect 53674 119144 54702 119513
rect 54870 119144 55990 119513
rect 56158 119144 57186 119513
rect 57354 119144 58382 119513
rect 58550 119144 59670 119513
rect 59838 119144 60866 119513
rect 61034 119144 62154 119513
rect 62322 119144 63350 119513
rect 63518 119144 64638 119513
rect 64806 119144 65834 119513
rect 66002 119144 67030 119513
rect 67198 119144 68318 119513
rect 68486 119144 69514 119513
rect 69682 119144 70802 119513
rect 70970 119144 71998 119513
rect 72166 119144 73194 119513
rect 73362 119144 74482 119513
rect 74650 119144 75678 119513
rect 75846 119144 76966 119513
rect 77134 119144 78162 119513
rect 78330 119144 79358 119513
rect 79526 119144 80646 119513
rect 80814 119144 81842 119513
rect 82010 119144 83130 119513
rect 83298 119144 84326 119513
rect 84494 119144 85522 119513
rect 85690 119144 86810 119513
rect 86978 119144 88006 119513
rect 88174 119144 89294 119513
rect 89462 119144 90490 119513
rect 90658 119144 91686 119513
rect 91854 119144 92974 119513
rect 93142 119144 94170 119513
rect 94338 119144 95458 119513
rect 95626 119144 96654 119513
rect 96822 119144 97850 119513
rect 98018 119144 99138 119513
rect 99306 119144 100334 119513
rect 100502 119144 101622 119513
rect 101790 119144 102818 119513
rect 102986 119144 104014 119513
rect 104182 119144 105302 119513
rect 105470 119144 106498 119513
rect 106666 119144 107786 119513
rect 107954 119144 108982 119513
rect 109150 119144 110178 119513
rect 110346 119144 111466 119513
rect 111634 119144 112662 119513
rect 112830 119144 113950 119513
rect 114118 119144 115146 119513
rect 115314 119144 116342 119513
rect 116510 119144 117630 119513
rect 117798 119144 118826 119513
rect 118994 119144 120114 119513
rect 120282 119144 121310 119513
rect 121478 119144 122598 119513
rect 122766 119144 123794 119513
rect 123962 119144 124990 119513
rect 125158 119144 126278 119513
rect 126446 119144 127474 119513
rect 127642 119144 128762 119513
rect 128930 119144 129958 119513
rect 130126 119144 131154 119513
rect 131322 119144 132442 119513
rect 132610 119144 133638 119513
rect 133806 119144 134926 119513
rect 135094 119144 136122 119513
rect 136290 119144 137318 119513
rect 137486 119144 138606 119513
rect 138774 119144 139802 119513
rect 139970 119144 141090 119513
rect 141258 119144 142286 119513
rect 142454 119144 143482 119513
rect 143650 119144 144770 119513
rect 144938 119144 145966 119513
rect 146134 119144 147254 119513
rect 147422 119144 148450 119513
rect 148618 119144 149646 119513
rect 149814 119144 150934 119513
rect 151102 119144 152130 119513
rect 152298 119144 153418 119513
rect 153586 119144 154614 119513
rect 154782 119144 155810 119513
rect 155978 119144 157098 119513
rect 157266 119144 158294 119513
rect 158462 119144 159582 119513
rect 159750 119144 160778 119513
rect 160946 119144 161974 119513
rect 162142 119144 163262 119513
rect 163430 119144 164458 119513
rect 164626 119144 165746 119513
rect 165914 119144 166942 119513
rect 167110 119144 168138 119513
rect 168306 119144 169426 119513
rect 169594 119144 170622 119513
rect 170790 119144 171910 119513
rect 172078 119144 173106 119513
rect 173274 119144 174302 119513
rect 174470 119144 175590 119513
rect 175758 119144 176786 119513
rect 176954 119144 178074 119513
rect 178242 119144 179270 119513
rect 572 856 179380 119144
rect 572 303 698 856
rect 866 303 2170 856
rect 2338 303 3642 856
rect 3810 303 5114 856
rect 5282 303 6586 856
rect 6754 303 8058 856
rect 8226 303 9622 856
rect 9790 303 11094 856
rect 11262 303 12566 856
rect 12734 303 14038 856
rect 14206 303 15510 856
rect 15678 303 16982 856
rect 17150 303 18546 856
rect 18714 303 20018 856
rect 20186 303 21490 856
rect 21658 303 22962 856
rect 23130 303 24434 856
rect 24602 303 25906 856
rect 26074 303 27470 856
rect 27638 303 28942 856
rect 29110 303 30414 856
rect 30582 303 31886 856
rect 32054 303 33358 856
rect 33526 303 34830 856
rect 34998 303 36394 856
rect 36562 303 37866 856
rect 38034 303 39338 856
rect 39506 303 40810 856
rect 40978 303 42282 856
rect 42450 303 43846 856
rect 44014 303 45318 856
rect 45486 303 46790 856
rect 46958 303 48262 856
rect 48430 303 49734 856
rect 49902 303 51206 856
rect 51374 303 52770 856
rect 52938 303 54242 856
rect 54410 303 55714 856
rect 55882 303 57186 856
rect 57354 303 58658 856
rect 58826 303 60130 856
rect 60298 303 61694 856
rect 61862 303 63166 856
rect 63334 303 64638 856
rect 64806 303 66110 856
rect 66278 303 67582 856
rect 67750 303 69054 856
rect 69222 303 70618 856
rect 70786 303 72090 856
rect 72258 303 73562 856
rect 73730 303 75034 856
rect 75202 303 76506 856
rect 76674 303 78070 856
rect 78238 303 79542 856
rect 79710 303 81014 856
rect 81182 303 82486 856
rect 82654 303 83958 856
rect 84126 303 85430 856
rect 85598 303 86994 856
rect 87162 303 88466 856
rect 88634 303 89938 856
rect 90106 303 91410 856
rect 91578 303 92882 856
rect 93050 303 94354 856
rect 94522 303 95918 856
rect 96086 303 97390 856
rect 97558 303 98862 856
rect 99030 303 100334 856
rect 100502 303 101806 856
rect 101974 303 103278 856
rect 103446 303 104842 856
rect 105010 303 106314 856
rect 106482 303 107786 856
rect 107954 303 109258 856
rect 109426 303 110730 856
rect 110898 303 112294 856
rect 112462 303 113766 856
rect 113934 303 115238 856
rect 115406 303 116710 856
rect 116878 303 118182 856
rect 118350 303 119654 856
rect 119822 303 121218 856
rect 121386 303 122690 856
rect 122858 303 124162 856
rect 124330 303 125634 856
rect 125802 303 127106 856
rect 127274 303 128578 856
rect 128746 303 130142 856
rect 130310 303 131614 856
rect 131782 303 133086 856
rect 133254 303 134558 856
rect 134726 303 136030 856
rect 136198 303 137502 856
rect 137670 303 139066 856
rect 139234 303 140538 856
rect 140706 303 142010 856
rect 142178 303 143482 856
rect 143650 303 144954 856
rect 145122 303 146518 856
rect 146686 303 147990 856
rect 148158 303 149462 856
rect 149630 303 150934 856
rect 151102 303 152406 856
rect 152574 303 153878 856
rect 154046 303 155442 856
rect 155610 303 156914 856
rect 157082 303 158386 856
rect 158554 303 159858 856
rect 160026 303 161330 856
rect 161498 303 162802 856
rect 162970 303 164366 856
rect 164534 303 165838 856
rect 166006 303 167310 856
rect 167478 303 168782 856
rect 168950 303 170254 856
rect 170422 303 171726 856
rect 171894 303 173290 856
rect 173458 303 174762 856
rect 174930 303 176234 856
rect 176402 303 177706 856
rect 177874 303 179178 856
rect 179346 303 179380 856
<< metal3 >>
rect 179200 119416 180000 119536
rect 0 118872 800 118992
rect 179200 118736 180000 118856
rect 179200 117920 180000 118040
rect 179200 117240 180000 117360
rect 0 116832 800 116952
rect 179200 116560 180000 116680
rect 179200 115744 180000 115864
rect 179200 115064 180000 115184
rect 0 114792 800 114912
rect 179200 114384 180000 114504
rect 179200 113568 180000 113688
rect 0 112888 800 113008
rect 179200 112888 180000 113008
rect 179200 112208 180000 112328
rect 179200 111392 180000 111512
rect 0 110848 800 110968
rect 179200 110712 180000 110832
rect 179200 110032 180000 110152
rect 179200 109216 180000 109336
rect 0 108808 800 108928
rect 179200 108536 180000 108656
rect 179200 107856 180000 107976
rect 0 106904 800 107024
rect 179200 107040 180000 107160
rect 179200 106360 180000 106480
rect 179200 105680 180000 105800
rect 0 104864 800 104984
rect 179200 104864 180000 104984
rect 179200 104184 180000 104304
rect 179200 103504 180000 103624
rect 0 102824 800 102944
rect 179200 102688 180000 102808
rect 179200 102008 180000 102128
rect 179200 101328 180000 101448
rect 0 100920 800 101040
rect 179200 100512 180000 100632
rect 179200 99832 180000 99952
rect 0 98880 800 99000
rect 179200 99016 180000 99136
rect 179200 98336 180000 98456
rect 179200 97656 180000 97776
rect 0 96840 800 96960
rect 179200 96840 180000 96960
rect 179200 96160 180000 96280
rect 179200 95480 180000 95600
rect 0 94800 800 94920
rect 179200 94664 180000 94784
rect 179200 93984 180000 94104
rect 179200 93304 180000 93424
rect 0 92896 800 93016
rect 179200 92488 180000 92608
rect 179200 91808 180000 91928
rect 179200 91128 180000 91248
rect 0 90856 800 90976
rect 179200 90312 180000 90432
rect 179200 89632 180000 89752
rect 0 88816 800 88936
rect 179200 88952 180000 89072
rect 179200 88136 180000 88256
rect 179200 87456 180000 87576
rect 0 86912 800 87032
rect 179200 86776 180000 86896
rect 179200 85960 180000 86080
rect 179200 85280 180000 85400
rect 0 84872 800 84992
rect 179200 84600 180000 84720
rect 179200 83784 180000 83904
rect 179200 83104 180000 83224
rect 0 82832 800 82952
rect 179200 82424 180000 82544
rect 179200 81608 180000 81728
rect 0 80928 800 81048
rect 179200 80928 180000 81048
rect 179200 80248 180000 80368
rect 179200 79432 180000 79552
rect 0 78888 800 79008
rect 179200 78752 180000 78872
rect 179200 77936 180000 78056
rect 179200 77256 180000 77376
rect 0 76848 800 76968
rect 179200 76576 180000 76696
rect 179200 75760 180000 75880
rect 179200 75080 180000 75200
rect 0 74808 800 74928
rect 179200 74400 180000 74520
rect 179200 73584 180000 73704
rect 0 72904 800 73024
rect 179200 72904 180000 73024
rect 179200 72224 180000 72344
rect 179200 71408 180000 71528
rect 0 70864 800 70984
rect 179200 70728 180000 70848
rect 179200 70048 180000 70168
rect 179200 69232 180000 69352
rect 0 68824 800 68944
rect 179200 68552 180000 68672
rect 179200 67872 180000 67992
rect 0 66920 800 67040
rect 179200 67056 180000 67176
rect 179200 66376 180000 66496
rect 179200 65696 180000 65816
rect 0 64880 800 65000
rect 179200 64880 180000 65000
rect 179200 64200 180000 64320
rect 179200 63520 180000 63640
rect 0 62840 800 62960
rect 179200 62704 180000 62824
rect 179200 62024 180000 62144
rect 179200 61344 180000 61464
rect 0 60936 800 61056
rect 179200 60528 180000 60648
rect 179200 59848 180000 59968
rect 0 58896 800 59016
rect 179200 59032 180000 59152
rect 179200 58352 180000 58472
rect 179200 57672 180000 57792
rect 0 56856 800 56976
rect 179200 56856 180000 56976
rect 179200 56176 180000 56296
rect 179200 55496 180000 55616
rect 0 54816 800 54936
rect 179200 54680 180000 54800
rect 179200 54000 180000 54120
rect 179200 53320 180000 53440
rect 0 52912 800 53032
rect 179200 52504 180000 52624
rect 179200 51824 180000 51944
rect 179200 51144 180000 51264
rect 0 50872 800 50992
rect 179200 50328 180000 50448
rect 179200 49648 180000 49768
rect 0 48832 800 48952
rect 179200 48968 180000 49088
rect 179200 48152 180000 48272
rect 179200 47472 180000 47592
rect 0 46928 800 47048
rect 179200 46792 180000 46912
rect 179200 45976 180000 46096
rect 179200 45296 180000 45416
rect 0 44888 800 45008
rect 179200 44616 180000 44736
rect 179200 43800 180000 43920
rect 179200 43120 180000 43240
rect 0 42848 800 42968
rect 179200 42440 180000 42560
rect 179200 41624 180000 41744
rect 0 40944 800 41064
rect 179200 40944 180000 41064
rect 179200 40264 180000 40384
rect 179200 39448 180000 39568
rect 0 38904 800 39024
rect 179200 38768 180000 38888
rect 179200 37952 180000 38072
rect 179200 37272 180000 37392
rect 0 36864 800 36984
rect 179200 36592 180000 36712
rect 179200 35776 180000 35896
rect 179200 35096 180000 35216
rect 0 34824 800 34944
rect 179200 34416 180000 34536
rect 179200 33600 180000 33720
rect 0 32920 800 33040
rect 179200 32920 180000 33040
rect 179200 32240 180000 32360
rect 179200 31424 180000 31544
rect 0 30880 800 31000
rect 179200 30744 180000 30864
rect 179200 30064 180000 30184
rect 179200 29248 180000 29368
rect 0 28840 800 28960
rect 179200 28568 180000 28688
rect 179200 27888 180000 28008
rect 0 26936 800 27056
rect 179200 27072 180000 27192
rect 179200 26392 180000 26512
rect 179200 25712 180000 25832
rect 0 24896 800 25016
rect 179200 24896 180000 25016
rect 179200 24216 180000 24336
rect 179200 23536 180000 23656
rect 0 22856 800 22976
rect 179200 22720 180000 22840
rect 179200 22040 180000 22160
rect 179200 21360 180000 21480
rect 0 20952 800 21072
rect 179200 20544 180000 20664
rect 179200 19864 180000 19984
rect 0 18912 800 19032
rect 179200 19048 180000 19168
rect 179200 18368 180000 18488
rect 179200 17688 180000 17808
rect 0 16872 800 16992
rect 179200 16872 180000 16992
rect 179200 16192 180000 16312
rect 179200 15512 180000 15632
rect 0 14832 800 14952
rect 179200 14696 180000 14816
rect 179200 14016 180000 14136
rect 179200 13336 180000 13456
rect 0 12928 800 13048
rect 179200 12520 180000 12640
rect 179200 11840 180000 11960
rect 179200 11160 180000 11280
rect 0 10888 800 11008
rect 179200 10344 180000 10464
rect 179200 9664 180000 9784
rect 0 8848 800 8968
rect 179200 8984 180000 9104
rect 179200 8168 180000 8288
rect 179200 7488 180000 7608
rect 0 6944 800 7064
rect 179200 6808 180000 6928
rect 179200 5992 180000 6112
rect 179200 5312 180000 5432
rect 0 4904 800 5024
rect 179200 4632 180000 4752
rect 179200 3816 180000 3936
rect 179200 3136 180000 3256
rect 0 2864 800 2984
rect 179200 2456 180000 2576
rect 179200 1640 180000 1760
rect 0 960 800 1080
rect 179200 960 180000 1080
rect 179200 280 180000 400
<< obsm3 >>
rect 800 119336 179120 119509
rect 800 119072 179200 119336
rect 880 118936 179200 119072
rect 880 118792 179120 118936
rect 800 118656 179120 118792
rect 800 118120 179200 118656
rect 800 117840 179120 118120
rect 800 117440 179200 117840
rect 800 117160 179120 117440
rect 800 117032 179200 117160
rect 880 116760 179200 117032
rect 880 116752 179120 116760
rect 800 116480 179120 116752
rect 800 115944 179200 116480
rect 800 115664 179120 115944
rect 800 115264 179200 115664
rect 800 114992 179120 115264
rect 880 114984 179120 114992
rect 880 114712 179200 114984
rect 800 114584 179200 114712
rect 800 114304 179120 114584
rect 800 113768 179200 114304
rect 800 113488 179120 113768
rect 800 113088 179200 113488
rect 880 112808 179120 113088
rect 800 112408 179200 112808
rect 800 112128 179120 112408
rect 800 111592 179200 112128
rect 800 111312 179120 111592
rect 800 111048 179200 111312
rect 880 110912 179200 111048
rect 880 110768 179120 110912
rect 800 110632 179120 110768
rect 800 110232 179200 110632
rect 800 109952 179120 110232
rect 800 109416 179200 109952
rect 800 109136 179120 109416
rect 800 109008 179200 109136
rect 880 108736 179200 109008
rect 880 108728 179120 108736
rect 800 108456 179120 108728
rect 800 108056 179200 108456
rect 800 107776 179120 108056
rect 800 107240 179200 107776
rect 800 107104 179120 107240
rect 880 106960 179120 107104
rect 880 106824 179200 106960
rect 800 106560 179200 106824
rect 800 106280 179120 106560
rect 800 105880 179200 106280
rect 800 105600 179120 105880
rect 800 105064 179200 105600
rect 880 104784 179120 105064
rect 800 104384 179200 104784
rect 800 104104 179120 104384
rect 800 103704 179200 104104
rect 800 103424 179120 103704
rect 800 103024 179200 103424
rect 880 102888 179200 103024
rect 880 102744 179120 102888
rect 800 102608 179120 102744
rect 800 102208 179200 102608
rect 800 101928 179120 102208
rect 800 101528 179200 101928
rect 800 101248 179120 101528
rect 800 101120 179200 101248
rect 880 100840 179200 101120
rect 800 100712 179200 100840
rect 800 100432 179120 100712
rect 800 100032 179200 100432
rect 800 99752 179120 100032
rect 800 99216 179200 99752
rect 800 99080 179120 99216
rect 880 98936 179120 99080
rect 880 98800 179200 98936
rect 800 98536 179200 98800
rect 800 98256 179120 98536
rect 800 97856 179200 98256
rect 800 97576 179120 97856
rect 800 97040 179200 97576
rect 880 96760 179120 97040
rect 800 96360 179200 96760
rect 800 96080 179120 96360
rect 800 95680 179200 96080
rect 800 95400 179120 95680
rect 800 95000 179200 95400
rect 880 94864 179200 95000
rect 880 94720 179120 94864
rect 800 94584 179120 94720
rect 800 94184 179200 94584
rect 800 93904 179120 94184
rect 800 93504 179200 93904
rect 800 93224 179120 93504
rect 800 93096 179200 93224
rect 880 92816 179200 93096
rect 800 92688 179200 92816
rect 800 92408 179120 92688
rect 800 92008 179200 92408
rect 800 91728 179120 92008
rect 800 91328 179200 91728
rect 800 91056 179120 91328
rect 880 91048 179120 91056
rect 880 90776 179200 91048
rect 800 90512 179200 90776
rect 800 90232 179120 90512
rect 800 89832 179200 90232
rect 800 89552 179120 89832
rect 800 89152 179200 89552
rect 800 89016 179120 89152
rect 880 88872 179120 89016
rect 880 88736 179200 88872
rect 800 88336 179200 88736
rect 800 88056 179120 88336
rect 800 87656 179200 88056
rect 800 87376 179120 87656
rect 800 87112 179200 87376
rect 880 86976 179200 87112
rect 880 86832 179120 86976
rect 800 86696 179120 86832
rect 800 86160 179200 86696
rect 800 85880 179120 86160
rect 800 85480 179200 85880
rect 800 85200 179120 85480
rect 800 85072 179200 85200
rect 880 84800 179200 85072
rect 880 84792 179120 84800
rect 800 84520 179120 84792
rect 800 83984 179200 84520
rect 800 83704 179120 83984
rect 800 83304 179200 83704
rect 800 83032 179120 83304
rect 880 83024 179120 83032
rect 880 82752 179200 83024
rect 800 82624 179200 82752
rect 800 82344 179120 82624
rect 800 81808 179200 82344
rect 800 81528 179120 81808
rect 800 81128 179200 81528
rect 880 80848 179120 81128
rect 800 80448 179200 80848
rect 800 80168 179120 80448
rect 800 79632 179200 80168
rect 800 79352 179120 79632
rect 800 79088 179200 79352
rect 880 78952 179200 79088
rect 880 78808 179120 78952
rect 800 78672 179120 78808
rect 800 78136 179200 78672
rect 800 77856 179120 78136
rect 800 77456 179200 77856
rect 800 77176 179120 77456
rect 800 77048 179200 77176
rect 880 76776 179200 77048
rect 880 76768 179120 76776
rect 800 76496 179120 76768
rect 800 75960 179200 76496
rect 800 75680 179120 75960
rect 800 75280 179200 75680
rect 800 75008 179120 75280
rect 880 75000 179120 75008
rect 880 74728 179200 75000
rect 800 74600 179200 74728
rect 800 74320 179120 74600
rect 800 73784 179200 74320
rect 800 73504 179120 73784
rect 800 73104 179200 73504
rect 880 72824 179120 73104
rect 800 72424 179200 72824
rect 800 72144 179120 72424
rect 800 71608 179200 72144
rect 800 71328 179120 71608
rect 800 71064 179200 71328
rect 880 70928 179200 71064
rect 880 70784 179120 70928
rect 800 70648 179120 70784
rect 800 70248 179200 70648
rect 800 69968 179120 70248
rect 800 69432 179200 69968
rect 800 69152 179120 69432
rect 800 69024 179200 69152
rect 880 68752 179200 69024
rect 880 68744 179120 68752
rect 800 68472 179120 68744
rect 800 68072 179200 68472
rect 800 67792 179120 68072
rect 800 67256 179200 67792
rect 800 67120 179120 67256
rect 880 66976 179120 67120
rect 880 66840 179200 66976
rect 800 66576 179200 66840
rect 800 66296 179120 66576
rect 800 65896 179200 66296
rect 800 65616 179120 65896
rect 800 65080 179200 65616
rect 880 64800 179120 65080
rect 800 64400 179200 64800
rect 800 64120 179120 64400
rect 800 63720 179200 64120
rect 800 63440 179120 63720
rect 800 63040 179200 63440
rect 880 62904 179200 63040
rect 880 62760 179120 62904
rect 800 62624 179120 62760
rect 800 62224 179200 62624
rect 800 61944 179120 62224
rect 800 61544 179200 61944
rect 800 61264 179120 61544
rect 800 61136 179200 61264
rect 880 60856 179200 61136
rect 800 60728 179200 60856
rect 800 60448 179120 60728
rect 800 60048 179200 60448
rect 800 59768 179120 60048
rect 800 59232 179200 59768
rect 800 59096 179120 59232
rect 880 58952 179120 59096
rect 880 58816 179200 58952
rect 800 58552 179200 58816
rect 800 58272 179120 58552
rect 800 57872 179200 58272
rect 800 57592 179120 57872
rect 800 57056 179200 57592
rect 880 56776 179120 57056
rect 800 56376 179200 56776
rect 800 56096 179120 56376
rect 800 55696 179200 56096
rect 800 55416 179120 55696
rect 800 55016 179200 55416
rect 880 54880 179200 55016
rect 880 54736 179120 54880
rect 800 54600 179120 54736
rect 800 54200 179200 54600
rect 800 53920 179120 54200
rect 800 53520 179200 53920
rect 800 53240 179120 53520
rect 800 53112 179200 53240
rect 880 52832 179200 53112
rect 800 52704 179200 52832
rect 800 52424 179120 52704
rect 800 52024 179200 52424
rect 800 51744 179120 52024
rect 800 51344 179200 51744
rect 800 51072 179120 51344
rect 880 51064 179120 51072
rect 880 50792 179200 51064
rect 800 50528 179200 50792
rect 800 50248 179120 50528
rect 800 49848 179200 50248
rect 800 49568 179120 49848
rect 800 49168 179200 49568
rect 800 49032 179120 49168
rect 880 48888 179120 49032
rect 880 48752 179200 48888
rect 800 48352 179200 48752
rect 800 48072 179120 48352
rect 800 47672 179200 48072
rect 800 47392 179120 47672
rect 800 47128 179200 47392
rect 880 46992 179200 47128
rect 880 46848 179120 46992
rect 800 46712 179120 46848
rect 800 46176 179200 46712
rect 800 45896 179120 46176
rect 800 45496 179200 45896
rect 800 45216 179120 45496
rect 800 45088 179200 45216
rect 880 44816 179200 45088
rect 880 44808 179120 44816
rect 800 44536 179120 44808
rect 800 44000 179200 44536
rect 800 43720 179120 44000
rect 800 43320 179200 43720
rect 800 43048 179120 43320
rect 880 43040 179120 43048
rect 880 42768 179200 43040
rect 800 42640 179200 42768
rect 800 42360 179120 42640
rect 800 41824 179200 42360
rect 800 41544 179120 41824
rect 800 41144 179200 41544
rect 880 40864 179120 41144
rect 800 40464 179200 40864
rect 800 40184 179120 40464
rect 800 39648 179200 40184
rect 800 39368 179120 39648
rect 800 39104 179200 39368
rect 880 38968 179200 39104
rect 880 38824 179120 38968
rect 800 38688 179120 38824
rect 800 38152 179200 38688
rect 800 37872 179120 38152
rect 800 37472 179200 37872
rect 800 37192 179120 37472
rect 800 37064 179200 37192
rect 880 36792 179200 37064
rect 880 36784 179120 36792
rect 800 36512 179120 36784
rect 800 35976 179200 36512
rect 800 35696 179120 35976
rect 800 35296 179200 35696
rect 800 35024 179120 35296
rect 880 35016 179120 35024
rect 880 34744 179200 35016
rect 800 34616 179200 34744
rect 800 34336 179120 34616
rect 800 33800 179200 34336
rect 800 33520 179120 33800
rect 800 33120 179200 33520
rect 880 32840 179120 33120
rect 800 32440 179200 32840
rect 800 32160 179120 32440
rect 800 31624 179200 32160
rect 800 31344 179120 31624
rect 800 31080 179200 31344
rect 880 30944 179200 31080
rect 880 30800 179120 30944
rect 800 30664 179120 30800
rect 800 30264 179200 30664
rect 800 29984 179120 30264
rect 800 29448 179200 29984
rect 800 29168 179120 29448
rect 800 29040 179200 29168
rect 880 28768 179200 29040
rect 880 28760 179120 28768
rect 800 28488 179120 28760
rect 800 28088 179200 28488
rect 800 27808 179120 28088
rect 800 27272 179200 27808
rect 800 27136 179120 27272
rect 880 26992 179120 27136
rect 880 26856 179200 26992
rect 800 26592 179200 26856
rect 800 26312 179120 26592
rect 800 25912 179200 26312
rect 800 25632 179120 25912
rect 800 25096 179200 25632
rect 880 24816 179120 25096
rect 800 24416 179200 24816
rect 800 24136 179120 24416
rect 800 23736 179200 24136
rect 800 23456 179120 23736
rect 800 23056 179200 23456
rect 880 22920 179200 23056
rect 880 22776 179120 22920
rect 800 22640 179120 22776
rect 800 22240 179200 22640
rect 800 21960 179120 22240
rect 800 21560 179200 21960
rect 800 21280 179120 21560
rect 800 21152 179200 21280
rect 880 20872 179200 21152
rect 800 20744 179200 20872
rect 800 20464 179120 20744
rect 800 20064 179200 20464
rect 800 19784 179120 20064
rect 800 19248 179200 19784
rect 800 19112 179120 19248
rect 880 18968 179120 19112
rect 880 18832 179200 18968
rect 800 18568 179200 18832
rect 800 18288 179120 18568
rect 800 17888 179200 18288
rect 800 17608 179120 17888
rect 800 17072 179200 17608
rect 880 16792 179120 17072
rect 800 16392 179200 16792
rect 800 16112 179120 16392
rect 800 15712 179200 16112
rect 800 15432 179120 15712
rect 800 15032 179200 15432
rect 880 14896 179200 15032
rect 880 14752 179120 14896
rect 800 14616 179120 14752
rect 800 14216 179200 14616
rect 800 13936 179120 14216
rect 800 13536 179200 13936
rect 800 13256 179120 13536
rect 800 13128 179200 13256
rect 880 12848 179200 13128
rect 800 12720 179200 12848
rect 800 12440 179120 12720
rect 800 12040 179200 12440
rect 800 11760 179120 12040
rect 800 11360 179200 11760
rect 800 11088 179120 11360
rect 880 11080 179120 11088
rect 880 10808 179200 11080
rect 800 10544 179200 10808
rect 800 10264 179120 10544
rect 800 9864 179200 10264
rect 800 9584 179120 9864
rect 800 9184 179200 9584
rect 800 9048 179120 9184
rect 880 8904 179120 9048
rect 880 8768 179200 8904
rect 800 8368 179200 8768
rect 800 8088 179120 8368
rect 800 7688 179200 8088
rect 800 7408 179120 7688
rect 800 7144 179200 7408
rect 880 7008 179200 7144
rect 880 6864 179120 7008
rect 800 6728 179120 6864
rect 800 6192 179200 6728
rect 800 5912 179120 6192
rect 800 5512 179200 5912
rect 800 5232 179120 5512
rect 800 5104 179200 5232
rect 880 4832 179200 5104
rect 880 4824 179120 4832
rect 800 4552 179120 4824
rect 800 4016 179200 4552
rect 800 3736 179120 4016
rect 800 3336 179200 3736
rect 800 3064 179120 3336
rect 880 3056 179120 3064
rect 880 2784 179200 3056
rect 800 2656 179200 2784
rect 800 2376 179120 2656
rect 800 1840 179200 2376
rect 800 1560 179120 1840
rect 800 1160 179200 1560
rect 880 880 179120 1160
rect 800 480 179200 880
rect 800 307 179120 480
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< labels >>
rlabel metal2 s 160834 119200 160890 120000 6 adc0_dat_i[0]
port 1 nsew signal input
rlabel metal3 s 179200 112208 180000 112328 6 adc0_dat_i[10]
port 2 nsew signal input
rlabel metal2 s 170310 0 170366 800 6 adc0_dat_i[11]
port 3 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 adc0_dat_i[12]
port 4 nsew signal input
rlabel metal3 s 0 94800 800 94920 6 adc0_dat_i[13]
port 5 nsew signal input
rlabel metal3 s 0 96840 800 96960 6 adc0_dat_i[14]
port 6 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 adc0_dat_i[15]
port 7 nsew signal input
rlabel metal2 s 168194 119200 168250 120000 6 adc0_dat_i[16]
port 8 nsew signal input
rlabel metal2 s 169482 119200 169538 120000 6 adc0_dat_i[17]
port 9 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 adc0_dat_i[18]
port 10 nsew signal input
rlabel metal3 s 179200 113568 180000 113688 6 adc0_dat_i[19]
port 11 nsew signal input
rlabel metal3 s 179200 110032 180000 110152 6 adc0_dat_i[1]
port 12 nsew signal input
rlabel metal3 s 0 104864 800 104984 6 adc0_dat_i[20]
port 13 nsew signal input
rlabel metal3 s 179200 114384 180000 114504 6 adc0_dat_i[21]
port 14 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 adc0_dat_i[22]
port 15 nsew signal input
rlabel metal2 s 176290 0 176346 800 6 adc0_dat_i[23]
port 16 nsew signal input
rlabel metal2 s 177762 0 177818 800 6 adc0_dat_i[24]
port 17 nsew signal input
rlabel metal2 s 175646 119200 175702 120000 6 adc0_dat_i[25]
port 18 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 adc0_dat_i[26]
port 19 nsew signal input
rlabel metal3 s 179200 117240 180000 117360 6 adc0_dat_i[27]
port 20 nsew signal input
rlabel metal2 s 178130 119200 178186 120000 6 adc0_dat_i[28]
port 21 nsew signal input
rlabel metal3 s 0 116832 800 116952 6 adc0_dat_i[29]
port 22 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 adc0_dat_i[2]
port 23 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 adc0_dat_i[30]
port 24 nsew signal input
rlabel metal3 s 179200 118736 180000 118856 6 adc0_dat_i[31]
port 25 nsew signal input
rlabel metal2 s 162858 0 162914 800 6 adc0_dat_i[3]
port 26 nsew signal input
rlabel metal3 s 0 76848 800 76968 6 adc0_dat_i[4]
port 27 nsew signal input
rlabel metal3 s 179200 111392 180000 111512 6 adc0_dat_i[5]
port 28 nsew signal input
rlabel metal2 s 167366 0 167422 800 6 adc0_dat_i[6]
port 29 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 adc0_dat_i[7]
port 30 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 adc0_dat_i[8]
port 31 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 adc0_dat_i[9]
port 32 nsew signal input
rlabel metal3 s 179200 109216 180000 109336 6 adc1_dat_i[0]
port 33 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 adc1_dat_i[10]
port 34 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 adc1_dat_i[11]
port 35 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 adc1_dat_i[12]
port 36 nsew signal input
rlabel metal3 s 179200 112888 180000 113008 6 adc1_dat_i[13]
port 37 nsew signal input
rlabel metal3 s 0 98880 800 99000 6 adc1_dat_i[14]
port 38 nsew signal input
rlabel metal2 s 173346 0 173402 800 6 adc1_dat_i[15]
port 39 nsew signal input
rlabel metal2 s 174818 0 174874 800 6 adc1_dat_i[16]
port 40 nsew signal input
rlabel metal2 s 170678 119200 170734 120000 6 adc1_dat_i[17]
port 41 nsew signal input
rlabel metal2 s 171966 119200 172022 120000 6 adc1_dat_i[18]
port 42 nsew signal input
rlabel metal2 s 173162 119200 173218 120000 6 adc1_dat_i[19]
port 43 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 adc1_dat_i[1]
port 44 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 adc1_dat_i[20]
port 45 nsew signal input
rlabel metal2 s 174358 119200 174414 120000 6 adc1_dat_i[21]
port 46 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 adc1_dat_i[22]
port 47 nsew signal input
rlabel metal3 s 179200 115064 180000 115184 6 adc1_dat_i[23]
port 48 nsew signal input
rlabel metal3 s 179200 115744 180000 115864 6 adc1_dat_i[24]
port 49 nsew signal input
rlabel metal3 s 179200 116560 180000 116680 6 adc1_dat_i[25]
port 50 nsew signal input
rlabel metal2 s 179234 0 179290 800 6 adc1_dat_i[26]
port 51 nsew signal input
rlabel metal2 s 176842 119200 176898 120000 6 adc1_dat_i[27]
port 52 nsew signal input
rlabel metal3 s 0 114792 800 114912 6 adc1_dat_i[28]
port 53 nsew signal input
rlabel metal2 s 179326 119200 179382 120000 6 adc1_dat_i[29]
port 54 nsew signal input
rlabel metal3 s 179200 110712 180000 110832 6 adc1_dat_i[2]
port 55 nsew signal input
rlabel metal3 s 179200 117920 180000 118040 6 adc1_dat_i[30]
port 56 nsew signal input
rlabel metal3 s 179200 119416 180000 119536 6 adc1_dat_i[31]
port 57 nsew signal input
rlabel metal2 s 164514 119200 164570 120000 6 adc1_dat_i[3]
port 58 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 adc1_dat_i[4]
port 59 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 adc1_dat_i[5]
port 60 nsew signal input
rlabel metal2 s 165802 119200 165858 120000 6 adc1_dat_i[6]
port 61 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 adc1_dat_i[7]
port 62 nsew signal input
rlabel metal2 s 168838 0 168894 800 6 adc1_dat_i[8]
port 63 nsew signal input
rlabel metal2 s 166998 119200 167054 120000 6 adc1_dat_i[9]
port 64 nsew signal input
rlabel metal3 s 0 960 800 1080 6 adc2_dat_i[0]
port 65 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 adc2_dat_i[10]
port 66 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 adc2_dat_i[11]
port 67 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 adc2_dat_i[12]
port 68 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 adc2_dat_i[13]
port 69 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 adc2_dat_i[14]
port 70 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 adc2_dat_i[15]
port 71 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 adc2_dat_i[16]
port 72 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 adc2_dat_i[17]
port 73 nsew signal input
rlabel metal3 s 0 36864 800 36984 6 adc2_dat_i[18]
port 74 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 adc2_dat_i[19]
port 75 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 adc2_dat_i[1]
port 76 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 adc2_dat_i[20]
port 77 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 adc2_dat_i[21]
port 78 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 adc2_dat_i[22]
port 79 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 adc2_dat_i[23]
port 80 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 adc2_dat_i[24]
port 81 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 adc2_dat_i[25]
port 82 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 adc2_dat_i[26]
port 83 nsew signal input
rlabel metal3 s 0 54816 800 54936 6 adc2_dat_i[27]
port 84 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 adc2_dat_i[28]
port 85 nsew signal input
rlabel metal3 s 0 58896 800 59016 6 adc2_dat_i[29]
port 86 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 adc2_dat_i[2]
port 87 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 adc2_dat_i[30]
port 88 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 adc2_dat_i[31]
port 89 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 adc2_dat_i[3]
port 90 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 adc2_dat_i[4]
port 91 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 adc2_dat_i[5]
port 92 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 adc2_dat_i[6]
port 93 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 adc2_dat_i[7]
port 94 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 adc2_dat_i[8]
port 95 nsew signal input
rlabel metal3 s 0 18912 800 19032 6 adc2_dat_i[9]
port 96 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 adc_dvalid_i[0]
port 97 nsew signal input
rlabel metal2 s 159914 0 159970 800 6 adc_dvalid_i[1]
port 98 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 adc_dvalid_i[2]
port 99 nsew signal input
rlabel metal2 s 570 119200 626 120000 6 io_in[0]
port 100 nsew signal input
rlabel metal2 s 37554 119200 37610 120000 6 io_in[10]
port 101 nsew signal input
rlabel metal2 s 41234 119200 41290 120000 6 io_in[11]
port 102 nsew signal input
rlabel metal2 s 44914 119200 44970 120000 6 io_in[12]
port 103 nsew signal input
rlabel metal2 s 48594 119200 48650 120000 6 io_in[13]
port 104 nsew signal input
rlabel metal2 s 52274 119200 52330 120000 6 io_in[14]
port 105 nsew signal input
rlabel metal2 s 56046 119200 56102 120000 6 io_in[15]
port 106 nsew signal input
rlabel metal2 s 59726 119200 59782 120000 6 io_in[16]
port 107 nsew signal input
rlabel metal2 s 63406 119200 63462 120000 6 io_in[17]
port 108 nsew signal input
rlabel metal2 s 67086 119200 67142 120000 6 io_in[18]
port 109 nsew signal input
rlabel metal2 s 70858 119200 70914 120000 6 io_in[19]
port 110 nsew signal input
rlabel metal2 s 4250 119200 4306 120000 6 io_in[1]
port 111 nsew signal input
rlabel metal2 s 74538 119200 74594 120000 6 io_in[20]
port 112 nsew signal input
rlabel metal2 s 78218 119200 78274 120000 6 io_in[21]
port 113 nsew signal input
rlabel metal2 s 81898 119200 81954 120000 6 io_in[22]
port 114 nsew signal input
rlabel metal2 s 85578 119200 85634 120000 6 io_in[23]
port 115 nsew signal input
rlabel metal2 s 89350 119200 89406 120000 6 io_in[24]
port 116 nsew signal input
rlabel metal2 s 93030 119200 93086 120000 6 io_in[25]
port 117 nsew signal input
rlabel metal2 s 96710 119200 96766 120000 6 io_in[26]
port 118 nsew signal input
rlabel metal2 s 100390 119200 100446 120000 6 io_in[27]
port 119 nsew signal input
rlabel metal2 s 104070 119200 104126 120000 6 io_in[28]
port 120 nsew signal input
rlabel metal2 s 107842 119200 107898 120000 6 io_in[29]
port 121 nsew signal input
rlabel metal2 s 7930 119200 7986 120000 6 io_in[2]
port 122 nsew signal input
rlabel metal2 s 111522 119200 111578 120000 6 io_in[30]
port 123 nsew signal input
rlabel metal2 s 115202 119200 115258 120000 6 io_in[31]
port 124 nsew signal input
rlabel metal2 s 118882 119200 118938 120000 6 io_in[32]
port 125 nsew signal input
rlabel metal2 s 122654 119200 122710 120000 6 io_in[33]
port 126 nsew signal input
rlabel metal2 s 126334 119200 126390 120000 6 io_in[34]
port 127 nsew signal input
rlabel metal2 s 130014 119200 130070 120000 6 io_in[35]
port 128 nsew signal input
rlabel metal2 s 133694 119200 133750 120000 6 io_in[36]
port 129 nsew signal input
rlabel metal2 s 137374 119200 137430 120000 6 io_in[37]
port 130 nsew signal input
rlabel metal2 s 11610 119200 11666 120000 6 io_in[3]
port 131 nsew signal input
rlabel metal2 s 15290 119200 15346 120000 6 io_in[4]
port 132 nsew signal input
rlabel metal2 s 19062 119200 19118 120000 6 io_in[5]
port 133 nsew signal input
rlabel metal2 s 22742 119200 22798 120000 6 io_in[6]
port 134 nsew signal input
rlabel metal2 s 26422 119200 26478 120000 6 io_in[7]
port 135 nsew signal input
rlabel metal2 s 30102 119200 30158 120000 6 io_in[8]
port 136 nsew signal input
rlabel metal2 s 33782 119200 33838 120000 6 io_in[9]
port 137 nsew signal input
rlabel metal2 s 1766 119200 1822 120000 6 io_oeb[0]
port 138 nsew signal output
rlabel metal2 s 38750 119200 38806 120000 6 io_oeb[10]
port 139 nsew signal output
rlabel metal2 s 42430 119200 42486 120000 6 io_oeb[11]
port 140 nsew signal output
rlabel metal2 s 46110 119200 46166 120000 6 io_oeb[12]
port 141 nsew signal output
rlabel metal2 s 49882 119200 49938 120000 6 io_oeb[13]
port 142 nsew signal output
rlabel metal2 s 53562 119200 53618 120000 6 io_oeb[14]
port 143 nsew signal output
rlabel metal2 s 57242 119200 57298 120000 6 io_oeb[15]
port 144 nsew signal output
rlabel metal2 s 60922 119200 60978 120000 6 io_oeb[16]
port 145 nsew signal output
rlabel metal2 s 64694 119200 64750 120000 6 io_oeb[17]
port 146 nsew signal output
rlabel metal2 s 68374 119200 68430 120000 6 io_oeb[18]
port 147 nsew signal output
rlabel metal2 s 72054 119200 72110 120000 6 io_oeb[19]
port 148 nsew signal output
rlabel metal2 s 5446 119200 5502 120000 6 io_oeb[1]
port 149 nsew signal output
rlabel metal2 s 75734 119200 75790 120000 6 io_oeb[20]
port 150 nsew signal output
rlabel metal2 s 79414 119200 79470 120000 6 io_oeb[21]
port 151 nsew signal output
rlabel metal2 s 83186 119200 83242 120000 6 io_oeb[22]
port 152 nsew signal output
rlabel metal2 s 86866 119200 86922 120000 6 io_oeb[23]
port 153 nsew signal output
rlabel metal2 s 90546 119200 90602 120000 6 io_oeb[24]
port 154 nsew signal output
rlabel metal2 s 94226 119200 94282 120000 6 io_oeb[25]
port 155 nsew signal output
rlabel metal2 s 97906 119200 97962 120000 6 io_oeb[26]
port 156 nsew signal output
rlabel metal2 s 101678 119200 101734 120000 6 io_oeb[27]
port 157 nsew signal output
rlabel metal2 s 105358 119200 105414 120000 6 io_oeb[28]
port 158 nsew signal output
rlabel metal2 s 109038 119200 109094 120000 6 io_oeb[29]
port 159 nsew signal output
rlabel metal2 s 9126 119200 9182 120000 6 io_oeb[2]
port 160 nsew signal output
rlabel metal2 s 112718 119200 112774 120000 6 io_oeb[30]
port 161 nsew signal output
rlabel metal2 s 116398 119200 116454 120000 6 io_oeb[31]
port 162 nsew signal output
rlabel metal2 s 120170 119200 120226 120000 6 io_oeb[32]
port 163 nsew signal output
rlabel metal2 s 123850 119200 123906 120000 6 io_oeb[33]
port 164 nsew signal output
rlabel metal2 s 127530 119200 127586 120000 6 io_oeb[34]
port 165 nsew signal output
rlabel metal2 s 131210 119200 131266 120000 6 io_oeb[35]
port 166 nsew signal output
rlabel metal2 s 134982 119200 135038 120000 6 io_oeb[36]
port 167 nsew signal output
rlabel metal2 s 138662 119200 138718 120000 6 io_oeb[37]
port 168 nsew signal output
rlabel metal2 s 12898 119200 12954 120000 6 io_oeb[3]
port 169 nsew signal output
rlabel metal2 s 16578 119200 16634 120000 6 io_oeb[4]
port 170 nsew signal output
rlabel metal2 s 20258 119200 20314 120000 6 io_oeb[5]
port 171 nsew signal output
rlabel metal2 s 23938 119200 23994 120000 6 io_oeb[6]
port 172 nsew signal output
rlabel metal2 s 27618 119200 27674 120000 6 io_oeb[7]
port 173 nsew signal output
rlabel metal2 s 31390 119200 31446 120000 6 io_oeb[8]
port 174 nsew signal output
rlabel metal2 s 35070 119200 35126 120000 6 io_oeb[9]
port 175 nsew signal output
rlabel metal2 s 2962 119200 3018 120000 6 io_out[0]
port 176 nsew signal output
rlabel metal2 s 39946 119200 40002 120000 6 io_out[10]
port 177 nsew signal output
rlabel metal2 s 43718 119200 43774 120000 6 io_out[11]
port 178 nsew signal output
rlabel metal2 s 47398 119200 47454 120000 6 io_out[12]
port 179 nsew signal output
rlabel metal2 s 51078 119200 51134 120000 6 io_out[13]
port 180 nsew signal output
rlabel metal2 s 54758 119200 54814 120000 6 io_out[14]
port 181 nsew signal output
rlabel metal2 s 58438 119200 58494 120000 6 io_out[15]
port 182 nsew signal output
rlabel metal2 s 62210 119200 62266 120000 6 io_out[16]
port 183 nsew signal output
rlabel metal2 s 65890 119200 65946 120000 6 io_out[17]
port 184 nsew signal output
rlabel metal2 s 69570 119200 69626 120000 6 io_out[18]
port 185 nsew signal output
rlabel metal2 s 73250 119200 73306 120000 6 io_out[19]
port 186 nsew signal output
rlabel metal2 s 6734 119200 6790 120000 6 io_out[1]
port 187 nsew signal output
rlabel metal2 s 77022 119200 77078 120000 6 io_out[20]
port 188 nsew signal output
rlabel metal2 s 80702 119200 80758 120000 6 io_out[21]
port 189 nsew signal output
rlabel metal2 s 84382 119200 84438 120000 6 io_out[22]
port 190 nsew signal output
rlabel metal2 s 88062 119200 88118 120000 6 io_out[23]
port 191 nsew signal output
rlabel metal2 s 91742 119200 91798 120000 6 io_out[24]
port 192 nsew signal output
rlabel metal2 s 95514 119200 95570 120000 6 io_out[25]
port 193 nsew signal output
rlabel metal2 s 99194 119200 99250 120000 6 io_out[26]
port 194 nsew signal output
rlabel metal2 s 102874 119200 102930 120000 6 io_out[27]
port 195 nsew signal output
rlabel metal2 s 106554 119200 106610 120000 6 io_out[28]
port 196 nsew signal output
rlabel metal2 s 110234 119200 110290 120000 6 io_out[29]
port 197 nsew signal output
rlabel metal2 s 10414 119200 10470 120000 6 io_out[2]
port 198 nsew signal output
rlabel metal2 s 114006 119200 114062 120000 6 io_out[30]
port 199 nsew signal output
rlabel metal2 s 117686 119200 117742 120000 6 io_out[31]
port 200 nsew signal output
rlabel metal2 s 121366 119200 121422 120000 6 io_out[32]
port 201 nsew signal output
rlabel metal2 s 125046 119200 125102 120000 6 io_out[33]
port 202 nsew signal output
rlabel metal2 s 128818 119200 128874 120000 6 io_out[34]
port 203 nsew signal output
rlabel metal2 s 132498 119200 132554 120000 6 io_out[35]
port 204 nsew signal output
rlabel metal2 s 136178 119200 136234 120000 6 io_out[36]
port 205 nsew signal output
rlabel metal2 s 139858 119200 139914 120000 6 io_out[37]
port 206 nsew signal output
rlabel metal2 s 14094 119200 14150 120000 6 io_out[3]
port 207 nsew signal output
rlabel metal2 s 17774 119200 17830 120000 6 io_out[4]
port 208 nsew signal output
rlabel metal2 s 21454 119200 21510 120000 6 io_out[5]
port 209 nsew signal output
rlabel metal2 s 25226 119200 25282 120000 6 io_out[6]
port 210 nsew signal output
rlabel metal2 s 28906 119200 28962 120000 6 io_out[7]
port 211 nsew signal output
rlabel metal2 s 32586 119200 32642 120000 6 io_out[8]
port 212 nsew signal output
rlabel metal2 s 36266 119200 36322 120000 6 io_out[9]
port 213 nsew signal output
rlabel metal2 s 162030 119200 162086 120000 6 irq[0]
port 214 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 irq[1]
port 215 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 irq[2]
port 216 nsew signal output
rlabel metal3 s 179200 280 180000 400 6 mem1_data_i[0]
port 217 nsew signal input
rlabel metal3 s 179200 45296 180000 45416 6 mem1_data_i[10]
port 218 nsew signal input
rlabel metal3 s 179200 48152 180000 48272 6 mem1_data_i[11]
port 219 nsew signal input
rlabel metal3 s 179200 51144 180000 51264 6 mem1_data_i[12]
port 220 nsew signal input
rlabel metal3 s 179200 54000 180000 54120 6 mem1_data_i[13]
port 221 nsew signal input
rlabel metal3 s 179200 56856 180000 56976 6 mem1_data_i[14]
port 222 nsew signal input
rlabel metal3 s 179200 59848 180000 59968 6 mem1_data_i[15]
port 223 nsew signal input
rlabel metal3 s 179200 62704 180000 62824 6 mem1_data_i[16]
port 224 nsew signal input
rlabel metal3 s 179200 65696 180000 65816 6 mem1_data_i[17]
port 225 nsew signal input
rlabel metal3 s 179200 68552 180000 68672 6 mem1_data_i[18]
port 226 nsew signal input
rlabel metal3 s 179200 71408 180000 71528 6 mem1_data_i[19]
port 227 nsew signal input
rlabel metal3 s 179200 5992 180000 6112 6 mem1_data_i[1]
port 228 nsew signal input
rlabel metal3 s 179200 74400 180000 74520 6 mem1_data_i[20]
port 229 nsew signal input
rlabel metal3 s 179200 77256 180000 77376 6 mem1_data_i[21]
port 230 nsew signal input
rlabel metal3 s 179200 80248 180000 80368 6 mem1_data_i[22]
port 231 nsew signal input
rlabel metal3 s 179200 83104 180000 83224 6 mem1_data_i[23]
port 232 nsew signal input
rlabel metal3 s 179200 85960 180000 86080 6 mem1_data_i[24]
port 233 nsew signal input
rlabel metal3 s 179200 88952 180000 89072 6 mem1_data_i[25]
port 234 nsew signal input
rlabel metal3 s 179200 91808 180000 91928 6 mem1_data_i[26]
port 235 nsew signal input
rlabel metal3 s 179200 94664 180000 94784 6 mem1_data_i[27]
port 236 nsew signal input
rlabel metal3 s 179200 97656 180000 97776 6 mem1_data_i[28]
port 237 nsew signal input
rlabel metal3 s 179200 100512 180000 100632 6 mem1_data_i[29]
port 238 nsew signal input
rlabel metal3 s 179200 11840 180000 11960 6 mem1_data_i[2]
port 239 nsew signal input
rlabel metal3 s 179200 103504 180000 103624 6 mem1_data_i[30]
port 240 nsew signal input
rlabel metal3 s 179200 106360 180000 106480 6 mem1_data_i[31]
port 241 nsew signal input
rlabel metal3 s 179200 16192 180000 16312 6 mem1_data_i[3]
port 242 nsew signal input
rlabel metal3 s 179200 20544 180000 20664 6 mem1_data_i[4]
port 243 nsew signal input
rlabel metal3 s 179200 24896 180000 25016 6 mem1_data_i[5]
port 244 nsew signal input
rlabel metal3 s 179200 29248 180000 29368 6 mem1_data_i[6]
port 245 nsew signal input
rlabel metal3 s 179200 33600 180000 33720 6 mem1_data_i[7]
port 246 nsew signal input
rlabel metal3 s 179200 37952 180000 38072 6 mem1_data_i[8]
port 247 nsew signal input
rlabel metal3 s 179200 42440 180000 42560 6 mem1_data_i[9]
port 248 nsew signal input
rlabel metal3 s 179200 960 180000 1080 6 mem_data2_i[0]
port 249 nsew signal input
rlabel metal3 s 179200 45976 180000 46096 6 mem_data2_i[10]
port 250 nsew signal input
rlabel metal3 s 179200 48968 180000 49088 6 mem_data2_i[11]
port 251 nsew signal input
rlabel metal3 s 179200 51824 180000 51944 6 mem_data2_i[12]
port 252 nsew signal input
rlabel metal3 s 179200 54680 180000 54800 6 mem_data2_i[13]
port 253 nsew signal input
rlabel metal3 s 179200 57672 180000 57792 6 mem_data2_i[14]
port 254 nsew signal input
rlabel metal3 s 179200 60528 180000 60648 6 mem_data2_i[15]
port 255 nsew signal input
rlabel metal3 s 179200 63520 180000 63640 6 mem_data2_i[16]
port 256 nsew signal input
rlabel metal3 s 179200 66376 180000 66496 6 mem_data2_i[17]
port 257 nsew signal input
rlabel metal3 s 179200 69232 180000 69352 6 mem_data2_i[18]
port 258 nsew signal input
rlabel metal3 s 179200 72224 180000 72344 6 mem_data2_i[19]
port 259 nsew signal input
rlabel metal3 s 179200 6808 180000 6928 6 mem_data2_i[1]
port 260 nsew signal input
rlabel metal3 s 179200 75080 180000 75200 6 mem_data2_i[20]
port 261 nsew signal input
rlabel metal3 s 179200 77936 180000 78056 6 mem_data2_i[21]
port 262 nsew signal input
rlabel metal3 s 179200 80928 180000 81048 6 mem_data2_i[22]
port 263 nsew signal input
rlabel metal3 s 179200 83784 180000 83904 6 mem_data2_i[23]
port 264 nsew signal input
rlabel metal3 s 179200 86776 180000 86896 6 mem_data2_i[24]
port 265 nsew signal input
rlabel metal3 s 179200 89632 180000 89752 6 mem_data2_i[25]
port 266 nsew signal input
rlabel metal3 s 179200 92488 180000 92608 6 mem_data2_i[26]
port 267 nsew signal input
rlabel metal3 s 179200 95480 180000 95600 6 mem_data2_i[27]
port 268 nsew signal input
rlabel metal3 s 179200 98336 180000 98456 6 mem_data2_i[28]
port 269 nsew signal input
rlabel metal3 s 179200 101328 180000 101448 6 mem_data2_i[29]
port 270 nsew signal input
rlabel metal3 s 179200 12520 180000 12640 6 mem_data2_i[2]
port 271 nsew signal input
rlabel metal3 s 179200 104184 180000 104304 6 mem_data2_i[30]
port 272 nsew signal input
rlabel metal3 s 179200 107040 180000 107160 6 mem_data2_i[31]
port 273 nsew signal input
rlabel metal3 s 179200 16872 180000 16992 6 mem_data2_i[3]
port 274 nsew signal input
rlabel metal3 s 179200 21360 180000 21480 6 mem_data2_i[4]
port 275 nsew signal input
rlabel metal3 s 179200 25712 180000 25832 6 mem_data2_i[5]
port 276 nsew signal input
rlabel metal3 s 179200 30064 180000 30184 6 mem_data2_i[6]
port 277 nsew signal input
rlabel metal3 s 179200 34416 180000 34536 6 mem_data2_i[7]
port 278 nsew signal input
rlabel metal3 s 179200 38768 180000 38888 6 mem_data2_i[8]
port 279 nsew signal input
rlabel metal3 s 179200 43120 180000 43240 6 mem_data2_i[9]
port 280 nsew signal input
rlabel metal3 s 179200 1640 180000 1760 6 mem_data_i[0]
port 281 nsew signal input
rlabel metal3 s 179200 46792 180000 46912 6 mem_data_i[10]
port 282 nsew signal input
rlabel metal3 s 179200 49648 180000 49768 6 mem_data_i[11]
port 283 nsew signal input
rlabel metal3 s 179200 52504 180000 52624 6 mem_data_i[12]
port 284 nsew signal input
rlabel metal3 s 179200 55496 180000 55616 6 mem_data_i[13]
port 285 nsew signal input
rlabel metal3 s 179200 58352 180000 58472 6 mem_data_i[14]
port 286 nsew signal input
rlabel metal3 s 179200 61344 180000 61464 6 mem_data_i[15]
port 287 nsew signal input
rlabel metal3 s 179200 64200 180000 64320 6 mem_data_i[16]
port 288 nsew signal input
rlabel metal3 s 179200 67056 180000 67176 6 mem_data_i[17]
port 289 nsew signal input
rlabel metal3 s 179200 70048 180000 70168 6 mem_data_i[18]
port 290 nsew signal input
rlabel metal3 s 179200 72904 180000 73024 6 mem_data_i[19]
port 291 nsew signal input
rlabel metal3 s 179200 7488 180000 7608 6 mem_data_i[1]
port 292 nsew signal input
rlabel metal3 s 179200 75760 180000 75880 6 mem_data_i[20]
port 293 nsew signal input
rlabel metal3 s 179200 78752 180000 78872 6 mem_data_i[21]
port 294 nsew signal input
rlabel metal3 s 179200 81608 180000 81728 6 mem_data_i[22]
port 295 nsew signal input
rlabel metal3 s 179200 84600 180000 84720 6 mem_data_i[23]
port 296 nsew signal input
rlabel metal3 s 179200 87456 180000 87576 6 mem_data_i[24]
port 297 nsew signal input
rlabel metal3 s 179200 90312 180000 90432 6 mem_data_i[25]
port 298 nsew signal input
rlabel metal3 s 179200 93304 180000 93424 6 mem_data_i[26]
port 299 nsew signal input
rlabel metal3 s 179200 96160 180000 96280 6 mem_data_i[27]
port 300 nsew signal input
rlabel metal3 s 179200 99016 180000 99136 6 mem_data_i[28]
port 301 nsew signal input
rlabel metal3 s 179200 102008 180000 102128 6 mem_data_i[29]
port 302 nsew signal input
rlabel metal3 s 179200 13336 180000 13456 6 mem_data_i[2]
port 303 nsew signal input
rlabel metal3 s 179200 104864 180000 104984 6 mem_data_i[30]
port 304 nsew signal input
rlabel metal3 s 179200 107856 180000 107976 6 mem_data_i[31]
port 305 nsew signal input
rlabel metal3 s 179200 17688 180000 17808 6 mem_data_i[3]
port 306 nsew signal input
rlabel metal3 s 179200 22040 180000 22160 6 mem_data_i[4]
port 307 nsew signal input
rlabel metal3 s 179200 26392 180000 26512 6 mem_data_i[5]
port 308 nsew signal input
rlabel metal3 s 179200 30744 180000 30864 6 mem_data_i[6]
port 309 nsew signal input
rlabel metal3 s 179200 35096 180000 35216 6 mem_data_i[7]
port 310 nsew signal input
rlabel metal3 s 179200 39448 180000 39568 6 mem_data_i[8]
port 311 nsew signal input
rlabel metal3 s 179200 43800 180000 43920 6 mem_data_i[9]
port 312 nsew signal input
rlabel metal3 s 179200 2456 180000 2576 6 mem_data_o[0]
port 313 nsew signal output
rlabel metal3 s 179200 47472 180000 47592 6 mem_data_o[10]
port 314 nsew signal output
rlabel metal3 s 179200 50328 180000 50448 6 mem_data_o[11]
port 315 nsew signal output
rlabel metal3 s 179200 53320 180000 53440 6 mem_data_o[12]
port 316 nsew signal output
rlabel metal3 s 179200 56176 180000 56296 6 mem_data_o[13]
port 317 nsew signal output
rlabel metal3 s 179200 59032 180000 59152 6 mem_data_o[14]
port 318 nsew signal output
rlabel metal3 s 179200 62024 180000 62144 6 mem_data_o[15]
port 319 nsew signal output
rlabel metal3 s 179200 64880 180000 65000 6 mem_data_o[16]
port 320 nsew signal output
rlabel metal3 s 179200 67872 180000 67992 6 mem_data_o[17]
port 321 nsew signal output
rlabel metal3 s 179200 70728 180000 70848 6 mem_data_o[18]
port 322 nsew signal output
rlabel metal3 s 179200 73584 180000 73704 6 mem_data_o[19]
port 323 nsew signal output
rlabel metal3 s 179200 8168 180000 8288 6 mem_data_o[1]
port 324 nsew signal output
rlabel metal3 s 179200 76576 180000 76696 6 mem_data_o[20]
port 325 nsew signal output
rlabel metal3 s 179200 79432 180000 79552 6 mem_data_o[21]
port 326 nsew signal output
rlabel metal3 s 179200 82424 180000 82544 6 mem_data_o[22]
port 327 nsew signal output
rlabel metal3 s 179200 85280 180000 85400 6 mem_data_o[23]
port 328 nsew signal output
rlabel metal3 s 179200 88136 180000 88256 6 mem_data_o[24]
port 329 nsew signal output
rlabel metal3 s 179200 91128 180000 91248 6 mem_data_o[25]
port 330 nsew signal output
rlabel metal3 s 179200 93984 180000 94104 6 mem_data_o[26]
port 331 nsew signal output
rlabel metal3 s 179200 96840 180000 96960 6 mem_data_o[27]
port 332 nsew signal output
rlabel metal3 s 179200 99832 180000 99952 6 mem_data_o[28]
port 333 nsew signal output
rlabel metal3 s 179200 102688 180000 102808 6 mem_data_o[29]
port 334 nsew signal output
rlabel metal3 s 179200 14016 180000 14136 6 mem_data_o[2]
port 335 nsew signal output
rlabel metal3 s 179200 105680 180000 105800 6 mem_data_o[30]
port 336 nsew signal output
rlabel metal3 s 179200 108536 180000 108656 6 mem_data_o[31]
port 337 nsew signal output
rlabel metal3 s 179200 18368 180000 18488 6 mem_data_o[3]
port 338 nsew signal output
rlabel metal3 s 179200 22720 180000 22840 6 mem_data_o[4]
port 339 nsew signal output
rlabel metal3 s 179200 27072 180000 27192 6 mem_data_o[5]
port 340 nsew signal output
rlabel metal3 s 179200 31424 180000 31544 6 mem_data_o[6]
port 341 nsew signal output
rlabel metal3 s 179200 35776 180000 35896 6 mem_data_o[7]
port 342 nsew signal output
rlabel metal3 s 179200 40264 180000 40384 6 mem_data_o[8]
port 343 nsew signal output
rlabel metal3 s 179200 44616 180000 44736 6 mem_data_o[9]
port 344 nsew signal output
rlabel metal3 s 179200 3136 180000 3256 6 mem_raddr_o[0]
port 345 nsew signal output
rlabel metal3 s 179200 8984 180000 9104 6 mem_raddr_o[1]
port 346 nsew signal output
rlabel metal3 s 179200 14696 180000 14816 6 mem_raddr_o[2]
port 347 nsew signal output
rlabel metal3 s 179200 19048 180000 19168 6 mem_raddr_o[3]
port 348 nsew signal output
rlabel metal3 s 179200 23536 180000 23656 6 mem_raddr_o[4]
port 349 nsew signal output
rlabel metal3 s 179200 27888 180000 28008 6 mem_raddr_o[5]
port 350 nsew signal output
rlabel metal3 s 179200 32240 180000 32360 6 mem_raddr_o[6]
port 351 nsew signal output
rlabel metal3 s 179200 36592 180000 36712 6 mem_raddr_o[7]
port 352 nsew signal output
rlabel metal3 s 179200 40944 180000 41064 6 mem_raddr_o[8]
port 353 nsew signal output
rlabel metal3 s 179200 3816 180000 3936 6 mem_renb_o[0]
port 354 nsew signal output
rlabel metal3 s 179200 9664 180000 9784 6 mem_renb_o[1]
port 355 nsew signal output
rlabel metal3 s 179200 4632 180000 4752 6 mem_waddr_o[0]
port 356 nsew signal output
rlabel metal3 s 179200 10344 180000 10464 6 mem_waddr_o[1]
port 357 nsew signal output
rlabel metal3 s 179200 15512 180000 15632 6 mem_waddr_o[2]
port 358 nsew signal output
rlabel metal3 s 179200 19864 180000 19984 6 mem_waddr_o[3]
port 359 nsew signal output
rlabel metal3 s 179200 24216 180000 24336 6 mem_waddr_o[4]
port 360 nsew signal output
rlabel metal3 s 179200 28568 180000 28688 6 mem_waddr_o[5]
port 361 nsew signal output
rlabel metal3 s 179200 32920 180000 33040 6 mem_waddr_o[6]
port 362 nsew signal output
rlabel metal3 s 179200 37272 180000 37392 6 mem_waddr_o[7]
port 363 nsew signal output
rlabel metal3 s 179200 41624 180000 41744 6 mem_waddr_o[8]
port 364 nsew signal output
rlabel metal3 s 179200 5312 180000 5432 6 mem_wenb_o[0]
port 365 nsew signal output
rlabel metal3 s 179200 11160 180000 11280 6 mem_wenb_o[1]
port 366 nsew signal output
rlabel metal2 s 141146 119200 141202 120000 6 oversample_o[0]
port 367 nsew signal output
rlabel metal2 s 142342 119200 142398 120000 6 oversample_o[1]
port 368 nsew signal output
rlabel metal2 s 143538 119200 143594 120000 6 oversample_o[2]
port 369 nsew signal output
rlabel metal2 s 144826 119200 144882 120000 6 oversample_o[3]
port 370 nsew signal output
rlabel metal2 s 146022 119200 146078 120000 6 oversample_o[4]
port 371 nsew signal output
rlabel metal2 s 147310 119200 147366 120000 6 oversample_o[5]
port 372 nsew signal output
rlabel metal2 s 148506 119200 148562 120000 6 oversample_o[6]
port 373 nsew signal output
rlabel metal2 s 149702 119200 149758 120000 6 oversample_o[7]
port 374 nsew signal output
rlabel metal2 s 150990 119200 151046 120000 6 oversample_o[8]
port 375 nsew signal output
rlabel metal2 s 152186 119200 152242 120000 6 oversample_o[9]
port 376 nsew signal output
rlabel metal2 s 157154 119200 157210 120000 6 sinc3_en_o[0]
port 377 nsew signal output
rlabel metal2 s 158350 119200 158406 120000 6 sinc3_en_o[1]
port 378 nsew signal output
rlabel metal2 s 159638 119200 159694 120000 6 sinc3_en_o[2]
port 379 nsew signal output
rlabel metal2 s 153474 119200 153530 120000 6 vco_enb_o[0]
port 380 nsew signal output
rlabel metal2 s 154670 119200 154726 120000 6 vco_enb_o[1]
port 381 nsew signal output
rlabel metal2 s 155866 119200 155922 120000 6 vco_enb_o[2]
port 382 nsew signal output
rlabel metal2 s 754 0 810 800 6 wb_clk_i
port 383 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wb_rst_i
port 384 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_ack_o
port 385 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 wbs_adr_i[0]
port 386 nsew signal input
rlabel metal2 s 60186 0 60242 800 6 wbs_adr_i[10]
port 387 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wbs_adr_i[11]
port 388 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 wbs_adr_i[12]
port 389 nsew signal input
rlabel metal2 s 73618 0 73674 800 6 wbs_adr_i[13]
port 390 nsew signal input
rlabel metal2 s 78126 0 78182 800 6 wbs_adr_i[14]
port 391 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 wbs_adr_i[15]
port 392 nsew signal input
rlabel metal2 s 87050 0 87106 800 6 wbs_adr_i[16]
port 393 nsew signal input
rlabel metal2 s 91466 0 91522 800 6 wbs_adr_i[17]
port 394 nsew signal input
rlabel metal2 s 95974 0 96030 800 6 wbs_adr_i[18]
port 395 nsew signal input
rlabel metal2 s 100390 0 100446 800 6 wbs_adr_i[19]
port 396 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wbs_adr_i[1]
port 397 nsew signal input
rlabel metal2 s 104898 0 104954 800 6 wbs_adr_i[20]
port 398 nsew signal input
rlabel metal2 s 109314 0 109370 800 6 wbs_adr_i[21]
port 399 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 wbs_adr_i[22]
port 400 nsew signal input
rlabel metal2 s 118238 0 118294 800 6 wbs_adr_i[23]
port 401 nsew signal input
rlabel metal2 s 122746 0 122802 800 6 wbs_adr_i[24]
port 402 nsew signal input
rlabel metal2 s 127162 0 127218 800 6 wbs_adr_i[25]
port 403 nsew signal input
rlabel metal2 s 131670 0 131726 800 6 wbs_adr_i[26]
port 404 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 wbs_adr_i[27]
port 405 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 wbs_adr_i[28]
port 406 nsew signal input
rlabel metal2 s 145010 0 145066 800 6 wbs_adr_i[29]
port 407 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 wbs_adr_i[2]
port 408 nsew signal input
rlabel metal2 s 149518 0 149574 800 6 wbs_adr_i[30]
port 409 nsew signal input
rlabel metal2 s 153934 0 153990 800 6 wbs_adr_i[31]
port 410 nsew signal input
rlabel metal2 s 27526 0 27582 800 6 wbs_adr_i[3]
port 411 nsew signal input
rlabel metal2 s 33414 0 33470 800 6 wbs_adr_i[4]
port 412 nsew signal input
rlabel metal2 s 37922 0 37978 800 6 wbs_adr_i[5]
port 413 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 wbs_adr_i[6]
port 414 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_adr_i[7]
port 415 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 wbs_adr_i[8]
port 416 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 wbs_adr_i[9]
port 417 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_cyc_i
port 418 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_i[0]
port 419 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_dat_i[10]
port 420 nsew signal input
rlabel metal2 s 66166 0 66222 800 6 wbs_dat_i[11]
port 421 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 wbs_dat_i[12]
port 422 nsew signal input
rlabel metal2 s 75090 0 75146 800 6 wbs_dat_i[13]
port 423 nsew signal input
rlabel metal2 s 79598 0 79654 800 6 wbs_dat_i[14]
port 424 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_dat_i[15]
port 425 nsew signal input
rlabel metal2 s 88522 0 88578 800 6 wbs_dat_i[16]
port 426 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 wbs_dat_i[17]
port 427 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_dat_i[18]
port 428 nsew signal input
rlabel metal2 s 101862 0 101918 800 6 wbs_dat_i[19]
port 429 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 wbs_dat_i[1]
port 430 nsew signal input
rlabel metal2 s 106370 0 106426 800 6 wbs_dat_i[20]
port 431 nsew signal input
rlabel metal2 s 110786 0 110842 800 6 wbs_dat_i[21]
port 432 nsew signal input
rlabel metal2 s 115294 0 115350 800 6 wbs_dat_i[22]
port 433 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 wbs_dat_i[23]
port 434 nsew signal input
rlabel metal2 s 124218 0 124274 800 6 wbs_dat_i[24]
port 435 nsew signal input
rlabel metal2 s 128634 0 128690 800 6 wbs_dat_i[25]
port 436 nsew signal input
rlabel metal2 s 133142 0 133198 800 6 wbs_dat_i[26]
port 437 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 wbs_dat_i[27]
port 438 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 wbs_dat_i[28]
port 439 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 wbs_dat_i[29]
port 440 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_i[2]
port 441 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 wbs_dat_i[30]
port 442 nsew signal input
rlabel metal2 s 155498 0 155554 800 6 wbs_dat_i[31]
port 443 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 wbs_dat_i[3]
port 444 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wbs_dat_i[4]
port 445 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 wbs_dat_i[5]
port 446 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 wbs_dat_i[6]
port 447 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[7]
port 448 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 wbs_dat_i[8]
port 449 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 wbs_dat_i[9]
port 450 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[0]
port 451 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 wbs_dat_o[10]
port 452 nsew signal output
rlabel metal2 s 67638 0 67694 800 6 wbs_dat_o[11]
port 453 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[12]
port 454 nsew signal output
rlabel metal2 s 76562 0 76618 800 6 wbs_dat_o[13]
port 455 nsew signal output
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_o[14]
port 456 nsew signal output
rlabel metal2 s 85486 0 85542 800 6 wbs_dat_o[15]
port 457 nsew signal output
rlabel metal2 s 89994 0 90050 800 6 wbs_dat_o[16]
port 458 nsew signal output
rlabel metal2 s 94410 0 94466 800 6 wbs_dat_o[17]
port 459 nsew signal output
rlabel metal2 s 98918 0 98974 800 6 wbs_dat_o[18]
port 460 nsew signal output
rlabel metal2 s 103334 0 103390 800 6 wbs_dat_o[19]
port 461 nsew signal output
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_o[1]
port 462 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 wbs_dat_o[20]
port 463 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 wbs_dat_o[21]
port 464 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 wbs_dat_o[22]
port 465 nsew signal output
rlabel metal2 s 121274 0 121330 800 6 wbs_dat_o[23]
port 466 nsew signal output
rlabel metal2 s 125690 0 125746 800 6 wbs_dat_o[24]
port 467 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 wbs_dat_o[25]
port 468 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 wbs_dat_o[26]
port 469 nsew signal output
rlabel metal2 s 139122 0 139178 800 6 wbs_dat_o[27]
port 470 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 wbs_dat_o[28]
port 471 nsew signal output
rlabel metal2 s 148046 0 148102 800 6 wbs_dat_o[29]
port 472 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 wbs_dat_o[2]
port 473 nsew signal output
rlabel metal2 s 152462 0 152518 800 6 wbs_dat_o[30]
port 474 nsew signal output
rlabel metal2 s 156970 0 157026 800 6 wbs_dat_o[31]
port 475 nsew signal output
rlabel metal2 s 30470 0 30526 800 6 wbs_dat_o[3]
port 476 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 wbs_dat_o[4]
port 477 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 wbs_dat_o[5]
port 478 nsew signal output
rlabel metal2 s 45374 0 45430 800 6 wbs_dat_o[6]
port 479 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 wbs_dat_o[7]
port 480 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 wbs_dat_o[8]
port 481 nsew signal output
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_o[9]
port 482 nsew signal output
rlabel metal2 s 14094 0 14150 800 6 wbs_sel_i[0]
port 483 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 wbs_sel_i[1]
port 484 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 wbs_sel_i[2]
port 485 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_sel_i[3]
port 486 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_stb_i
port 487 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_we_i
port 488 nsew signal input
rlabel metal3 s 0 64880 800 65000 6 wmask_o[0]
port 489 nsew signal output
rlabel metal2 s 161386 0 161442 800 6 wmask_o[1]
port 490 nsew signal output
rlabel metal2 s 163318 119200 163374 120000 6 wmask_o[2]
port 491 nsew signal output
rlabel metal2 s 164422 0 164478 800 6 wmask_o[3]
port 492 nsew signal output
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 493 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 494 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 495 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 496 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 497 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 498 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 499 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 500 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 501 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 502 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 503 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 504 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 505 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 506 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 507 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 508 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 509 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 510 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 511 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 512 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 513 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 514 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 515 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 516 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 517 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 518 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 519 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 520 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 521 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 522 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 523 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 524 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 525 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 526 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 527 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 528 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 529 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 530 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 531 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 532 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 533 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 534 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 535 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 536 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 538 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 539 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 540 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 8663362
string GDS_START 689282
<< end >>

