VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_adc_wrapper
  CLASS BLOCK ;
  FOREIGN vco_adc_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 700.000 BY 700.000 ;
  PIN adc0_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 696.000 2.670 700.000 ;
    END
  END adc0_dat_i[0]
  PIN adc0_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 696.000 176.090 700.000 ;
    END
  END adc0_dat_i[10]
  PIN adc0_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 696.000 191.730 700.000 ;
    END
  END adc0_dat_i[11]
  PIN adc0_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 696.000 207.830 700.000 ;
    END
  END adc0_dat_i[12]
  PIN adc0_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.190 696.000 223.470 700.000 ;
    END
  END adc0_dat_i[13]
  PIN adc0_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 696.000 239.110 700.000 ;
    END
  END adc0_dat_i[14]
  PIN adc0_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.930 696.000 255.210 700.000 ;
    END
  END adc0_dat_i[15]
  PIN adc0_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 696.000 270.850 700.000 ;
    END
  END adc0_dat_i[16]
  PIN adc0_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.210 696.000 286.490 700.000 ;
    END
  END adc0_dat_i[17]
  PIN adc0_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.310 696.000 302.590 700.000 ;
    END
  END adc0_dat_i[18]
  PIN adc0_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 696.000 318.230 700.000 ;
    END
  END adc0_dat_i[19]
  PIN adc0_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 696.000 23.370 700.000 ;
    END
  END adc0_dat_i[1]
  PIN adc0_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.590 696.000 333.870 700.000 ;
    END
  END adc0_dat_i[20]
  PIN adc0_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.690 696.000 349.970 700.000 ;
    END
  END adc0_dat_i[21]
  PIN adc0_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.330 696.000 365.610 700.000 ;
    END
  END adc0_dat_i[22]
  PIN adc0_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.970 696.000 381.250 700.000 ;
    END
  END adc0_dat_i[23]
  PIN adc0_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 397.070 696.000 397.350 700.000 ;
    END
  END adc0_dat_i[24]
  PIN adc0_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 696.000 412.990 700.000 ;
    END
  END adc0_dat_i[25]
  PIN adc0_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 696.000 428.630 700.000 ;
    END
  END adc0_dat_i[26]
  PIN adc0_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 696.000 444.730 700.000 ;
    END
  END adc0_dat_i[27]
  PIN adc0_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.090 696.000 460.370 700.000 ;
    END
  END adc0_dat_i[28]
  PIN adc0_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 696.000 476.010 700.000 ;
    END
  END adc0_dat_i[29]
  PIN adc0_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 696.000 44.530 700.000 ;
    END
  END adc0_dat_i[2]
  PIN adc0_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 696.000 492.110 700.000 ;
    END
  END adc0_dat_i[30]
  PIN adc0_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.470 696.000 507.750 700.000 ;
    END
  END adc0_dat_i[31]
  PIN adc0_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 65.410 696.000 65.690 700.000 ;
    END
  END adc0_dat_i[3]
  PIN adc0_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 696.000 81.330 700.000 ;
    END
  END adc0_dat_i[4]
  PIN adc0_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 696.000 96.970 700.000 ;
    END
  END adc0_dat_i[5]
  PIN adc0_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 696.000 113.070 700.000 ;
    END
  END adc0_dat_i[6]
  PIN adc0_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 696.000 128.710 700.000 ;
    END
  END adc0_dat_i[7]
  PIN adc0_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 696.000 144.350 700.000 ;
    END
  END adc0_dat_i[8]
  PIN adc0_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 696.000 160.450 700.000 ;
    END
  END adc0_dat_i[9]
  PIN adc1_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 7.450 696.000 7.730 700.000 ;
    END
  END adc1_dat_i[0]
  PIN adc1_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 696.000 181.610 700.000 ;
    END
  END adc1_dat_i[10]
  PIN adc1_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.970 696.000 197.250 700.000 ;
    END
  END adc1_dat_i[11]
  PIN adc1_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 696.000 212.890 700.000 ;
    END
  END adc1_dat_i[12]
  PIN adc1_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 696.000 228.990 700.000 ;
    END
  END adc1_dat_i[13]
  PIN adc1_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 696.000 244.630 700.000 ;
    END
  END adc1_dat_i[14]
  PIN adc1_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 259.990 696.000 260.270 700.000 ;
    END
  END adc1_dat_i[15]
  PIN adc1_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 696.000 276.370 700.000 ;
    END
  END adc1_dat_i[16]
  PIN adc1_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.730 696.000 292.010 700.000 ;
    END
  END adc1_dat_i[17]
  PIN adc1_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 307.370 696.000 307.650 700.000 ;
    END
  END adc1_dat_i[18]
  PIN adc1_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 696.000 323.750 700.000 ;
    END
  END adc1_dat_i[19]
  PIN adc1_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.610 696.000 28.890 700.000 ;
    END
  END adc1_dat_i[1]
  PIN adc1_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.110 696.000 339.390 700.000 ;
    END
  END adc1_dat_i[20]
  PIN adc1_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.750 696.000 355.030 700.000 ;
    END
  END adc1_dat_i[21]
  PIN adc1_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 696.000 371.130 700.000 ;
    END
  END adc1_dat_i[22]
  PIN adc1_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 696.000 386.770 700.000 ;
    END
  END adc1_dat_i[23]
  PIN adc1_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.130 696.000 402.410 700.000 ;
    END
  END adc1_dat_i[24]
  PIN adc1_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 696.000 418.510 700.000 ;
    END
  END adc1_dat_i[25]
  PIN adc1_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 433.870 696.000 434.150 700.000 ;
    END
  END adc1_dat_i[26]
  PIN adc1_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 449.510 696.000 449.790 700.000 ;
    END
  END adc1_dat_i[27]
  PIN adc1_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 696.000 465.890 700.000 ;
    END
  END adc1_dat_i[28]
  PIN adc1_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.250 696.000 481.530 700.000 ;
    END
  END adc1_dat_i[29]
  PIN adc1_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 696.000 49.590 700.000 ;
    END
  END adc1_dat_i[2]
  PIN adc1_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.890 696.000 497.170 700.000 ;
    END
  END adc1_dat_i[30]
  PIN adc1_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 696.000 513.270 700.000 ;
    END
  END adc1_dat_i[31]
  PIN adc1_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.470 696.000 70.750 700.000 ;
    END
  END adc1_dat_i[3]
  PIN adc1_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 86.570 696.000 86.850 700.000 ;
    END
  END adc1_dat_i[4]
  PIN adc1_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 696.000 102.490 700.000 ;
    END
  END adc1_dat_i[5]
  PIN adc1_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 696.000 118.130 700.000 ;
    END
  END adc1_dat_i[6]
  PIN adc1_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 696.000 134.230 700.000 ;
    END
  END adc1_dat_i[7]
  PIN adc1_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 149.590 696.000 149.870 700.000 ;
    END
  END adc1_dat_i[8]
  PIN adc1_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 696.000 165.510 700.000 ;
    END
  END adc1_dat_i[9]
  PIN adc2_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 696.000 12.790 700.000 ;
    END
  END adc2_dat_i[0]
  PIN adc2_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 696.000 186.670 700.000 ;
    END
  END adc2_dat_i[10]
  PIN adc2_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.030 696.000 202.310 700.000 ;
    END
  END adc2_dat_i[11]
  PIN adc2_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 218.130 696.000 218.410 700.000 ;
    END
  END adc2_dat_i[12]
  PIN adc2_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 696.000 234.050 700.000 ;
    END
  END adc2_dat_i[13]
  PIN adc2_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 249.410 696.000 249.690 700.000 ;
    END
  END adc2_dat_i[14]
  PIN adc2_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 696.000 265.790 700.000 ;
    END
  END adc2_dat_i[15]
  PIN adc2_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 696.000 281.430 700.000 ;
    END
  END adc2_dat_i[16]
  PIN adc2_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.790 696.000 297.070 700.000 ;
    END
  END adc2_dat_i[17]
  PIN adc2_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.890 696.000 313.170 700.000 ;
    END
  END adc2_dat_i[18]
  PIN adc2_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 696.000 328.810 700.000 ;
    END
  END adc2_dat_i[19]
  PIN adc2_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 33.670 696.000 33.950 700.000 ;
    END
  END adc2_dat_i[1]
  PIN adc2_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.170 696.000 344.450 700.000 ;
    END
  END adc2_dat_i[20]
  PIN adc2_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.270 696.000 360.550 700.000 ;
    END
  END adc2_dat_i[21]
  PIN adc2_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 696.000 376.190 700.000 ;
    END
  END adc2_dat_i[22]
  PIN adc2_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.550 696.000 391.830 700.000 ;
    END
  END adc2_dat_i[23]
  PIN adc2_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.650 696.000 407.930 700.000 ;
    END
  END adc2_dat_i[24]
  PIN adc2_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 696.000 423.570 700.000 ;
    END
  END adc2_dat_i[25]
  PIN adc2_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 696.000 439.210 700.000 ;
    END
  END adc2_dat_i[26]
  PIN adc2_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 696.000 455.310 700.000 ;
    END
  END adc2_dat_i[27]
  PIN adc2_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.670 696.000 470.950 700.000 ;
    END
  END adc2_dat_i[28]
  PIN adc2_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 486.310 696.000 486.590 700.000 ;
    END
  END adc2_dat_i[29]
  PIN adc2_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 696.000 55.110 700.000 ;
    END
  END adc2_dat_i[2]
  PIN adc2_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 696.000 502.690 700.000 ;
    END
  END adc2_dat_i[30]
  PIN adc2_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 696.000 518.330 700.000 ;
    END
  END adc2_dat_i[31]
  PIN adc2_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.990 696.000 76.270 700.000 ;
    END
  END adc2_dat_i[3]
  PIN adc2_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.630 696.000 91.910 700.000 ;
    END
  END adc2_dat_i[4]
  PIN adc2_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 696.000 107.550 700.000 ;
    END
  END adc2_dat_i[5]
  PIN adc2_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.370 696.000 123.650 700.000 ;
    END
  END adc2_dat_i[6]
  PIN adc2_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.010 696.000 139.290 700.000 ;
    END
  END adc2_dat_i[7]
  PIN adc2_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 696.000 154.930 700.000 ;
    END
  END adc2_dat_i[8]
  PIN adc2_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 696.000 171.030 700.000 ;
    END
  END adc2_dat_i[9]
  PIN adc_dvalid_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.030 696.000 18.310 700.000 ;
    END
  END adc_dvalid_i[0]
  PIN adc_dvalid_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 696.000 39.470 700.000 ;
    END
  END adc_dvalid_i[1]
  PIN adc_dvalid_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 696.000 60.170 700.000 ;
    END
  END adc_dvalid_i[2]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 34.720 700.000 35.320 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 501.200 700.000 501.800 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 547.440 700.000 548.040 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 594.360 700.000 594.960 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 641.280 700.000 641.880 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 687.520 700.000 688.120 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.990 696.000 697.270 700.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 696.000 686.690 700.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.830 696.000 676.110 700.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 665.250 696.000 665.530 700.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.130 696.000 655.410 700.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 80.960 700.000 81.560 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.550 696.000 644.830 700.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.970 696.000 634.250 700.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.390 696.000 623.670 700.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.810 696.000 613.090 700.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 614.080 4.000 614.680 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 620.200 4.000 620.800 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.000 4.000 627.600 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.920 4.000 640.520 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 127.880 700.000 128.480 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 652.840 4.000 653.440 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 4.000 659.560 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 665.760 4.000 666.360 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 671.880 4.000 672.480 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 678.000 4.000 678.600 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 697.720 4.000 698.320 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 174.800 700.000 175.400 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 221.040 700.000 221.640 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 267.960 700.000 268.560 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 314.200 700.000 314.800 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 361.120 700.000 361.720 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 408.040 700.000 408.640 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 454.280 700.000 454.880 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 11.600 700.000 12.200 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 478.080 700.000 478.680 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 524.320 700.000 524.920 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 571.240 700.000 571.840 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 617.480 700.000 618.080 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 664.400 700.000 665.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 696.000 692.210 700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 696.000 681.630 700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.770 696.000 671.050 700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 660.190 696.000 660.470 700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 696.000 649.890 700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 57.840 700.000 58.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.030 696.000 639.310 700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.450 696.000 628.730 700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.870 696.000 618.150 700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 696.000 608.030 700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 617.480 4.000 618.080 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 630.400 4.000 631.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 636.520 4.000 637.120 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 643.320 4.000 643.920 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 104.760 700.000 105.360 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 649.440 4.000 650.040 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 655.560 4.000 656.160 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 662.360 4.000 662.960 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.280 4.000 675.880 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 681.400 4.000 682.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 688.200 4.000 688.800 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 694.320 4.000 694.920 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 151.000 700.000 151.600 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 197.920 700.000 198.520 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 244.840 700.000 245.440 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 291.080 700.000 291.680 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 338.000 700.000 338.600 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 384.240 700.000 384.840 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 696.000 431.160 700.000 431.760 ;
    END
  END io_out[9]
  PIN mem0_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 199.960 4.000 200.560 ;
    END
  END mem0_data_i[0]
  PIN mem0_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 328.480 4.000 329.080 ;
    END
  END mem0_data_i[10]
  PIN mem0_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 341.400 4.000 342.000 ;
    END
  END mem0_data_i[11]
  PIN mem0_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END mem0_data_i[12]
  PIN mem0_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END mem0_data_i[13]
  PIN mem0_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 379.480 4.000 380.080 ;
    END
  END mem0_data_i[14]
  PIN mem0_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END mem0_data_i[15]
  PIN mem0_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 405.320 4.000 405.920 ;
    END
  END mem0_data_i[16]
  PIN mem0_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END mem0_data_i[17]
  PIN mem0_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.160 4.000 431.760 ;
    END
  END mem0_data_i[18]
  PIN mem0_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END mem0_data_i[19]
  PIN mem0_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.880 4.000 213.480 ;
    END
  END mem0_data_i[1]
  PIN mem0_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.000 4.000 457.600 ;
    END
  END mem0_data_i[20]
  PIN mem0_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END mem0_data_i[21]
  PIN mem0_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END mem0_data_i[22]
  PIN mem0_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.080 4.000 495.680 ;
    END
  END mem0_data_i[23]
  PIN mem0_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END mem0_data_i[24]
  PIN mem0_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 520.920 4.000 521.520 ;
    END
  END mem0_data_i[25]
  PIN mem0_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END mem0_data_i[26]
  PIN mem0_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 546.760 4.000 547.360 ;
    END
  END mem0_data_i[27]
  PIN mem0_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.680 4.000 560.280 ;
    END
  END mem0_data_i[28]
  PIN mem0_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 572.600 4.000 573.200 ;
    END
  END mem0_data_i[29]
  PIN mem0_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END mem0_data_i[2]
  PIN mem0_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 585.520 4.000 586.120 ;
    END
  END mem0_data_i[30]
  PIN mem0_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 597.760 4.000 598.360 ;
    END
  END mem0_data_i[31]
  PIN mem0_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END mem0_data_i[3]
  PIN mem0_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END mem0_data_i[4]
  PIN mem0_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END mem0_data_i[5]
  PIN mem0_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.800 4.000 277.400 ;
    END
  END mem0_data_i[6]
  PIN mem0_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.720 4.000 290.320 ;
    END
  END mem0_data_i[7]
  PIN mem0_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END mem0_data_i[8]
  PIN mem0_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 315.560 4.000 316.160 ;
    END
  END mem0_data_i[9]
  PIN mem1_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END mem1_data_i[0]
  PIN mem1_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END mem1_data_i[10]
  PIN mem1_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 344.800 4.000 345.400 ;
    END
  END mem1_data_i[11]
  PIN mem1_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END mem1_data_i[12]
  PIN mem1_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END mem1_data_i[13]
  PIN mem1_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 382.880 4.000 383.480 ;
    END
  END mem1_data_i[14]
  PIN mem1_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 395.800 4.000 396.400 ;
    END
  END mem1_data_i[15]
  PIN mem1_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END mem1_data_i[16]
  PIN mem1_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END mem1_data_i[17]
  PIN mem1_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END mem1_data_i[18]
  PIN mem1_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 447.480 4.000 448.080 ;
    END
  END mem1_data_i[19]
  PIN mem1_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 216.280 4.000 216.880 ;
    END
  END mem1_data_i[1]
  PIN mem1_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.720 4.000 460.320 ;
    END
  END mem1_data_i[20]
  PIN mem1_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END mem1_data_i[21]
  PIN mem1_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 485.560 4.000 486.160 ;
    END
  END mem1_data_i[22]
  PIN mem1_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 498.480 4.000 499.080 ;
    END
  END mem1_data_i[23]
  PIN mem1_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END mem1_data_i[24]
  PIN mem1_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END mem1_data_i[25]
  PIN mem1_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.240 4.000 537.840 ;
    END
  END mem1_data_i[26]
  PIN mem1_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 550.160 4.000 550.760 ;
    END
  END mem1_data_i[27]
  PIN mem1_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.080 4.000 563.680 ;
    END
  END mem1_data_i[28]
  PIN mem1_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 575.320 4.000 575.920 ;
    END
  END mem1_data_i[29]
  PIN mem1_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 229.200 4.000 229.800 ;
    END
  END mem1_data_i[2]
  PIN mem1_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END mem1_data_i[30]
  PIN mem1_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END mem1_data_i[31]
  PIN mem1_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END mem1_data_i[3]
  PIN mem1_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END mem1_data_i[4]
  PIN mem1_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 267.280 4.000 267.880 ;
    END
  END mem1_data_i[5]
  PIN mem1_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END mem1_data_i[6]
  PIN mem1_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 293.120 4.000 293.720 ;
    END
  END mem1_data_i[7]
  PIN mem1_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END mem1_data_i[8]
  PIN mem1_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.960 4.000 319.560 ;
    END
  END mem1_data_i[9]
  PIN mem2_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END mem2_data_i[0]
  PIN mem2_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 334.600 4.000 335.200 ;
    END
  END mem2_data_i[10]
  PIN mem2_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 347.520 4.000 348.120 ;
    END
  END mem2_data_i[11]
  PIN mem2_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END mem2_data_i[12]
  PIN mem2_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 373.360 4.000 373.960 ;
    END
  END mem2_data_i[13]
  PIN mem2_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END mem2_data_i[14]
  PIN mem2_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END mem2_data_i[15]
  PIN mem2_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.120 4.000 412.720 ;
    END
  END mem2_data_i[16]
  PIN mem2_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END mem2_data_i[17]
  PIN mem2_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END mem2_data_i[18]
  PIN mem2_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.200 4.000 450.800 ;
    END
  END mem2_data_i[19]
  PIN mem2_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.000 4.000 219.600 ;
    END
  END mem2_data_i[1]
  PIN mem2_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END mem2_data_i[20]
  PIN mem2_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END mem2_data_i[21]
  PIN mem2_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END mem2_data_i[22]
  PIN mem2_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.880 4.000 502.480 ;
    END
  END mem2_data_i[23]
  PIN mem2_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 514.800 4.000 515.400 ;
    END
  END mem2_data_i[24]
  PIN mem2_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 527.720 4.000 528.320 ;
    END
  END mem2_data_i[25]
  PIN mem2_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 539.960 4.000 540.560 ;
    END
  END mem2_data_i[26]
  PIN mem2_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END mem2_data_i[27]
  PIN mem2_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 565.800 4.000 566.400 ;
    END
  END mem2_data_i[28]
  PIN mem2_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END mem2_data_i[29]
  PIN mem2_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END mem2_data_i[2]
  PIN mem2_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 591.640 4.000 592.240 ;
    END
  END mem2_data_i[30]
  PIN mem2_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END mem2_data_i[31]
  PIN mem2_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END mem2_data_i[3]
  PIN mem2_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.760 4.000 258.360 ;
    END
  END mem2_data_i[4]
  PIN mem2_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END mem2_data_i[5]
  PIN mem2_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END mem2_data_i[6]
  PIN mem2_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END mem2_data_i[7]
  PIN mem2_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END mem2_data_i[8]
  PIN mem2_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END mem2_data_i[9]
  PIN mem3_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END mem3_data_i[0]
  PIN mem3_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.000 4.000 338.600 ;
    END
  END mem3_data_i[10]
  PIN mem3_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.920 4.000 351.520 ;
    END
  END mem3_data_i[11]
  PIN mem3_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END mem3_data_i[12]
  PIN mem3_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END mem3_data_i[13]
  PIN mem3_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 389.680 4.000 390.280 ;
    END
  END mem3_data_i[14]
  PIN mem3_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 402.600 4.000 403.200 ;
    END
  END mem3_data_i[15]
  PIN mem3_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END mem3_data_i[16]
  PIN mem3_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END mem3_data_i[17]
  PIN mem3_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.680 4.000 441.280 ;
    END
  END mem3_data_i[18]
  PIN mem3_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END mem3_data_i[19]
  PIN mem3_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END mem3_data_i[1]
  PIN mem3_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END mem3_data_i[20]
  PIN mem3_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END mem3_data_i[21]
  PIN mem3_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END mem3_data_i[22]
  PIN mem3_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END mem3_data_i[23]
  PIN mem3_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 517.520 4.000 518.120 ;
    END
  END mem3_data_i[24]
  PIN mem3_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END mem3_data_i[25]
  PIN mem3_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 543.360 4.000 543.960 ;
    END
  END mem3_data_i[26]
  PIN mem3_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END mem3_data_i[27]
  PIN mem3_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 569.200 4.000 569.800 ;
    END
  END mem3_data_i[28]
  PIN mem3_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 582.120 4.000 582.720 ;
    END
  END mem3_data_i[29]
  PIN mem3_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END mem3_data_i[2]
  PIN mem3_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END mem3_data_i[30]
  PIN mem3_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 607.960 4.000 608.560 ;
    END
  END mem3_data_i[31]
  PIN mem3_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END mem3_data_i[3]
  PIN mem3_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.160 4.000 261.760 ;
    END
  END mem3_data_i[4]
  PIN mem3_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 274.080 4.000 274.680 ;
    END
  END mem3_data_i[5]
  PIN mem3_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END mem3_data_i[6]
  PIN mem3_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END mem3_data_i[7]
  PIN mem3_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END mem3_data_i[8]
  PIN mem3_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.080 4.000 325.680 ;
    END
  END mem3_data_i[9]
  PIN mem_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END mem_data_o[0]
  PIN mem_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 116.320 4.000 116.920 ;
    END
  END mem_data_o[10]
  PIN mem_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.720 4.000 120.320 ;
    END
  END mem_data_o[11]
  PIN mem_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END mem_data_o[12]
  PIN mem_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 126.520 4.000 127.120 ;
    END
  END mem_data_o[13]
  PIN mem_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END mem_data_o[14]
  PIN mem_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END mem_data_o[15]
  PIN mem_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END mem_data_o[16]
  PIN mem_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END mem_data_o[17]
  PIN mem_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.160 4.000 142.760 ;
    END
  END mem_data_o[18]
  PIN mem_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END mem_data_o[19]
  PIN mem_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.760 4.000 88.360 ;
    END
  END mem_data_o[1]
  PIN mem_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END mem_data_o[20]
  PIN mem_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END mem_data_o[21]
  PIN mem_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END mem_data_o[22]
  PIN mem_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END mem_data_o[23]
  PIN mem_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 161.880 4.000 162.480 ;
    END
  END mem_data_o[24]
  PIN mem_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END mem_data_o[25]
  PIN mem_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.000 4.000 168.600 ;
    END
  END mem_data_o[26]
  PIN mem_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END mem_data_o[27]
  PIN mem_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END mem_data_o[28]
  PIN mem_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 177.520 4.000 178.120 ;
    END
  END mem_data_o[29]
  PIN mem_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END mem_data_o[2]
  PIN mem_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END mem_data_o[30]
  PIN mem_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 184.320 4.000 184.920 ;
    END
  END mem_data_o[31]
  PIN mem_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END mem_data_o[3]
  PIN mem_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.280 4.000 97.880 ;
    END
  END mem_data_o[4]
  PIN mem_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.680 4.000 101.280 ;
    END
  END mem_data_o[5]
  PIN mem_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.080 4.000 104.680 ;
    END
  END mem_data_o[6]
  PIN mem_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END mem_data_o[7]
  PIN mem_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 110.200 4.000 110.800 ;
    END
  END mem_data_o[8]
  PIN mem_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END mem_data_o[9]
  PIN mem_raddr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 1.400 4.000 2.000 ;
    END
  END mem_raddr_o[0]
  PIN mem_raddr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 4.120 4.000 4.720 ;
    END
  END mem_raddr_o[1]
  PIN mem_raddr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END mem_raddr_o[2]
  PIN mem_raddr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.920 4.000 11.520 ;
    END
  END mem_raddr_o[3]
  PIN mem_raddr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END mem_raddr_o[4]
  PIN mem_raddr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END mem_raddr_o[5]
  PIN mem_raddr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END mem_raddr_o[6]
  PIN mem_raddr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END mem_raddr_o[7]
  PIN mem_raddr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 26.560 4.000 27.160 ;
    END
  END mem_raddr_o[8]
  PIN mem_renb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 58.520 4.000 59.120 ;
    END
  END mem_renb_o[0]
  PIN mem_renb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.920 4.000 62.520 ;
    END
  END mem_renb_o[1]
  PIN mem_renb_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END mem_renb_o[2]
  PIN mem_renb_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.720 4.000 69.320 ;
    END
  END mem_renb_o[3]
  PIN mem_waddr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END mem_waddr_o[0]
  PIN mem_waddr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END mem_waddr_o[1]
  PIN mem_waddr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.080 4.000 36.680 ;
    END
  END mem_waddr_o[2]
  PIN mem_waddr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 39.480 4.000 40.080 ;
    END
  END mem_waddr_o[3]
  PIN mem_waddr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END mem_waddr_o[4]
  PIN mem_waddr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 46.280 4.000 46.880 ;
    END
  END mem_waddr_o[5]
  PIN mem_waddr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END mem_waddr_o[6]
  PIN mem_waddr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END mem_waddr_o[7]
  PIN mem_waddr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.800 4.000 56.400 ;
    END
  END mem_waddr_o[8]
  PIN mem_wenb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END mem_wenb_o[0]
  PIN mem_wenb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END mem_wenb_o[1]
  PIN mem_wenb_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END mem_wenb_o[2]
  PIN mem_wenb_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END mem_wenb_o[3]
  PIN oversample_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.110 696.000 523.390 700.000 ;
    END
  END oversample_o[0]
  PIN oversample_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 696.000 528.910 700.000 ;
    END
  END oversample_o[1]
  PIN oversample_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.690 696.000 533.970 700.000 ;
    END
  END oversample_o[2]
  PIN oversample_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 696.000 539.490 700.000 ;
    END
  END oversample_o[3]
  PIN oversample_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 696.000 544.550 700.000 ;
    END
  END oversample_o[4]
  PIN oversample_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 549.790 696.000 550.070 700.000 ;
    END
  END oversample_o[5]
  PIN oversample_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 554.850 696.000 555.130 700.000 ;
    END
  END oversample_o[6]
  PIN oversample_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 696.000 560.650 700.000 ;
    END
  END oversample_o[7]
  PIN oversample_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 565.430 696.000 565.710 700.000 ;
    END
  END oversample_o[8]
  PIN oversample_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.490 696.000 570.770 700.000 ;
    END
  END oversample_o[9]
  PIN sinc3_en_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 591.650 696.000 591.930 700.000 ;
    END
  END sinc3_en_o[0]
  PIN sinc3_en_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.170 696.000 597.450 700.000 ;
    END
  END sinc3_en_o[1]
  PIN sinc3_en_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.230 696.000 602.510 700.000 ;
    END
  END sinc3_en_o[2]
  PIN vco_enb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 696.000 576.290 700.000 ;
    END
  END vco_enb_o[0]
  PIN vco_enb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 696.000 581.350 700.000 ;
    END
  END vco_enb_o[1]
  PIN vco_enb_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 696.000 586.870 700.000 ;
    END
  END vco_enb_o[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 306.910 0.000 307.190 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 0.000 366.530 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.590 0.000 425.870 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 0.000 465.890 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.730 0.000 545.010 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.290 0.000 584.570 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.070 0.000 604.350 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.630 0.000 643.910 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 0.000 663.690 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.990 0.000 168.270 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.230 0.000 188.510 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.570 0.000 247.850 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 0.000 49.590 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.570 0.000 293.850 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 0.000 333.410 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 373.150 0.000 373.430 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.710 0.000 412.990 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 0.000 432.770 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.270 0.000 452.550 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 75.530 0.000 75.810 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 472.050 0.000 472.330 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 491.830 0.000 492.110 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.610 0.000 511.890 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.390 0.000 531.670 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.170 0.000 551.450 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.950 0.000 571.230 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 0.000 631.030 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.530 0.000 650.810 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.310 0.000 670.590 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.890 0.000 175.170 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 0.000 214.730 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 234.230 0.000 234.510 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 0.000 56.030 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.690 0.000 280.970 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.470 0.000 300.750 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 340.030 0.000 340.310 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 359.810 0.000 360.090 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.590 0.000 379.870 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.150 0.000 419.430 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 458.710 0.000 458.990 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 0.000 82.710 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 478.490 0.000 478.770 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.270 0.000 498.550 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.050 0.000 518.330 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 538.290 0.000 538.570 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 558.070 0.000 558.350 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 577.850 0.000 578.130 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 0.000 597.910 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.410 0.000 617.690 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 637.190 0.000 637.470 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.970 0.000 657.250 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 0.000 696.810 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.330 0.000 181.610 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 201.110 0.000 201.390 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 0.000 115.830 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 4.000 ;
    END
  END wbs_we_i
  PIN wmask_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END wmask_o[0]
  PIN wmask_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END wmask_o[1]
  PIN wmask_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END wmask_o[2]
  PIN wmask_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END wmask_o[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 694.140 688.245 ;
      LAYER met1 ;
        RECT 2.370 9.220 697.290 688.400 ;
      LAYER met2 ;
        RECT 2.950 695.720 7.170 698.205 ;
        RECT 8.010 695.720 12.230 698.205 ;
        RECT 13.070 695.720 17.750 698.205 ;
        RECT 18.590 695.720 22.810 698.205 ;
        RECT 23.650 695.720 28.330 698.205 ;
        RECT 29.170 695.720 33.390 698.205 ;
        RECT 34.230 695.720 38.910 698.205 ;
        RECT 39.750 695.720 43.970 698.205 ;
        RECT 44.810 695.720 49.030 698.205 ;
        RECT 49.870 695.720 54.550 698.205 ;
        RECT 55.390 695.720 59.610 698.205 ;
        RECT 60.450 695.720 65.130 698.205 ;
        RECT 65.970 695.720 70.190 698.205 ;
        RECT 71.030 695.720 75.710 698.205 ;
        RECT 76.550 695.720 80.770 698.205 ;
        RECT 81.610 695.720 86.290 698.205 ;
        RECT 87.130 695.720 91.350 698.205 ;
        RECT 92.190 695.720 96.410 698.205 ;
        RECT 97.250 695.720 101.930 698.205 ;
        RECT 102.770 695.720 106.990 698.205 ;
        RECT 107.830 695.720 112.510 698.205 ;
        RECT 113.350 695.720 117.570 698.205 ;
        RECT 118.410 695.720 123.090 698.205 ;
        RECT 123.930 695.720 128.150 698.205 ;
        RECT 128.990 695.720 133.670 698.205 ;
        RECT 134.510 695.720 138.730 698.205 ;
        RECT 139.570 695.720 143.790 698.205 ;
        RECT 144.630 695.720 149.310 698.205 ;
        RECT 150.150 695.720 154.370 698.205 ;
        RECT 155.210 695.720 159.890 698.205 ;
        RECT 160.730 695.720 164.950 698.205 ;
        RECT 165.790 695.720 170.470 698.205 ;
        RECT 171.310 695.720 175.530 698.205 ;
        RECT 176.370 695.720 181.050 698.205 ;
        RECT 181.890 695.720 186.110 698.205 ;
        RECT 186.950 695.720 191.170 698.205 ;
        RECT 192.010 695.720 196.690 698.205 ;
        RECT 197.530 695.720 201.750 698.205 ;
        RECT 202.590 695.720 207.270 698.205 ;
        RECT 208.110 695.720 212.330 698.205 ;
        RECT 213.170 695.720 217.850 698.205 ;
        RECT 218.690 695.720 222.910 698.205 ;
        RECT 223.750 695.720 228.430 698.205 ;
        RECT 229.270 695.720 233.490 698.205 ;
        RECT 234.330 695.720 238.550 698.205 ;
        RECT 239.390 695.720 244.070 698.205 ;
        RECT 244.910 695.720 249.130 698.205 ;
        RECT 249.970 695.720 254.650 698.205 ;
        RECT 255.490 695.720 259.710 698.205 ;
        RECT 260.550 695.720 265.230 698.205 ;
        RECT 266.070 695.720 270.290 698.205 ;
        RECT 271.130 695.720 275.810 698.205 ;
        RECT 276.650 695.720 280.870 698.205 ;
        RECT 281.710 695.720 285.930 698.205 ;
        RECT 286.770 695.720 291.450 698.205 ;
        RECT 292.290 695.720 296.510 698.205 ;
        RECT 297.350 695.720 302.030 698.205 ;
        RECT 302.870 695.720 307.090 698.205 ;
        RECT 307.930 695.720 312.610 698.205 ;
        RECT 313.450 695.720 317.670 698.205 ;
        RECT 318.510 695.720 323.190 698.205 ;
        RECT 324.030 695.720 328.250 698.205 ;
        RECT 329.090 695.720 333.310 698.205 ;
        RECT 334.150 695.720 338.830 698.205 ;
        RECT 339.670 695.720 343.890 698.205 ;
        RECT 344.730 695.720 349.410 698.205 ;
        RECT 350.250 695.720 354.470 698.205 ;
        RECT 355.310 695.720 359.990 698.205 ;
        RECT 360.830 695.720 365.050 698.205 ;
        RECT 365.890 695.720 370.570 698.205 ;
        RECT 371.410 695.720 375.630 698.205 ;
        RECT 376.470 695.720 380.690 698.205 ;
        RECT 381.530 695.720 386.210 698.205 ;
        RECT 387.050 695.720 391.270 698.205 ;
        RECT 392.110 695.720 396.790 698.205 ;
        RECT 397.630 695.720 401.850 698.205 ;
        RECT 402.690 695.720 407.370 698.205 ;
        RECT 408.210 695.720 412.430 698.205 ;
        RECT 413.270 695.720 417.950 698.205 ;
        RECT 418.790 695.720 423.010 698.205 ;
        RECT 423.850 695.720 428.070 698.205 ;
        RECT 428.910 695.720 433.590 698.205 ;
        RECT 434.430 695.720 438.650 698.205 ;
        RECT 439.490 695.720 444.170 698.205 ;
        RECT 445.010 695.720 449.230 698.205 ;
        RECT 450.070 695.720 454.750 698.205 ;
        RECT 455.590 695.720 459.810 698.205 ;
        RECT 460.650 695.720 465.330 698.205 ;
        RECT 466.170 695.720 470.390 698.205 ;
        RECT 471.230 695.720 475.450 698.205 ;
        RECT 476.290 695.720 480.970 698.205 ;
        RECT 481.810 695.720 486.030 698.205 ;
        RECT 486.870 695.720 491.550 698.205 ;
        RECT 492.390 695.720 496.610 698.205 ;
        RECT 497.450 695.720 502.130 698.205 ;
        RECT 502.970 695.720 507.190 698.205 ;
        RECT 508.030 695.720 512.710 698.205 ;
        RECT 513.550 695.720 517.770 698.205 ;
        RECT 518.610 695.720 522.830 698.205 ;
        RECT 523.670 695.720 528.350 698.205 ;
        RECT 529.190 695.720 533.410 698.205 ;
        RECT 534.250 695.720 538.930 698.205 ;
        RECT 539.770 695.720 543.990 698.205 ;
        RECT 544.830 695.720 549.510 698.205 ;
        RECT 550.350 695.720 554.570 698.205 ;
        RECT 555.410 695.720 560.090 698.205 ;
        RECT 560.930 695.720 565.150 698.205 ;
        RECT 565.990 695.720 570.210 698.205 ;
        RECT 571.050 695.720 575.730 698.205 ;
        RECT 576.570 695.720 580.790 698.205 ;
        RECT 581.630 695.720 586.310 698.205 ;
        RECT 587.150 695.720 591.370 698.205 ;
        RECT 592.210 695.720 596.890 698.205 ;
        RECT 597.730 695.720 601.950 698.205 ;
        RECT 602.790 695.720 607.470 698.205 ;
        RECT 608.310 695.720 612.530 698.205 ;
        RECT 613.370 695.720 617.590 698.205 ;
        RECT 618.430 695.720 623.110 698.205 ;
        RECT 623.950 695.720 628.170 698.205 ;
        RECT 629.010 695.720 633.690 698.205 ;
        RECT 634.530 695.720 638.750 698.205 ;
        RECT 639.590 695.720 644.270 698.205 ;
        RECT 645.110 695.720 649.330 698.205 ;
        RECT 650.170 695.720 654.850 698.205 ;
        RECT 655.690 695.720 659.910 698.205 ;
        RECT 660.750 695.720 664.970 698.205 ;
        RECT 665.810 695.720 670.490 698.205 ;
        RECT 671.330 695.720 675.550 698.205 ;
        RECT 676.390 695.720 681.070 698.205 ;
        RECT 681.910 695.720 686.130 698.205 ;
        RECT 686.970 695.720 691.650 698.205 ;
        RECT 692.490 695.720 696.710 698.205 ;
        RECT 2.400 4.280 697.260 695.720 ;
        RECT 2.400 1.515 3.030 4.280 ;
        RECT 3.870 1.515 9.470 4.280 ;
        RECT 10.310 1.515 15.910 4.280 ;
        RECT 16.750 1.515 22.810 4.280 ;
        RECT 23.650 1.515 29.250 4.280 ;
        RECT 30.090 1.515 35.690 4.280 ;
        RECT 36.530 1.515 42.590 4.280 ;
        RECT 43.430 1.515 49.030 4.280 ;
        RECT 49.870 1.515 55.470 4.280 ;
        RECT 56.310 1.515 62.370 4.280 ;
        RECT 63.210 1.515 68.810 4.280 ;
        RECT 69.650 1.515 75.250 4.280 ;
        RECT 76.090 1.515 82.150 4.280 ;
        RECT 82.990 1.515 88.590 4.280 ;
        RECT 89.430 1.515 95.490 4.280 ;
        RECT 96.330 1.515 101.930 4.280 ;
        RECT 102.770 1.515 108.370 4.280 ;
        RECT 109.210 1.515 115.270 4.280 ;
        RECT 116.110 1.515 121.710 4.280 ;
        RECT 122.550 1.515 128.150 4.280 ;
        RECT 128.990 1.515 135.050 4.280 ;
        RECT 135.890 1.515 141.490 4.280 ;
        RECT 142.330 1.515 147.930 4.280 ;
        RECT 148.770 1.515 154.830 4.280 ;
        RECT 155.670 1.515 161.270 4.280 ;
        RECT 162.110 1.515 167.710 4.280 ;
        RECT 168.550 1.515 174.610 4.280 ;
        RECT 175.450 1.515 181.050 4.280 ;
        RECT 181.890 1.515 187.950 4.280 ;
        RECT 188.790 1.515 194.390 4.280 ;
        RECT 195.230 1.515 200.830 4.280 ;
        RECT 201.670 1.515 207.730 4.280 ;
        RECT 208.570 1.515 214.170 4.280 ;
        RECT 215.010 1.515 220.610 4.280 ;
        RECT 221.450 1.515 227.510 4.280 ;
        RECT 228.350 1.515 233.950 4.280 ;
        RECT 234.790 1.515 240.390 4.280 ;
        RECT 241.230 1.515 247.290 4.280 ;
        RECT 248.130 1.515 253.730 4.280 ;
        RECT 254.570 1.515 260.170 4.280 ;
        RECT 261.010 1.515 267.070 4.280 ;
        RECT 267.910 1.515 273.510 4.280 ;
        RECT 274.350 1.515 280.410 4.280 ;
        RECT 281.250 1.515 286.850 4.280 ;
        RECT 287.690 1.515 293.290 4.280 ;
        RECT 294.130 1.515 300.190 4.280 ;
        RECT 301.030 1.515 306.630 4.280 ;
        RECT 307.470 1.515 313.070 4.280 ;
        RECT 313.910 1.515 319.970 4.280 ;
        RECT 320.810 1.515 326.410 4.280 ;
        RECT 327.250 1.515 332.850 4.280 ;
        RECT 333.690 1.515 339.750 4.280 ;
        RECT 340.590 1.515 346.190 4.280 ;
        RECT 347.030 1.515 353.090 4.280 ;
        RECT 353.930 1.515 359.530 4.280 ;
        RECT 360.370 1.515 365.970 4.280 ;
        RECT 366.810 1.515 372.870 4.280 ;
        RECT 373.710 1.515 379.310 4.280 ;
        RECT 380.150 1.515 385.750 4.280 ;
        RECT 386.590 1.515 392.650 4.280 ;
        RECT 393.490 1.515 399.090 4.280 ;
        RECT 399.930 1.515 405.530 4.280 ;
        RECT 406.370 1.515 412.430 4.280 ;
        RECT 413.270 1.515 418.870 4.280 ;
        RECT 419.710 1.515 425.310 4.280 ;
        RECT 426.150 1.515 432.210 4.280 ;
        RECT 433.050 1.515 438.650 4.280 ;
        RECT 439.490 1.515 445.550 4.280 ;
        RECT 446.390 1.515 451.990 4.280 ;
        RECT 452.830 1.515 458.430 4.280 ;
        RECT 459.270 1.515 465.330 4.280 ;
        RECT 466.170 1.515 471.770 4.280 ;
        RECT 472.610 1.515 478.210 4.280 ;
        RECT 479.050 1.515 485.110 4.280 ;
        RECT 485.950 1.515 491.550 4.280 ;
        RECT 492.390 1.515 497.990 4.280 ;
        RECT 498.830 1.515 504.890 4.280 ;
        RECT 505.730 1.515 511.330 4.280 ;
        RECT 512.170 1.515 517.770 4.280 ;
        RECT 518.610 1.515 524.670 4.280 ;
        RECT 525.510 1.515 531.110 4.280 ;
        RECT 531.950 1.515 538.010 4.280 ;
        RECT 538.850 1.515 544.450 4.280 ;
        RECT 545.290 1.515 550.890 4.280 ;
        RECT 551.730 1.515 557.790 4.280 ;
        RECT 558.630 1.515 564.230 4.280 ;
        RECT 565.070 1.515 570.670 4.280 ;
        RECT 571.510 1.515 577.570 4.280 ;
        RECT 578.410 1.515 584.010 4.280 ;
        RECT 584.850 1.515 590.450 4.280 ;
        RECT 591.290 1.515 597.350 4.280 ;
        RECT 598.190 1.515 603.790 4.280 ;
        RECT 604.630 1.515 610.230 4.280 ;
        RECT 611.070 1.515 617.130 4.280 ;
        RECT 617.970 1.515 623.570 4.280 ;
        RECT 624.410 1.515 630.470 4.280 ;
        RECT 631.310 1.515 636.910 4.280 ;
        RECT 637.750 1.515 643.350 4.280 ;
        RECT 644.190 1.515 650.250 4.280 ;
        RECT 651.090 1.515 656.690 4.280 ;
        RECT 657.530 1.515 663.130 4.280 ;
        RECT 663.970 1.515 670.030 4.280 ;
        RECT 670.870 1.515 676.470 4.280 ;
        RECT 677.310 1.515 682.910 4.280 ;
        RECT 683.750 1.515 689.810 4.280 ;
        RECT 690.650 1.515 696.250 4.280 ;
        RECT 697.090 1.515 697.260 4.280 ;
      LAYER met3 ;
        RECT 4.400 697.320 696.000 698.185 ;
        RECT 4.000 695.320 696.000 697.320 ;
        RECT 4.400 693.920 696.000 695.320 ;
        RECT 4.000 691.920 696.000 693.920 ;
        RECT 4.400 690.520 696.000 691.920 ;
        RECT 4.000 689.200 696.000 690.520 ;
        RECT 4.400 688.520 696.000 689.200 ;
        RECT 4.400 687.800 695.600 688.520 ;
        RECT 4.000 687.120 695.600 687.800 ;
        RECT 4.000 685.800 696.000 687.120 ;
        RECT 4.400 684.400 696.000 685.800 ;
        RECT 4.000 682.400 696.000 684.400 ;
        RECT 4.400 681.000 696.000 682.400 ;
        RECT 4.000 679.000 696.000 681.000 ;
        RECT 4.400 677.600 696.000 679.000 ;
        RECT 4.000 676.280 696.000 677.600 ;
        RECT 4.400 674.880 696.000 676.280 ;
        RECT 4.000 672.880 696.000 674.880 ;
        RECT 4.400 671.480 696.000 672.880 ;
        RECT 4.000 669.480 696.000 671.480 ;
        RECT 4.400 668.080 696.000 669.480 ;
        RECT 4.000 666.760 696.000 668.080 ;
        RECT 4.400 665.400 696.000 666.760 ;
        RECT 4.400 665.360 695.600 665.400 ;
        RECT 4.000 664.000 695.600 665.360 ;
        RECT 4.000 663.360 696.000 664.000 ;
        RECT 4.400 661.960 696.000 663.360 ;
        RECT 4.000 659.960 696.000 661.960 ;
        RECT 4.400 658.560 696.000 659.960 ;
        RECT 4.000 656.560 696.000 658.560 ;
        RECT 4.400 655.160 696.000 656.560 ;
        RECT 4.000 653.840 696.000 655.160 ;
        RECT 4.400 652.440 696.000 653.840 ;
        RECT 4.000 650.440 696.000 652.440 ;
        RECT 4.400 649.040 696.000 650.440 ;
        RECT 4.000 647.040 696.000 649.040 ;
        RECT 4.400 645.640 696.000 647.040 ;
        RECT 4.000 644.320 696.000 645.640 ;
        RECT 4.400 642.920 696.000 644.320 ;
        RECT 4.000 642.280 696.000 642.920 ;
        RECT 4.000 640.920 695.600 642.280 ;
        RECT 4.400 640.880 695.600 640.920 ;
        RECT 4.400 639.520 696.000 640.880 ;
        RECT 4.000 637.520 696.000 639.520 ;
        RECT 4.400 636.120 696.000 637.520 ;
        RECT 4.000 634.120 696.000 636.120 ;
        RECT 4.400 632.720 696.000 634.120 ;
        RECT 4.000 631.400 696.000 632.720 ;
        RECT 4.400 630.000 696.000 631.400 ;
        RECT 4.000 628.000 696.000 630.000 ;
        RECT 4.400 626.600 696.000 628.000 ;
        RECT 4.000 624.600 696.000 626.600 ;
        RECT 4.400 623.200 696.000 624.600 ;
        RECT 4.000 621.200 696.000 623.200 ;
        RECT 4.400 619.800 696.000 621.200 ;
        RECT 4.000 618.480 696.000 619.800 ;
        RECT 4.400 617.080 695.600 618.480 ;
        RECT 4.000 615.080 696.000 617.080 ;
        RECT 4.400 613.680 696.000 615.080 ;
        RECT 4.000 611.680 696.000 613.680 ;
        RECT 4.400 610.280 696.000 611.680 ;
        RECT 4.000 608.960 696.000 610.280 ;
        RECT 4.400 607.560 696.000 608.960 ;
        RECT 4.000 605.560 696.000 607.560 ;
        RECT 4.400 604.160 696.000 605.560 ;
        RECT 4.000 602.160 696.000 604.160 ;
        RECT 4.400 600.760 696.000 602.160 ;
        RECT 4.000 598.760 696.000 600.760 ;
        RECT 4.400 597.360 696.000 598.760 ;
        RECT 4.000 596.040 696.000 597.360 ;
        RECT 4.400 595.360 696.000 596.040 ;
        RECT 4.400 594.640 695.600 595.360 ;
        RECT 4.000 593.960 695.600 594.640 ;
        RECT 4.000 592.640 696.000 593.960 ;
        RECT 4.400 591.240 696.000 592.640 ;
        RECT 4.000 589.240 696.000 591.240 ;
        RECT 4.400 587.840 696.000 589.240 ;
        RECT 4.000 586.520 696.000 587.840 ;
        RECT 4.400 585.120 696.000 586.520 ;
        RECT 4.000 583.120 696.000 585.120 ;
        RECT 4.400 581.720 696.000 583.120 ;
        RECT 4.000 579.720 696.000 581.720 ;
        RECT 4.400 578.320 696.000 579.720 ;
        RECT 4.000 576.320 696.000 578.320 ;
        RECT 4.400 574.920 696.000 576.320 ;
        RECT 4.000 573.600 696.000 574.920 ;
        RECT 4.400 572.240 696.000 573.600 ;
        RECT 4.400 572.200 695.600 572.240 ;
        RECT 4.000 570.840 695.600 572.200 ;
        RECT 4.000 570.200 696.000 570.840 ;
        RECT 4.400 568.800 696.000 570.200 ;
        RECT 4.000 566.800 696.000 568.800 ;
        RECT 4.400 565.400 696.000 566.800 ;
        RECT 4.000 564.080 696.000 565.400 ;
        RECT 4.400 562.680 696.000 564.080 ;
        RECT 4.000 560.680 696.000 562.680 ;
        RECT 4.400 559.280 696.000 560.680 ;
        RECT 4.000 557.280 696.000 559.280 ;
        RECT 4.400 555.880 696.000 557.280 ;
        RECT 4.000 553.880 696.000 555.880 ;
        RECT 4.400 552.480 696.000 553.880 ;
        RECT 4.000 551.160 696.000 552.480 ;
        RECT 4.400 549.760 696.000 551.160 ;
        RECT 4.000 548.440 696.000 549.760 ;
        RECT 4.000 547.760 695.600 548.440 ;
        RECT 4.400 547.040 695.600 547.760 ;
        RECT 4.400 546.360 696.000 547.040 ;
        RECT 4.000 544.360 696.000 546.360 ;
        RECT 4.400 542.960 696.000 544.360 ;
        RECT 4.000 540.960 696.000 542.960 ;
        RECT 4.400 539.560 696.000 540.960 ;
        RECT 4.000 538.240 696.000 539.560 ;
        RECT 4.400 536.840 696.000 538.240 ;
        RECT 4.000 534.840 696.000 536.840 ;
        RECT 4.400 533.440 696.000 534.840 ;
        RECT 4.000 531.440 696.000 533.440 ;
        RECT 4.400 530.040 696.000 531.440 ;
        RECT 4.000 528.720 696.000 530.040 ;
        RECT 4.400 527.320 696.000 528.720 ;
        RECT 4.000 525.320 696.000 527.320 ;
        RECT 4.400 523.920 695.600 525.320 ;
        RECT 4.000 521.920 696.000 523.920 ;
        RECT 4.400 520.520 696.000 521.920 ;
        RECT 4.000 518.520 696.000 520.520 ;
        RECT 4.400 517.120 696.000 518.520 ;
        RECT 4.000 515.800 696.000 517.120 ;
        RECT 4.400 514.400 696.000 515.800 ;
        RECT 4.000 512.400 696.000 514.400 ;
        RECT 4.400 511.000 696.000 512.400 ;
        RECT 4.000 509.000 696.000 511.000 ;
        RECT 4.400 507.600 696.000 509.000 ;
        RECT 4.000 506.280 696.000 507.600 ;
        RECT 4.400 504.880 696.000 506.280 ;
        RECT 4.000 502.880 696.000 504.880 ;
        RECT 4.400 502.200 696.000 502.880 ;
        RECT 4.400 501.480 695.600 502.200 ;
        RECT 4.000 500.800 695.600 501.480 ;
        RECT 4.000 499.480 696.000 500.800 ;
        RECT 4.400 498.080 696.000 499.480 ;
        RECT 4.000 496.080 696.000 498.080 ;
        RECT 4.400 494.680 696.000 496.080 ;
        RECT 4.000 493.360 696.000 494.680 ;
        RECT 4.400 491.960 696.000 493.360 ;
        RECT 4.000 489.960 696.000 491.960 ;
        RECT 4.400 488.560 696.000 489.960 ;
        RECT 4.000 486.560 696.000 488.560 ;
        RECT 4.400 485.160 696.000 486.560 ;
        RECT 4.000 483.840 696.000 485.160 ;
        RECT 4.400 482.440 696.000 483.840 ;
        RECT 4.000 480.440 696.000 482.440 ;
        RECT 4.400 479.080 696.000 480.440 ;
        RECT 4.400 479.040 695.600 479.080 ;
        RECT 4.000 477.680 695.600 479.040 ;
        RECT 4.000 477.040 696.000 477.680 ;
        RECT 4.400 475.640 696.000 477.040 ;
        RECT 4.000 473.640 696.000 475.640 ;
        RECT 4.400 472.240 696.000 473.640 ;
        RECT 4.000 470.920 696.000 472.240 ;
        RECT 4.400 469.520 696.000 470.920 ;
        RECT 4.000 467.520 696.000 469.520 ;
        RECT 4.400 466.120 696.000 467.520 ;
        RECT 4.000 464.120 696.000 466.120 ;
        RECT 4.400 462.720 696.000 464.120 ;
        RECT 4.000 460.720 696.000 462.720 ;
        RECT 4.400 459.320 696.000 460.720 ;
        RECT 4.000 458.000 696.000 459.320 ;
        RECT 4.400 456.600 696.000 458.000 ;
        RECT 4.000 455.280 696.000 456.600 ;
        RECT 4.000 454.600 695.600 455.280 ;
        RECT 4.400 453.880 695.600 454.600 ;
        RECT 4.400 453.200 696.000 453.880 ;
        RECT 4.000 451.200 696.000 453.200 ;
        RECT 4.400 449.800 696.000 451.200 ;
        RECT 4.000 448.480 696.000 449.800 ;
        RECT 4.400 447.080 696.000 448.480 ;
        RECT 4.000 445.080 696.000 447.080 ;
        RECT 4.400 443.680 696.000 445.080 ;
        RECT 4.000 441.680 696.000 443.680 ;
        RECT 4.400 440.280 696.000 441.680 ;
        RECT 4.000 438.280 696.000 440.280 ;
        RECT 4.400 436.880 696.000 438.280 ;
        RECT 4.000 435.560 696.000 436.880 ;
        RECT 4.400 434.160 696.000 435.560 ;
        RECT 4.000 432.160 696.000 434.160 ;
        RECT 4.400 430.760 695.600 432.160 ;
        RECT 4.000 428.760 696.000 430.760 ;
        RECT 4.400 427.360 696.000 428.760 ;
        RECT 4.000 426.040 696.000 427.360 ;
        RECT 4.400 424.640 696.000 426.040 ;
        RECT 4.000 422.640 696.000 424.640 ;
        RECT 4.400 421.240 696.000 422.640 ;
        RECT 4.000 419.240 696.000 421.240 ;
        RECT 4.400 417.840 696.000 419.240 ;
        RECT 4.000 415.840 696.000 417.840 ;
        RECT 4.400 414.440 696.000 415.840 ;
        RECT 4.000 413.120 696.000 414.440 ;
        RECT 4.400 411.720 696.000 413.120 ;
        RECT 4.000 409.720 696.000 411.720 ;
        RECT 4.400 409.040 696.000 409.720 ;
        RECT 4.400 408.320 695.600 409.040 ;
        RECT 4.000 407.640 695.600 408.320 ;
        RECT 4.000 406.320 696.000 407.640 ;
        RECT 4.400 404.920 696.000 406.320 ;
        RECT 4.000 403.600 696.000 404.920 ;
        RECT 4.400 402.200 696.000 403.600 ;
        RECT 4.000 400.200 696.000 402.200 ;
        RECT 4.400 398.800 696.000 400.200 ;
        RECT 4.000 396.800 696.000 398.800 ;
        RECT 4.400 395.400 696.000 396.800 ;
        RECT 4.000 393.400 696.000 395.400 ;
        RECT 4.400 392.000 696.000 393.400 ;
        RECT 4.000 390.680 696.000 392.000 ;
        RECT 4.400 389.280 696.000 390.680 ;
        RECT 4.000 387.280 696.000 389.280 ;
        RECT 4.400 385.880 696.000 387.280 ;
        RECT 4.000 385.240 696.000 385.880 ;
        RECT 4.000 383.880 695.600 385.240 ;
        RECT 4.400 383.840 695.600 383.880 ;
        RECT 4.400 382.480 696.000 383.840 ;
        RECT 4.000 380.480 696.000 382.480 ;
        RECT 4.400 379.080 696.000 380.480 ;
        RECT 4.000 377.760 696.000 379.080 ;
        RECT 4.400 376.360 696.000 377.760 ;
        RECT 4.000 374.360 696.000 376.360 ;
        RECT 4.400 372.960 696.000 374.360 ;
        RECT 4.000 370.960 696.000 372.960 ;
        RECT 4.400 369.560 696.000 370.960 ;
        RECT 4.000 368.240 696.000 369.560 ;
        RECT 4.400 366.840 696.000 368.240 ;
        RECT 4.000 364.840 696.000 366.840 ;
        RECT 4.400 363.440 696.000 364.840 ;
        RECT 4.000 362.120 696.000 363.440 ;
        RECT 4.000 361.440 695.600 362.120 ;
        RECT 4.400 360.720 695.600 361.440 ;
        RECT 4.400 360.040 696.000 360.720 ;
        RECT 4.000 358.040 696.000 360.040 ;
        RECT 4.400 356.640 696.000 358.040 ;
        RECT 4.000 355.320 696.000 356.640 ;
        RECT 4.400 353.920 696.000 355.320 ;
        RECT 4.000 351.920 696.000 353.920 ;
        RECT 4.400 350.520 696.000 351.920 ;
        RECT 4.000 348.520 696.000 350.520 ;
        RECT 4.400 347.120 696.000 348.520 ;
        RECT 4.000 345.800 696.000 347.120 ;
        RECT 4.400 344.400 696.000 345.800 ;
        RECT 4.000 342.400 696.000 344.400 ;
        RECT 4.400 341.000 696.000 342.400 ;
        RECT 4.000 339.000 696.000 341.000 ;
        RECT 4.400 337.600 695.600 339.000 ;
        RECT 4.000 335.600 696.000 337.600 ;
        RECT 4.400 334.200 696.000 335.600 ;
        RECT 4.000 332.880 696.000 334.200 ;
        RECT 4.400 331.480 696.000 332.880 ;
        RECT 4.000 329.480 696.000 331.480 ;
        RECT 4.400 328.080 696.000 329.480 ;
        RECT 4.000 326.080 696.000 328.080 ;
        RECT 4.400 324.680 696.000 326.080 ;
        RECT 4.000 323.360 696.000 324.680 ;
        RECT 4.400 321.960 696.000 323.360 ;
        RECT 4.000 319.960 696.000 321.960 ;
        RECT 4.400 318.560 696.000 319.960 ;
        RECT 4.000 316.560 696.000 318.560 ;
        RECT 4.400 315.200 696.000 316.560 ;
        RECT 4.400 315.160 695.600 315.200 ;
        RECT 4.000 313.800 695.600 315.160 ;
        RECT 4.000 313.160 696.000 313.800 ;
        RECT 4.400 311.760 696.000 313.160 ;
        RECT 4.000 310.440 696.000 311.760 ;
        RECT 4.400 309.040 696.000 310.440 ;
        RECT 4.000 307.040 696.000 309.040 ;
        RECT 4.400 305.640 696.000 307.040 ;
        RECT 4.000 303.640 696.000 305.640 ;
        RECT 4.400 302.240 696.000 303.640 ;
        RECT 4.000 300.240 696.000 302.240 ;
        RECT 4.400 298.840 696.000 300.240 ;
        RECT 4.000 297.520 696.000 298.840 ;
        RECT 4.400 296.120 696.000 297.520 ;
        RECT 4.000 294.120 696.000 296.120 ;
        RECT 4.400 292.720 696.000 294.120 ;
        RECT 4.000 292.080 696.000 292.720 ;
        RECT 4.000 290.720 695.600 292.080 ;
        RECT 4.400 290.680 695.600 290.720 ;
        RECT 4.400 289.320 696.000 290.680 ;
        RECT 4.000 288.000 696.000 289.320 ;
        RECT 4.400 286.600 696.000 288.000 ;
        RECT 4.000 284.600 696.000 286.600 ;
        RECT 4.400 283.200 696.000 284.600 ;
        RECT 4.000 281.200 696.000 283.200 ;
        RECT 4.400 279.800 696.000 281.200 ;
        RECT 4.000 277.800 696.000 279.800 ;
        RECT 4.400 276.400 696.000 277.800 ;
        RECT 4.000 275.080 696.000 276.400 ;
        RECT 4.400 273.680 696.000 275.080 ;
        RECT 4.000 271.680 696.000 273.680 ;
        RECT 4.400 270.280 696.000 271.680 ;
        RECT 4.000 268.960 696.000 270.280 ;
        RECT 4.000 268.280 695.600 268.960 ;
        RECT 4.400 267.560 695.600 268.280 ;
        RECT 4.400 266.880 696.000 267.560 ;
        RECT 4.000 265.560 696.000 266.880 ;
        RECT 4.400 264.160 696.000 265.560 ;
        RECT 4.000 262.160 696.000 264.160 ;
        RECT 4.400 260.760 696.000 262.160 ;
        RECT 4.000 258.760 696.000 260.760 ;
        RECT 4.400 257.360 696.000 258.760 ;
        RECT 4.000 255.360 696.000 257.360 ;
        RECT 4.400 253.960 696.000 255.360 ;
        RECT 4.000 252.640 696.000 253.960 ;
        RECT 4.400 251.240 696.000 252.640 ;
        RECT 4.000 249.240 696.000 251.240 ;
        RECT 4.400 247.840 696.000 249.240 ;
        RECT 4.000 245.840 696.000 247.840 ;
        RECT 4.400 244.440 695.600 245.840 ;
        RECT 4.000 243.120 696.000 244.440 ;
        RECT 4.400 241.720 696.000 243.120 ;
        RECT 4.000 239.720 696.000 241.720 ;
        RECT 4.400 238.320 696.000 239.720 ;
        RECT 4.000 236.320 696.000 238.320 ;
        RECT 4.400 234.920 696.000 236.320 ;
        RECT 4.000 232.920 696.000 234.920 ;
        RECT 4.400 231.520 696.000 232.920 ;
        RECT 4.000 230.200 696.000 231.520 ;
        RECT 4.400 228.800 696.000 230.200 ;
        RECT 4.000 226.800 696.000 228.800 ;
        RECT 4.400 225.400 696.000 226.800 ;
        RECT 4.000 223.400 696.000 225.400 ;
        RECT 4.400 222.040 696.000 223.400 ;
        RECT 4.400 222.000 695.600 222.040 ;
        RECT 4.000 220.640 695.600 222.000 ;
        RECT 4.000 220.000 696.000 220.640 ;
        RECT 4.400 218.600 696.000 220.000 ;
        RECT 4.000 217.280 696.000 218.600 ;
        RECT 4.400 215.880 696.000 217.280 ;
        RECT 4.000 213.880 696.000 215.880 ;
        RECT 4.400 212.480 696.000 213.880 ;
        RECT 4.000 210.480 696.000 212.480 ;
        RECT 4.400 209.080 696.000 210.480 ;
        RECT 4.000 207.760 696.000 209.080 ;
        RECT 4.400 206.360 696.000 207.760 ;
        RECT 4.000 204.360 696.000 206.360 ;
        RECT 4.400 202.960 696.000 204.360 ;
        RECT 4.000 200.960 696.000 202.960 ;
        RECT 4.400 199.560 696.000 200.960 ;
        RECT 4.000 198.920 696.000 199.560 ;
        RECT 4.000 197.560 695.600 198.920 ;
        RECT 4.400 197.520 695.600 197.560 ;
        RECT 4.400 196.160 696.000 197.520 ;
        RECT 4.000 194.840 696.000 196.160 ;
        RECT 4.400 193.440 696.000 194.840 ;
        RECT 4.000 191.440 696.000 193.440 ;
        RECT 4.400 190.040 696.000 191.440 ;
        RECT 4.000 188.040 696.000 190.040 ;
        RECT 4.400 186.640 696.000 188.040 ;
        RECT 4.000 185.320 696.000 186.640 ;
        RECT 4.400 183.920 696.000 185.320 ;
        RECT 4.000 181.920 696.000 183.920 ;
        RECT 4.400 180.520 696.000 181.920 ;
        RECT 4.000 178.520 696.000 180.520 ;
        RECT 4.400 177.120 696.000 178.520 ;
        RECT 4.000 175.800 696.000 177.120 ;
        RECT 4.000 175.120 695.600 175.800 ;
        RECT 4.400 174.400 695.600 175.120 ;
        RECT 4.400 173.720 696.000 174.400 ;
        RECT 4.000 172.400 696.000 173.720 ;
        RECT 4.400 171.000 696.000 172.400 ;
        RECT 4.000 169.000 696.000 171.000 ;
        RECT 4.400 167.600 696.000 169.000 ;
        RECT 4.000 165.600 696.000 167.600 ;
        RECT 4.400 164.200 696.000 165.600 ;
        RECT 4.000 162.880 696.000 164.200 ;
        RECT 4.400 161.480 696.000 162.880 ;
        RECT 4.000 159.480 696.000 161.480 ;
        RECT 4.400 158.080 696.000 159.480 ;
        RECT 4.000 156.080 696.000 158.080 ;
        RECT 4.400 154.680 696.000 156.080 ;
        RECT 4.000 152.680 696.000 154.680 ;
        RECT 4.400 152.000 696.000 152.680 ;
        RECT 4.400 151.280 695.600 152.000 ;
        RECT 4.000 150.600 695.600 151.280 ;
        RECT 4.000 149.960 696.000 150.600 ;
        RECT 4.400 148.560 696.000 149.960 ;
        RECT 4.000 146.560 696.000 148.560 ;
        RECT 4.400 145.160 696.000 146.560 ;
        RECT 4.000 143.160 696.000 145.160 ;
        RECT 4.400 141.760 696.000 143.160 ;
        RECT 4.000 139.760 696.000 141.760 ;
        RECT 4.400 138.360 696.000 139.760 ;
        RECT 4.000 137.040 696.000 138.360 ;
        RECT 4.400 135.640 696.000 137.040 ;
        RECT 4.000 133.640 696.000 135.640 ;
        RECT 4.400 132.240 696.000 133.640 ;
        RECT 4.000 130.240 696.000 132.240 ;
        RECT 4.400 128.880 696.000 130.240 ;
        RECT 4.400 128.840 695.600 128.880 ;
        RECT 4.000 127.520 695.600 128.840 ;
        RECT 4.400 127.480 695.600 127.520 ;
        RECT 4.400 126.120 696.000 127.480 ;
        RECT 4.000 124.120 696.000 126.120 ;
        RECT 4.400 122.720 696.000 124.120 ;
        RECT 4.000 120.720 696.000 122.720 ;
        RECT 4.400 119.320 696.000 120.720 ;
        RECT 4.000 117.320 696.000 119.320 ;
        RECT 4.400 115.920 696.000 117.320 ;
        RECT 4.000 114.600 696.000 115.920 ;
        RECT 4.400 113.200 696.000 114.600 ;
        RECT 4.000 111.200 696.000 113.200 ;
        RECT 4.400 109.800 696.000 111.200 ;
        RECT 4.000 107.800 696.000 109.800 ;
        RECT 4.400 106.400 696.000 107.800 ;
        RECT 4.000 105.760 696.000 106.400 ;
        RECT 4.000 105.080 695.600 105.760 ;
        RECT 4.400 104.360 695.600 105.080 ;
        RECT 4.400 103.680 696.000 104.360 ;
        RECT 4.000 101.680 696.000 103.680 ;
        RECT 4.400 100.280 696.000 101.680 ;
        RECT 4.000 98.280 696.000 100.280 ;
        RECT 4.400 96.880 696.000 98.280 ;
        RECT 4.000 94.880 696.000 96.880 ;
        RECT 4.400 93.480 696.000 94.880 ;
        RECT 4.000 92.160 696.000 93.480 ;
        RECT 4.400 90.760 696.000 92.160 ;
        RECT 4.000 88.760 696.000 90.760 ;
        RECT 4.400 87.360 696.000 88.760 ;
        RECT 4.000 85.360 696.000 87.360 ;
        RECT 4.400 83.960 696.000 85.360 ;
        RECT 4.000 82.640 696.000 83.960 ;
        RECT 4.400 81.960 696.000 82.640 ;
        RECT 4.400 81.240 695.600 81.960 ;
        RECT 4.000 80.560 695.600 81.240 ;
        RECT 4.000 79.240 696.000 80.560 ;
        RECT 4.400 77.840 696.000 79.240 ;
        RECT 4.000 75.840 696.000 77.840 ;
        RECT 4.400 74.440 696.000 75.840 ;
        RECT 4.000 72.440 696.000 74.440 ;
        RECT 4.400 71.040 696.000 72.440 ;
        RECT 4.000 69.720 696.000 71.040 ;
        RECT 4.400 68.320 696.000 69.720 ;
        RECT 4.000 66.320 696.000 68.320 ;
        RECT 4.400 64.920 696.000 66.320 ;
        RECT 4.000 62.920 696.000 64.920 ;
        RECT 4.400 61.520 696.000 62.920 ;
        RECT 4.000 59.520 696.000 61.520 ;
        RECT 4.400 58.840 696.000 59.520 ;
        RECT 4.400 58.120 695.600 58.840 ;
        RECT 4.000 57.440 695.600 58.120 ;
        RECT 4.000 56.800 696.000 57.440 ;
        RECT 4.400 55.400 696.000 56.800 ;
        RECT 4.000 53.400 696.000 55.400 ;
        RECT 4.400 52.000 696.000 53.400 ;
        RECT 4.000 50.000 696.000 52.000 ;
        RECT 4.400 48.600 696.000 50.000 ;
        RECT 4.000 47.280 696.000 48.600 ;
        RECT 4.400 45.880 696.000 47.280 ;
        RECT 4.000 43.880 696.000 45.880 ;
        RECT 4.400 42.480 696.000 43.880 ;
        RECT 4.000 40.480 696.000 42.480 ;
        RECT 4.400 39.080 696.000 40.480 ;
        RECT 4.000 37.080 696.000 39.080 ;
        RECT 4.400 35.720 696.000 37.080 ;
        RECT 4.400 35.680 695.600 35.720 ;
        RECT 4.000 34.360 695.600 35.680 ;
        RECT 4.400 34.320 695.600 34.360 ;
        RECT 4.400 32.960 696.000 34.320 ;
        RECT 4.000 30.960 696.000 32.960 ;
        RECT 4.400 29.560 696.000 30.960 ;
        RECT 4.000 27.560 696.000 29.560 ;
        RECT 4.400 26.160 696.000 27.560 ;
        RECT 4.000 24.840 696.000 26.160 ;
        RECT 4.400 23.440 696.000 24.840 ;
        RECT 4.000 21.440 696.000 23.440 ;
        RECT 4.400 20.040 696.000 21.440 ;
        RECT 4.000 18.040 696.000 20.040 ;
        RECT 4.400 16.640 696.000 18.040 ;
        RECT 4.000 14.640 696.000 16.640 ;
        RECT 4.400 13.240 696.000 14.640 ;
        RECT 4.000 12.600 696.000 13.240 ;
        RECT 4.000 11.920 695.600 12.600 ;
        RECT 4.400 11.200 695.600 11.920 ;
        RECT 4.400 10.520 696.000 11.200 ;
        RECT 4.000 8.520 696.000 10.520 ;
        RECT 4.400 7.120 696.000 8.520 ;
        RECT 4.000 5.120 696.000 7.120 ;
        RECT 4.400 3.720 696.000 5.120 ;
        RECT 4.000 2.400 696.000 3.720 ;
        RECT 4.400 1.535 696.000 2.400 ;
  END
END vco_adc_wrapper
END LIBRARY

