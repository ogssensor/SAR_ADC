magic
tech sky130A
magscale 1 2
timestamp 1624100228
<< obsli1 >>
rect 1104 1445 178848 117521
<< obsm1 >>
rect 750 212 179294 117552
<< metal2 >>
rect 754 119200 810 120000
rect 2226 119200 2282 120000
rect 3698 119200 3754 120000
rect 5170 119200 5226 120000
rect 6642 119200 6698 120000
rect 8114 119200 8170 120000
rect 9586 119200 9642 120000
rect 11058 119200 11114 120000
rect 12530 119200 12586 120000
rect 14002 119200 14058 120000
rect 15474 119200 15530 120000
rect 16946 119200 17002 120000
rect 18418 119200 18474 120000
rect 19890 119200 19946 120000
rect 21362 119200 21418 120000
rect 22834 119200 22890 120000
rect 24306 119200 24362 120000
rect 25778 119200 25834 120000
rect 27250 119200 27306 120000
rect 28722 119200 28778 120000
rect 30194 119200 30250 120000
rect 31666 119200 31722 120000
rect 33138 119200 33194 120000
rect 34610 119200 34666 120000
rect 36082 119200 36138 120000
rect 37646 119200 37702 120000
rect 39118 119200 39174 120000
rect 40590 119200 40646 120000
rect 42062 119200 42118 120000
rect 43534 119200 43590 120000
rect 45006 119200 45062 120000
rect 46478 119200 46534 120000
rect 47950 119200 48006 120000
rect 49422 119200 49478 120000
rect 50894 119200 50950 120000
rect 52366 119200 52422 120000
rect 53838 119200 53894 120000
rect 55310 119200 55366 120000
rect 56782 119200 56838 120000
rect 58254 119200 58310 120000
rect 59726 119200 59782 120000
rect 61198 119200 61254 120000
rect 62670 119200 62726 120000
rect 64142 119200 64198 120000
rect 65614 119200 65670 120000
rect 67086 119200 67142 120000
rect 68558 119200 68614 120000
rect 70030 119200 70086 120000
rect 71502 119200 71558 120000
rect 73066 119200 73122 120000
rect 74538 119200 74594 120000
rect 76010 119200 76066 120000
rect 77482 119200 77538 120000
rect 78954 119200 79010 120000
rect 80426 119200 80482 120000
rect 81898 119200 81954 120000
rect 83370 119200 83426 120000
rect 84842 119200 84898 120000
rect 86314 119200 86370 120000
rect 87786 119200 87842 120000
rect 89258 119200 89314 120000
rect 90730 119200 90786 120000
rect 92202 119200 92258 120000
rect 93674 119200 93730 120000
rect 95146 119200 95202 120000
rect 96618 119200 96674 120000
rect 98090 119200 98146 120000
rect 99562 119200 99618 120000
rect 101034 119200 101090 120000
rect 102506 119200 102562 120000
rect 103978 119200 104034 120000
rect 105450 119200 105506 120000
rect 106922 119200 106978 120000
rect 108394 119200 108450 120000
rect 109958 119200 110014 120000
rect 111430 119200 111486 120000
rect 112902 119200 112958 120000
rect 114374 119200 114430 120000
rect 115846 119200 115902 120000
rect 117318 119200 117374 120000
rect 118790 119200 118846 120000
rect 120262 119200 120318 120000
rect 121734 119200 121790 120000
rect 123206 119200 123262 120000
rect 124678 119200 124734 120000
rect 126150 119200 126206 120000
rect 127622 119200 127678 120000
rect 129094 119200 129150 120000
rect 130566 119200 130622 120000
rect 132038 119200 132094 120000
rect 133510 119200 133566 120000
rect 134982 119200 135038 120000
rect 136454 119200 136510 120000
rect 137926 119200 137982 120000
rect 139398 119200 139454 120000
rect 140870 119200 140926 120000
rect 142342 119200 142398 120000
rect 143814 119200 143870 120000
rect 145378 119200 145434 120000
rect 146850 119200 146906 120000
rect 148322 119200 148378 120000
rect 149794 119200 149850 120000
rect 151266 119200 151322 120000
rect 152738 119200 152794 120000
rect 154210 119200 154266 120000
rect 155682 119200 155738 120000
rect 157154 119200 157210 120000
rect 158626 119200 158682 120000
rect 160098 119200 160154 120000
rect 161570 119200 161626 120000
rect 163042 119200 163098 120000
rect 164514 119200 164570 120000
rect 165986 119200 166042 120000
rect 167458 119200 167514 120000
rect 168930 119200 168986 120000
rect 170402 119200 170458 120000
rect 171874 119200 171930 120000
rect 173346 119200 173402 120000
rect 174818 119200 174874 120000
rect 176290 119200 176346 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5906 0 5962 800
rect 7562 0 7618 800
rect 9310 0 9366 800
rect 10966 0 11022 800
rect 12714 0 12770 800
rect 14370 0 14426 800
rect 16118 0 16174 800
rect 17774 0 17830 800
rect 19522 0 19578 800
rect 21178 0 21234 800
rect 22926 0 22982 800
rect 24582 0 24638 800
rect 26238 0 26294 800
rect 27986 0 28042 800
rect 29642 0 29698 800
rect 31390 0 31446 800
rect 33046 0 33102 800
rect 34794 0 34850 800
rect 36450 0 36506 800
rect 38198 0 38254 800
rect 39854 0 39910 800
rect 41602 0 41658 800
rect 43258 0 43314 800
rect 45006 0 45062 800
rect 46662 0 46718 800
rect 48318 0 48374 800
rect 50066 0 50122 800
rect 51722 0 51778 800
rect 53470 0 53526 800
rect 55126 0 55182 800
rect 56874 0 56930 800
rect 58530 0 58586 800
rect 60278 0 60334 800
rect 61934 0 61990 800
rect 63682 0 63738 800
rect 65338 0 65394 800
rect 67086 0 67142 800
rect 68742 0 68798 800
rect 70398 0 70454 800
rect 72146 0 72202 800
rect 73802 0 73858 800
rect 75550 0 75606 800
rect 77206 0 77262 800
rect 78954 0 79010 800
rect 80610 0 80666 800
rect 82358 0 82414 800
rect 84014 0 84070 800
rect 85762 0 85818 800
rect 87418 0 87474 800
rect 89166 0 89222 800
rect 90822 0 90878 800
rect 92478 0 92534 800
rect 94226 0 94282 800
rect 95882 0 95938 800
rect 97630 0 97686 800
rect 99286 0 99342 800
rect 101034 0 101090 800
rect 102690 0 102746 800
rect 104438 0 104494 800
rect 106094 0 106150 800
rect 107842 0 107898 800
rect 109498 0 109554 800
rect 111246 0 111302 800
rect 112902 0 112958 800
rect 114558 0 114614 800
rect 116306 0 116362 800
rect 117962 0 118018 800
rect 119710 0 119766 800
rect 121366 0 121422 800
rect 123114 0 123170 800
rect 124770 0 124826 800
rect 126518 0 126574 800
rect 128174 0 128230 800
rect 129922 0 129978 800
rect 131578 0 131634 800
rect 133326 0 133382 800
rect 134982 0 135038 800
rect 136638 0 136694 800
rect 138386 0 138442 800
rect 140042 0 140098 800
rect 141790 0 141846 800
rect 143446 0 143502 800
rect 145194 0 145250 800
rect 146850 0 146906 800
rect 148598 0 148654 800
rect 150254 0 150310 800
rect 152002 0 152058 800
rect 153658 0 153714 800
rect 155406 0 155462 800
rect 157062 0 157118 800
rect 158718 0 158774 800
rect 160466 0 160522 800
rect 162122 0 162178 800
rect 163870 0 163926 800
rect 165526 0 165582 800
rect 167274 0 167330 800
rect 168930 0 168986 800
rect 170678 0 170734 800
rect 172334 0 172390 800
rect 174082 0 174138 800
rect 175738 0 175794 800
rect 177486 0 177542 800
rect 179142 0 179198 800
<< obsm2 >>
rect 866 119144 2170 119377
rect 2338 119144 3642 119377
rect 3810 119144 5114 119377
rect 5282 119144 6586 119377
rect 6754 119144 8058 119377
rect 8226 119144 9530 119377
rect 9698 119144 11002 119377
rect 11170 119144 12474 119377
rect 12642 119144 13946 119377
rect 14114 119144 15418 119377
rect 15586 119144 16890 119377
rect 17058 119144 18362 119377
rect 18530 119144 19834 119377
rect 20002 119144 21306 119377
rect 21474 119144 22778 119377
rect 22946 119144 24250 119377
rect 24418 119144 25722 119377
rect 25890 119144 27194 119377
rect 27362 119144 28666 119377
rect 28834 119144 30138 119377
rect 30306 119144 31610 119377
rect 31778 119144 33082 119377
rect 33250 119144 34554 119377
rect 34722 119144 36026 119377
rect 36194 119144 37590 119377
rect 37758 119144 39062 119377
rect 39230 119144 40534 119377
rect 40702 119144 42006 119377
rect 42174 119144 43478 119377
rect 43646 119144 44950 119377
rect 45118 119144 46422 119377
rect 46590 119144 47894 119377
rect 48062 119144 49366 119377
rect 49534 119144 50838 119377
rect 51006 119144 52310 119377
rect 52478 119144 53782 119377
rect 53950 119144 55254 119377
rect 55422 119144 56726 119377
rect 56894 119144 58198 119377
rect 58366 119144 59670 119377
rect 59838 119144 61142 119377
rect 61310 119144 62614 119377
rect 62782 119144 64086 119377
rect 64254 119144 65558 119377
rect 65726 119144 67030 119377
rect 67198 119144 68502 119377
rect 68670 119144 69974 119377
rect 70142 119144 71446 119377
rect 71614 119144 73010 119377
rect 73178 119144 74482 119377
rect 74650 119144 75954 119377
rect 76122 119144 77426 119377
rect 77594 119144 78898 119377
rect 79066 119144 80370 119377
rect 80538 119144 81842 119377
rect 82010 119144 83314 119377
rect 83482 119144 84786 119377
rect 84954 119144 86258 119377
rect 86426 119144 87730 119377
rect 87898 119144 89202 119377
rect 89370 119144 90674 119377
rect 90842 119144 92146 119377
rect 92314 119144 93618 119377
rect 93786 119144 95090 119377
rect 95258 119144 96562 119377
rect 96730 119144 98034 119377
rect 98202 119144 99506 119377
rect 99674 119144 100978 119377
rect 101146 119144 102450 119377
rect 102618 119144 103922 119377
rect 104090 119144 105394 119377
rect 105562 119144 106866 119377
rect 107034 119144 108338 119377
rect 108506 119144 109902 119377
rect 110070 119144 111374 119377
rect 111542 119144 112846 119377
rect 113014 119144 114318 119377
rect 114486 119144 115790 119377
rect 115958 119144 117262 119377
rect 117430 119144 118734 119377
rect 118902 119144 120206 119377
rect 120374 119144 121678 119377
rect 121846 119144 123150 119377
rect 123318 119144 124622 119377
rect 124790 119144 126094 119377
rect 126262 119144 127566 119377
rect 127734 119144 129038 119377
rect 129206 119144 130510 119377
rect 130678 119144 131982 119377
rect 132150 119144 133454 119377
rect 133622 119144 134926 119377
rect 135094 119144 136398 119377
rect 136566 119144 137870 119377
rect 138038 119144 139342 119377
rect 139510 119144 140814 119377
rect 140982 119144 142286 119377
rect 142454 119144 143758 119377
rect 143926 119144 145322 119377
rect 145490 119144 146794 119377
rect 146962 119144 148266 119377
rect 148434 119144 149738 119377
rect 149906 119144 151210 119377
rect 151378 119144 152682 119377
rect 152850 119144 154154 119377
rect 154322 119144 155626 119377
rect 155794 119144 157098 119377
rect 157266 119144 158570 119377
rect 158738 119144 160042 119377
rect 160210 119144 161514 119377
rect 161682 119144 162986 119377
rect 163154 119144 164458 119377
rect 164626 119144 165930 119377
rect 166098 119144 167402 119377
rect 167570 119144 168874 119377
rect 169042 119144 170346 119377
rect 170514 119144 171818 119377
rect 171986 119144 173290 119377
rect 173458 119144 174762 119377
rect 174930 119144 176234 119377
rect 176402 119144 177706 119377
rect 177874 119144 179178 119377
rect 756 856 179288 119144
rect 756 206 790 856
rect 958 206 2446 856
rect 2614 206 4102 856
rect 4270 206 5850 856
rect 6018 206 7506 856
rect 7674 206 9254 856
rect 9422 206 10910 856
rect 11078 206 12658 856
rect 12826 206 14314 856
rect 14482 206 16062 856
rect 16230 206 17718 856
rect 17886 206 19466 856
rect 19634 206 21122 856
rect 21290 206 22870 856
rect 23038 206 24526 856
rect 24694 206 26182 856
rect 26350 206 27930 856
rect 28098 206 29586 856
rect 29754 206 31334 856
rect 31502 206 32990 856
rect 33158 206 34738 856
rect 34906 206 36394 856
rect 36562 206 38142 856
rect 38310 206 39798 856
rect 39966 206 41546 856
rect 41714 206 43202 856
rect 43370 206 44950 856
rect 45118 206 46606 856
rect 46774 206 48262 856
rect 48430 206 50010 856
rect 50178 206 51666 856
rect 51834 206 53414 856
rect 53582 206 55070 856
rect 55238 206 56818 856
rect 56986 206 58474 856
rect 58642 206 60222 856
rect 60390 206 61878 856
rect 62046 206 63626 856
rect 63794 206 65282 856
rect 65450 206 67030 856
rect 67198 206 68686 856
rect 68854 206 70342 856
rect 70510 206 72090 856
rect 72258 206 73746 856
rect 73914 206 75494 856
rect 75662 206 77150 856
rect 77318 206 78898 856
rect 79066 206 80554 856
rect 80722 206 82302 856
rect 82470 206 83958 856
rect 84126 206 85706 856
rect 85874 206 87362 856
rect 87530 206 89110 856
rect 89278 206 90766 856
rect 90934 206 92422 856
rect 92590 206 94170 856
rect 94338 206 95826 856
rect 95994 206 97574 856
rect 97742 206 99230 856
rect 99398 206 100978 856
rect 101146 206 102634 856
rect 102802 206 104382 856
rect 104550 206 106038 856
rect 106206 206 107786 856
rect 107954 206 109442 856
rect 109610 206 111190 856
rect 111358 206 112846 856
rect 113014 206 114502 856
rect 114670 206 116250 856
rect 116418 206 117906 856
rect 118074 206 119654 856
rect 119822 206 121310 856
rect 121478 206 123058 856
rect 123226 206 124714 856
rect 124882 206 126462 856
rect 126630 206 128118 856
rect 128286 206 129866 856
rect 130034 206 131522 856
rect 131690 206 133270 856
rect 133438 206 134926 856
rect 135094 206 136582 856
rect 136750 206 138330 856
rect 138498 206 139986 856
rect 140154 206 141734 856
rect 141902 206 143390 856
rect 143558 206 145138 856
rect 145306 206 146794 856
rect 146962 206 148542 856
rect 148710 206 150198 856
rect 150366 206 151946 856
rect 152114 206 153602 856
rect 153770 206 155350 856
rect 155518 206 157006 856
rect 157174 206 158662 856
rect 158830 206 160410 856
rect 160578 206 162066 856
rect 162234 206 163814 856
rect 163982 206 165470 856
rect 165638 206 167218 856
rect 167386 206 168874 856
rect 169042 206 170622 856
rect 170790 206 172278 856
rect 172446 206 174026 856
rect 174194 206 175682 856
rect 175850 206 177430 856
rect 177598 206 179086 856
rect 179254 206 179288 856
<< metal3 >>
rect 0 119280 800 119400
rect 179200 119280 180000 119400
rect 0 118328 800 118448
rect 179200 118192 180000 118312
rect 0 117376 800 117496
rect 179200 117104 180000 117224
rect 0 116424 800 116544
rect 179200 116016 180000 116136
rect 0 115336 800 115456
rect 179200 114928 180000 115048
rect 0 114384 800 114504
rect 179200 113840 180000 113960
rect 0 113432 800 113552
rect 179200 112752 180000 112872
rect 0 112480 800 112600
rect 179200 111664 180000 111784
rect 0 111392 800 111512
rect 0 110440 800 110560
rect 179200 110576 180000 110696
rect 0 109488 800 109608
rect 179200 109488 180000 109608
rect 0 108536 800 108656
rect 179200 108400 180000 108520
rect 0 107584 800 107704
rect 179200 107312 180000 107432
rect 0 106496 800 106616
rect 179200 106224 180000 106344
rect 0 105544 800 105664
rect 179200 105136 180000 105256
rect 0 104592 800 104712
rect 179200 104048 180000 104168
rect 0 103640 800 103760
rect 179200 102960 180000 103080
rect 0 102552 800 102672
rect 179200 101872 180000 101992
rect 0 101600 800 101720
rect 0 100648 800 100768
rect 179200 100784 180000 100904
rect 0 99696 800 99816
rect 179200 99696 180000 99816
rect 0 98608 800 98728
rect 179200 98608 180000 98728
rect 0 97656 800 97776
rect 179200 97520 180000 97640
rect 0 96704 800 96824
rect 179200 96432 180000 96552
rect 0 95752 800 95872
rect 179200 95344 180000 95464
rect 0 94800 800 94920
rect 179200 94256 180000 94376
rect 0 93712 800 93832
rect 179200 93168 180000 93288
rect 0 92760 800 92880
rect 179200 92080 180000 92200
rect 0 91808 800 91928
rect 0 90856 800 90976
rect 179200 90992 180000 91112
rect 0 89768 800 89888
rect 179200 89904 180000 90024
rect 0 88816 800 88936
rect 179200 88816 180000 88936
rect 0 87864 800 87984
rect 179200 87728 180000 87848
rect 0 86912 800 87032
rect 179200 86640 180000 86760
rect 0 85824 800 85944
rect 179200 85552 180000 85672
rect 0 84872 800 84992
rect 179200 84464 180000 84584
rect 0 83920 800 84040
rect 179200 83376 180000 83496
rect 0 82968 800 83088
rect 179200 82288 180000 82408
rect 0 82016 800 82136
rect 179200 81200 180000 81320
rect 0 80928 800 81048
rect 0 79976 800 80096
rect 179200 80112 180000 80232
rect 0 79024 800 79144
rect 179200 79024 180000 79144
rect 0 78072 800 78192
rect 179200 77936 180000 78056
rect 0 76984 800 77104
rect 179200 76848 180000 76968
rect 0 76032 800 76152
rect 179200 75760 180000 75880
rect 0 75080 800 75200
rect 179200 74672 180000 74792
rect 0 74128 800 74248
rect 179200 73584 180000 73704
rect 0 73040 800 73160
rect 179200 72496 180000 72616
rect 0 72088 800 72208
rect 179200 71408 180000 71528
rect 0 71136 800 71256
rect 0 70184 800 70304
rect 179200 70320 180000 70440
rect 0 69232 800 69352
rect 179200 69232 180000 69352
rect 0 68144 800 68264
rect 179200 68144 180000 68264
rect 0 67192 800 67312
rect 179200 67056 180000 67176
rect 0 66240 800 66360
rect 179200 65968 180000 66088
rect 0 65288 800 65408
rect 179200 64880 180000 65000
rect 0 64200 800 64320
rect 179200 63792 180000 63912
rect 0 63248 800 63368
rect 179200 62704 180000 62824
rect 0 62296 800 62416
rect 179200 61616 180000 61736
rect 0 61344 800 61464
rect 0 60392 800 60512
rect 179200 60528 180000 60648
rect 0 59304 800 59424
rect 179200 59304 180000 59424
rect 0 58352 800 58472
rect 179200 58216 180000 58336
rect 0 57400 800 57520
rect 179200 57128 180000 57248
rect 0 56448 800 56568
rect 179200 56040 180000 56160
rect 0 55360 800 55480
rect 179200 54952 180000 55072
rect 0 54408 800 54528
rect 179200 53864 180000 53984
rect 0 53456 800 53576
rect 179200 52776 180000 52896
rect 0 52504 800 52624
rect 179200 51688 180000 51808
rect 0 51416 800 51536
rect 0 50464 800 50584
rect 179200 50600 180000 50720
rect 0 49512 800 49632
rect 179200 49512 180000 49632
rect 0 48560 800 48680
rect 179200 48424 180000 48544
rect 0 47608 800 47728
rect 179200 47336 180000 47456
rect 0 46520 800 46640
rect 179200 46248 180000 46368
rect 0 45568 800 45688
rect 179200 45160 180000 45280
rect 0 44616 800 44736
rect 179200 44072 180000 44192
rect 0 43664 800 43784
rect 179200 42984 180000 43104
rect 0 42576 800 42696
rect 179200 41896 180000 42016
rect 0 41624 800 41744
rect 0 40672 800 40792
rect 179200 40808 180000 40928
rect 0 39720 800 39840
rect 179200 39720 180000 39840
rect 0 38632 800 38752
rect 179200 38632 180000 38752
rect 0 37680 800 37800
rect 179200 37544 180000 37664
rect 0 36728 800 36848
rect 179200 36456 180000 36576
rect 0 35776 800 35896
rect 179200 35368 180000 35488
rect 0 34824 800 34944
rect 179200 34280 180000 34400
rect 0 33736 800 33856
rect 179200 33192 180000 33312
rect 0 32784 800 32904
rect 179200 32104 180000 32224
rect 0 31832 800 31952
rect 0 30880 800 31000
rect 179200 31016 180000 31136
rect 0 29792 800 29912
rect 179200 29928 180000 30048
rect 0 28840 800 28960
rect 179200 28840 180000 28960
rect 0 27888 800 28008
rect 179200 27752 180000 27872
rect 0 26936 800 27056
rect 179200 26664 180000 26784
rect 0 25848 800 25968
rect 179200 25576 180000 25696
rect 0 24896 800 25016
rect 179200 24488 180000 24608
rect 0 23944 800 24064
rect 179200 23400 180000 23520
rect 0 22992 800 23112
rect 179200 22312 180000 22432
rect 0 22040 800 22160
rect 179200 21224 180000 21344
rect 0 20952 800 21072
rect 0 20000 800 20120
rect 179200 20136 180000 20256
rect 0 19048 800 19168
rect 179200 19048 180000 19168
rect 0 18096 800 18216
rect 179200 17960 180000 18080
rect 0 17008 800 17128
rect 179200 16872 180000 16992
rect 0 16056 800 16176
rect 179200 15784 180000 15904
rect 0 15104 800 15224
rect 179200 14696 180000 14816
rect 0 14152 800 14272
rect 179200 13608 180000 13728
rect 0 13064 800 13184
rect 179200 12520 180000 12640
rect 0 12112 800 12232
rect 179200 11432 180000 11552
rect 0 11160 800 11280
rect 0 10208 800 10328
rect 179200 10344 180000 10464
rect 0 9256 800 9376
rect 179200 9256 180000 9376
rect 0 8168 800 8288
rect 179200 8168 180000 8288
rect 0 7216 800 7336
rect 179200 7080 180000 7200
rect 0 6264 800 6384
rect 179200 5992 180000 6112
rect 0 5312 800 5432
rect 179200 4904 180000 5024
rect 0 4224 800 4344
rect 179200 3816 180000 3936
rect 0 3272 800 3392
rect 179200 2728 180000 2848
rect 0 2320 800 2440
rect 179200 1640 180000 1760
rect 0 1368 800 1488
rect 0 416 800 536
rect 179200 552 180000 672
<< obsm3 >>
rect 880 119200 179120 119373
rect 800 118528 179200 119200
rect 880 118392 179200 118528
rect 880 118248 179120 118392
rect 800 118112 179120 118248
rect 800 117576 179200 118112
rect 880 117304 179200 117576
rect 880 117296 179120 117304
rect 800 117024 179120 117296
rect 800 116624 179200 117024
rect 880 116344 179200 116624
rect 800 116216 179200 116344
rect 800 115936 179120 116216
rect 800 115536 179200 115936
rect 880 115256 179200 115536
rect 800 115128 179200 115256
rect 800 114848 179120 115128
rect 800 114584 179200 114848
rect 880 114304 179200 114584
rect 800 114040 179200 114304
rect 800 113760 179120 114040
rect 800 113632 179200 113760
rect 880 113352 179200 113632
rect 800 112952 179200 113352
rect 800 112680 179120 112952
rect 880 112672 179120 112680
rect 880 112400 179200 112672
rect 800 111864 179200 112400
rect 800 111592 179120 111864
rect 880 111584 179120 111592
rect 880 111312 179200 111584
rect 800 110776 179200 111312
rect 800 110640 179120 110776
rect 880 110496 179120 110640
rect 880 110360 179200 110496
rect 800 109688 179200 110360
rect 880 109408 179120 109688
rect 800 108736 179200 109408
rect 880 108600 179200 108736
rect 880 108456 179120 108600
rect 800 108320 179120 108456
rect 800 107784 179200 108320
rect 880 107512 179200 107784
rect 880 107504 179120 107512
rect 800 107232 179120 107504
rect 800 106696 179200 107232
rect 880 106424 179200 106696
rect 880 106416 179120 106424
rect 800 106144 179120 106416
rect 800 105744 179200 106144
rect 880 105464 179200 105744
rect 800 105336 179200 105464
rect 800 105056 179120 105336
rect 800 104792 179200 105056
rect 880 104512 179200 104792
rect 800 104248 179200 104512
rect 800 103968 179120 104248
rect 800 103840 179200 103968
rect 880 103560 179200 103840
rect 800 103160 179200 103560
rect 800 102880 179120 103160
rect 800 102752 179200 102880
rect 880 102472 179200 102752
rect 800 102072 179200 102472
rect 800 101800 179120 102072
rect 880 101792 179120 101800
rect 880 101520 179200 101792
rect 800 100984 179200 101520
rect 800 100848 179120 100984
rect 880 100704 179120 100848
rect 880 100568 179200 100704
rect 800 99896 179200 100568
rect 880 99616 179120 99896
rect 800 98808 179200 99616
rect 880 98528 179120 98808
rect 800 97856 179200 98528
rect 880 97720 179200 97856
rect 880 97576 179120 97720
rect 800 97440 179120 97576
rect 800 96904 179200 97440
rect 880 96632 179200 96904
rect 880 96624 179120 96632
rect 800 96352 179120 96624
rect 800 95952 179200 96352
rect 880 95672 179200 95952
rect 800 95544 179200 95672
rect 800 95264 179120 95544
rect 800 95000 179200 95264
rect 880 94720 179200 95000
rect 800 94456 179200 94720
rect 800 94176 179120 94456
rect 800 93912 179200 94176
rect 880 93632 179200 93912
rect 800 93368 179200 93632
rect 800 93088 179120 93368
rect 800 92960 179200 93088
rect 880 92680 179200 92960
rect 800 92280 179200 92680
rect 800 92008 179120 92280
rect 880 92000 179120 92008
rect 880 91728 179200 92000
rect 800 91192 179200 91728
rect 800 91056 179120 91192
rect 880 90912 179120 91056
rect 880 90776 179200 90912
rect 800 90104 179200 90776
rect 800 89968 179120 90104
rect 880 89824 179120 89968
rect 880 89688 179200 89824
rect 800 89016 179200 89688
rect 880 88736 179120 89016
rect 800 88064 179200 88736
rect 880 87928 179200 88064
rect 880 87784 179120 87928
rect 800 87648 179120 87784
rect 800 87112 179200 87648
rect 880 86840 179200 87112
rect 880 86832 179120 86840
rect 800 86560 179120 86832
rect 800 86024 179200 86560
rect 880 85752 179200 86024
rect 880 85744 179120 85752
rect 800 85472 179120 85744
rect 800 85072 179200 85472
rect 880 84792 179200 85072
rect 800 84664 179200 84792
rect 800 84384 179120 84664
rect 800 84120 179200 84384
rect 880 83840 179200 84120
rect 800 83576 179200 83840
rect 800 83296 179120 83576
rect 800 83168 179200 83296
rect 880 82888 179200 83168
rect 800 82488 179200 82888
rect 800 82216 179120 82488
rect 880 82208 179120 82216
rect 880 81936 179200 82208
rect 800 81400 179200 81936
rect 800 81128 179120 81400
rect 880 81120 179120 81128
rect 880 80848 179200 81120
rect 800 80312 179200 80848
rect 800 80176 179120 80312
rect 880 80032 179120 80176
rect 880 79896 179200 80032
rect 800 79224 179200 79896
rect 880 78944 179120 79224
rect 800 78272 179200 78944
rect 880 78136 179200 78272
rect 880 77992 179120 78136
rect 800 77856 179120 77992
rect 800 77184 179200 77856
rect 880 77048 179200 77184
rect 880 76904 179120 77048
rect 800 76768 179120 76904
rect 800 76232 179200 76768
rect 880 75960 179200 76232
rect 880 75952 179120 75960
rect 800 75680 179120 75952
rect 800 75280 179200 75680
rect 880 75000 179200 75280
rect 800 74872 179200 75000
rect 800 74592 179120 74872
rect 800 74328 179200 74592
rect 880 74048 179200 74328
rect 800 73784 179200 74048
rect 800 73504 179120 73784
rect 800 73240 179200 73504
rect 880 72960 179200 73240
rect 800 72696 179200 72960
rect 800 72416 179120 72696
rect 800 72288 179200 72416
rect 880 72008 179200 72288
rect 800 71608 179200 72008
rect 800 71336 179120 71608
rect 880 71328 179120 71336
rect 880 71056 179200 71328
rect 800 70520 179200 71056
rect 800 70384 179120 70520
rect 880 70240 179120 70384
rect 880 70104 179200 70240
rect 800 69432 179200 70104
rect 880 69152 179120 69432
rect 800 68344 179200 69152
rect 880 68064 179120 68344
rect 800 67392 179200 68064
rect 880 67256 179200 67392
rect 880 67112 179120 67256
rect 800 66976 179120 67112
rect 800 66440 179200 66976
rect 880 66168 179200 66440
rect 880 66160 179120 66168
rect 800 65888 179120 66160
rect 800 65488 179200 65888
rect 880 65208 179200 65488
rect 800 65080 179200 65208
rect 800 64800 179120 65080
rect 800 64400 179200 64800
rect 880 64120 179200 64400
rect 800 63992 179200 64120
rect 800 63712 179120 63992
rect 800 63448 179200 63712
rect 880 63168 179200 63448
rect 800 62904 179200 63168
rect 800 62624 179120 62904
rect 800 62496 179200 62624
rect 880 62216 179200 62496
rect 800 61816 179200 62216
rect 800 61544 179120 61816
rect 880 61536 179120 61544
rect 880 61264 179200 61536
rect 800 60728 179200 61264
rect 800 60592 179120 60728
rect 880 60448 179120 60592
rect 880 60312 179200 60448
rect 800 59504 179200 60312
rect 880 59224 179120 59504
rect 800 58552 179200 59224
rect 880 58416 179200 58552
rect 880 58272 179120 58416
rect 800 58136 179120 58272
rect 800 57600 179200 58136
rect 880 57328 179200 57600
rect 880 57320 179120 57328
rect 800 57048 179120 57320
rect 800 56648 179200 57048
rect 880 56368 179200 56648
rect 800 56240 179200 56368
rect 800 55960 179120 56240
rect 800 55560 179200 55960
rect 880 55280 179200 55560
rect 800 55152 179200 55280
rect 800 54872 179120 55152
rect 800 54608 179200 54872
rect 880 54328 179200 54608
rect 800 54064 179200 54328
rect 800 53784 179120 54064
rect 800 53656 179200 53784
rect 880 53376 179200 53656
rect 800 52976 179200 53376
rect 800 52704 179120 52976
rect 880 52696 179120 52704
rect 880 52424 179200 52696
rect 800 51888 179200 52424
rect 800 51616 179120 51888
rect 880 51608 179120 51616
rect 880 51336 179200 51608
rect 800 50800 179200 51336
rect 800 50664 179120 50800
rect 880 50520 179120 50664
rect 880 50384 179200 50520
rect 800 49712 179200 50384
rect 880 49432 179120 49712
rect 800 48760 179200 49432
rect 880 48624 179200 48760
rect 880 48480 179120 48624
rect 800 48344 179120 48480
rect 800 47808 179200 48344
rect 880 47536 179200 47808
rect 880 47528 179120 47536
rect 800 47256 179120 47528
rect 800 46720 179200 47256
rect 880 46448 179200 46720
rect 880 46440 179120 46448
rect 800 46168 179120 46440
rect 800 45768 179200 46168
rect 880 45488 179200 45768
rect 800 45360 179200 45488
rect 800 45080 179120 45360
rect 800 44816 179200 45080
rect 880 44536 179200 44816
rect 800 44272 179200 44536
rect 800 43992 179120 44272
rect 800 43864 179200 43992
rect 880 43584 179200 43864
rect 800 43184 179200 43584
rect 800 42904 179120 43184
rect 800 42776 179200 42904
rect 880 42496 179200 42776
rect 800 42096 179200 42496
rect 800 41824 179120 42096
rect 880 41816 179120 41824
rect 880 41544 179200 41816
rect 800 41008 179200 41544
rect 800 40872 179120 41008
rect 880 40728 179120 40872
rect 880 40592 179200 40728
rect 800 39920 179200 40592
rect 880 39640 179120 39920
rect 800 38832 179200 39640
rect 880 38552 179120 38832
rect 800 37880 179200 38552
rect 880 37744 179200 37880
rect 880 37600 179120 37744
rect 800 37464 179120 37600
rect 800 36928 179200 37464
rect 880 36656 179200 36928
rect 880 36648 179120 36656
rect 800 36376 179120 36648
rect 800 35976 179200 36376
rect 880 35696 179200 35976
rect 800 35568 179200 35696
rect 800 35288 179120 35568
rect 800 35024 179200 35288
rect 880 34744 179200 35024
rect 800 34480 179200 34744
rect 800 34200 179120 34480
rect 800 33936 179200 34200
rect 880 33656 179200 33936
rect 800 33392 179200 33656
rect 800 33112 179120 33392
rect 800 32984 179200 33112
rect 880 32704 179200 32984
rect 800 32304 179200 32704
rect 800 32032 179120 32304
rect 880 32024 179120 32032
rect 880 31752 179200 32024
rect 800 31216 179200 31752
rect 800 31080 179120 31216
rect 880 30936 179120 31080
rect 880 30800 179200 30936
rect 800 30128 179200 30800
rect 800 29992 179120 30128
rect 880 29848 179120 29992
rect 880 29712 179200 29848
rect 800 29040 179200 29712
rect 880 28760 179120 29040
rect 800 28088 179200 28760
rect 880 27952 179200 28088
rect 880 27808 179120 27952
rect 800 27672 179120 27808
rect 800 27136 179200 27672
rect 880 26864 179200 27136
rect 880 26856 179120 26864
rect 800 26584 179120 26856
rect 800 26048 179200 26584
rect 880 25776 179200 26048
rect 880 25768 179120 25776
rect 800 25496 179120 25768
rect 800 25096 179200 25496
rect 880 24816 179200 25096
rect 800 24688 179200 24816
rect 800 24408 179120 24688
rect 800 24144 179200 24408
rect 880 23864 179200 24144
rect 800 23600 179200 23864
rect 800 23320 179120 23600
rect 800 23192 179200 23320
rect 880 22912 179200 23192
rect 800 22512 179200 22912
rect 800 22240 179120 22512
rect 880 22232 179120 22240
rect 880 21960 179200 22232
rect 800 21424 179200 21960
rect 800 21152 179120 21424
rect 880 21144 179120 21152
rect 880 20872 179200 21144
rect 800 20336 179200 20872
rect 800 20200 179120 20336
rect 880 20056 179120 20200
rect 880 19920 179200 20056
rect 800 19248 179200 19920
rect 880 18968 179120 19248
rect 800 18296 179200 18968
rect 880 18160 179200 18296
rect 880 18016 179120 18160
rect 800 17880 179120 18016
rect 800 17208 179200 17880
rect 880 17072 179200 17208
rect 880 16928 179120 17072
rect 800 16792 179120 16928
rect 800 16256 179200 16792
rect 880 15984 179200 16256
rect 880 15976 179120 15984
rect 800 15704 179120 15976
rect 800 15304 179200 15704
rect 880 15024 179200 15304
rect 800 14896 179200 15024
rect 800 14616 179120 14896
rect 800 14352 179200 14616
rect 880 14072 179200 14352
rect 800 13808 179200 14072
rect 800 13528 179120 13808
rect 800 13264 179200 13528
rect 880 12984 179200 13264
rect 800 12720 179200 12984
rect 800 12440 179120 12720
rect 800 12312 179200 12440
rect 880 12032 179200 12312
rect 800 11632 179200 12032
rect 800 11360 179120 11632
rect 880 11352 179120 11360
rect 880 11080 179200 11352
rect 800 10544 179200 11080
rect 800 10408 179120 10544
rect 880 10264 179120 10408
rect 880 10128 179200 10264
rect 800 9456 179200 10128
rect 880 9176 179120 9456
rect 800 8368 179200 9176
rect 880 8088 179120 8368
rect 800 7416 179200 8088
rect 880 7280 179200 7416
rect 880 7136 179120 7280
rect 800 7000 179120 7136
rect 800 6464 179200 7000
rect 880 6192 179200 6464
rect 880 6184 179120 6192
rect 800 5912 179120 6184
rect 800 5512 179200 5912
rect 880 5232 179200 5512
rect 800 5104 179200 5232
rect 800 4824 179120 5104
rect 800 4424 179200 4824
rect 880 4144 179200 4424
rect 800 4016 179200 4144
rect 800 3736 179120 4016
rect 800 3472 179200 3736
rect 880 3192 179200 3472
rect 800 2928 179200 3192
rect 800 2648 179120 2928
rect 800 2520 179200 2648
rect 880 2240 179200 2520
rect 800 1840 179200 2240
rect 800 1568 179120 1840
rect 880 1560 179120 1568
rect 880 1288 179200 1560
rect 800 752 179200 1288
rect 800 616 179120 752
rect 880 472 179120 616
rect 880 443 179200 472
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 76419 6427 80928 10437
rect 81408 6427 81588 10437
rect 82068 6427 82248 10437
rect 82728 6427 82908 10437
rect 83388 6427 86605 10437
<< labels >>
rlabel metal3 s 179200 11432 180000 11552 6 adc0_dat_i[0]
port 1 nsew signal input
rlabel metal3 s 179200 47336 180000 47456 6 adc0_dat_i[10]
port 2 nsew signal input
rlabel metal3 s 179200 50600 180000 50720 6 adc0_dat_i[11]
port 3 nsew signal input
rlabel metal3 s 179200 53864 180000 53984 6 adc0_dat_i[12]
port 4 nsew signal input
rlabel metal3 s 179200 57128 180000 57248 6 adc0_dat_i[13]
port 5 nsew signal input
rlabel metal3 s 179200 60528 180000 60648 6 adc0_dat_i[14]
port 6 nsew signal input
rlabel metal3 s 179200 63792 180000 63912 6 adc0_dat_i[15]
port 7 nsew signal input
rlabel metal3 s 179200 67056 180000 67176 6 adc0_dat_i[16]
port 8 nsew signal input
rlabel metal3 s 179200 70320 180000 70440 6 adc0_dat_i[17]
port 9 nsew signal input
rlabel metal3 s 179200 73584 180000 73704 6 adc0_dat_i[18]
port 10 nsew signal input
rlabel metal3 s 179200 76848 180000 76968 6 adc0_dat_i[19]
port 11 nsew signal input
rlabel metal3 s 179200 15784 180000 15904 6 adc0_dat_i[1]
port 12 nsew signal input
rlabel metal3 s 179200 80112 180000 80232 6 adc0_dat_i[20]
port 13 nsew signal input
rlabel metal3 s 179200 83376 180000 83496 6 adc0_dat_i[21]
port 14 nsew signal input
rlabel metal3 s 179200 86640 180000 86760 6 adc0_dat_i[22]
port 15 nsew signal input
rlabel metal3 s 179200 89904 180000 90024 6 adc0_dat_i[23]
port 16 nsew signal input
rlabel metal3 s 179200 93168 180000 93288 6 adc0_dat_i[24]
port 17 nsew signal input
rlabel metal3 s 179200 96432 180000 96552 6 adc0_dat_i[25]
port 18 nsew signal input
rlabel metal3 s 179200 99696 180000 99816 6 adc0_dat_i[26]
port 19 nsew signal input
rlabel metal3 s 179200 102960 180000 103080 6 adc0_dat_i[27]
port 20 nsew signal input
rlabel metal3 s 179200 106224 180000 106344 6 adc0_dat_i[28]
port 21 nsew signal input
rlabel metal3 s 179200 109488 180000 109608 6 adc0_dat_i[29]
port 22 nsew signal input
rlabel metal3 s 179200 20136 180000 20256 6 adc0_dat_i[2]
port 23 nsew signal input
rlabel metal3 s 179200 112752 180000 112872 6 adc0_dat_i[30]
port 24 nsew signal input
rlabel metal3 s 179200 116016 180000 116136 6 adc0_dat_i[31]
port 25 nsew signal input
rlabel metal3 s 179200 24488 180000 24608 6 adc0_dat_i[3]
port 26 nsew signal input
rlabel metal3 s 179200 27752 180000 27872 6 adc0_dat_i[4]
port 27 nsew signal input
rlabel metal3 s 179200 31016 180000 31136 6 adc0_dat_i[5]
port 28 nsew signal input
rlabel metal3 s 179200 34280 180000 34400 6 adc0_dat_i[6]
port 29 nsew signal input
rlabel metal3 s 179200 37544 180000 37664 6 adc0_dat_i[7]
port 30 nsew signal input
rlabel metal3 s 179200 40808 180000 40928 6 adc0_dat_i[8]
port 31 nsew signal input
rlabel metal3 s 179200 44072 180000 44192 6 adc0_dat_i[9]
port 32 nsew signal input
rlabel metal3 s 179200 12520 180000 12640 6 adc1_dat_i[0]
port 33 nsew signal input
rlabel metal3 s 179200 48424 180000 48544 6 adc1_dat_i[10]
port 34 nsew signal input
rlabel metal3 s 179200 51688 180000 51808 6 adc1_dat_i[11]
port 35 nsew signal input
rlabel metal3 s 179200 54952 180000 55072 6 adc1_dat_i[12]
port 36 nsew signal input
rlabel metal3 s 179200 58216 180000 58336 6 adc1_dat_i[13]
port 37 nsew signal input
rlabel metal3 s 179200 61616 180000 61736 6 adc1_dat_i[14]
port 38 nsew signal input
rlabel metal3 s 179200 64880 180000 65000 6 adc1_dat_i[15]
port 39 nsew signal input
rlabel metal3 s 179200 68144 180000 68264 6 adc1_dat_i[16]
port 40 nsew signal input
rlabel metal3 s 179200 71408 180000 71528 6 adc1_dat_i[17]
port 41 nsew signal input
rlabel metal3 s 179200 74672 180000 74792 6 adc1_dat_i[18]
port 42 nsew signal input
rlabel metal3 s 179200 77936 180000 78056 6 adc1_dat_i[19]
port 43 nsew signal input
rlabel metal3 s 179200 16872 180000 16992 6 adc1_dat_i[1]
port 44 nsew signal input
rlabel metal3 s 179200 81200 180000 81320 6 adc1_dat_i[20]
port 45 nsew signal input
rlabel metal3 s 179200 84464 180000 84584 6 adc1_dat_i[21]
port 46 nsew signal input
rlabel metal3 s 179200 87728 180000 87848 6 adc1_dat_i[22]
port 47 nsew signal input
rlabel metal3 s 179200 90992 180000 91112 6 adc1_dat_i[23]
port 48 nsew signal input
rlabel metal3 s 179200 94256 180000 94376 6 adc1_dat_i[24]
port 49 nsew signal input
rlabel metal3 s 179200 97520 180000 97640 6 adc1_dat_i[25]
port 50 nsew signal input
rlabel metal3 s 179200 100784 180000 100904 6 adc1_dat_i[26]
port 51 nsew signal input
rlabel metal3 s 179200 104048 180000 104168 6 adc1_dat_i[27]
port 52 nsew signal input
rlabel metal3 s 179200 107312 180000 107432 6 adc1_dat_i[28]
port 53 nsew signal input
rlabel metal3 s 179200 110576 180000 110696 6 adc1_dat_i[29]
port 54 nsew signal input
rlabel metal3 s 179200 21224 180000 21344 6 adc1_dat_i[2]
port 55 nsew signal input
rlabel metal3 s 179200 113840 180000 113960 6 adc1_dat_i[30]
port 56 nsew signal input
rlabel metal3 s 179200 117104 180000 117224 6 adc1_dat_i[31]
port 57 nsew signal input
rlabel metal3 s 179200 25576 180000 25696 6 adc1_dat_i[3]
port 58 nsew signal input
rlabel metal3 s 179200 28840 180000 28960 6 adc1_dat_i[4]
port 59 nsew signal input
rlabel metal3 s 179200 32104 180000 32224 6 adc1_dat_i[5]
port 60 nsew signal input
rlabel metal3 s 179200 35368 180000 35488 6 adc1_dat_i[6]
port 61 nsew signal input
rlabel metal3 s 179200 38632 180000 38752 6 adc1_dat_i[7]
port 62 nsew signal input
rlabel metal3 s 179200 41896 180000 42016 6 adc1_dat_i[8]
port 63 nsew signal input
rlabel metal3 s 179200 45160 180000 45280 6 adc1_dat_i[9]
port 64 nsew signal input
rlabel metal3 s 179200 13608 180000 13728 6 adc2_dat_i[0]
port 65 nsew signal input
rlabel metal3 s 179200 49512 180000 49632 6 adc2_dat_i[10]
port 66 nsew signal input
rlabel metal3 s 179200 52776 180000 52896 6 adc2_dat_i[11]
port 67 nsew signal input
rlabel metal3 s 179200 56040 180000 56160 6 adc2_dat_i[12]
port 68 nsew signal input
rlabel metal3 s 179200 59304 180000 59424 6 adc2_dat_i[13]
port 69 nsew signal input
rlabel metal3 s 179200 62704 180000 62824 6 adc2_dat_i[14]
port 70 nsew signal input
rlabel metal3 s 179200 65968 180000 66088 6 adc2_dat_i[15]
port 71 nsew signal input
rlabel metal3 s 179200 69232 180000 69352 6 adc2_dat_i[16]
port 72 nsew signal input
rlabel metal3 s 179200 72496 180000 72616 6 adc2_dat_i[17]
port 73 nsew signal input
rlabel metal3 s 179200 75760 180000 75880 6 adc2_dat_i[18]
port 74 nsew signal input
rlabel metal3 s 179200 79024 180000 79144 6 adc2_dat_i[19]
port 75 nsew signal input
rlabel metal3 s 179200 17960 180000 18080 6 adc2_dat_i[1]
port 76 nsew signal input
rlabel metal3 s 179200 82288 180000 82408 6 adc2_dat_i[20]
port 77 nsew signal input
rlabel metal3 s 179200 85552 180000 85672 6 adc2_dat_i[21]
port 78 nsew signal input
rlabel metal3 s 179200 88816 180000 88936 6 adc2_dat_i[22]
port 79 nsew signal input
rlabel metal3 s 179200 92080 180000 92200 6 adc2_dat_i[23]
port 80 nsew signal input
rlabel metal3 s 179200 95344 180000 95464 6 adc2_dat_i[24]
port 81 nsew signal input
rlabel metal3 s 179200 98608 180000 98728 6 adc2_dat_i[25]
port 82 nsew signal input
rlabel metal3 s 179200 101872 180000 101992 6 adc2_dat_i[26]
port 83 nsew signal input
rlabel metal3 s 179200 105136 180000 105256 6 adc2_dat_i[27]
port 84 nsew signal input
rlabel metal3 s 179200 108400 180000 108520 6 adc2_dat_i[28]
port 85 nsew signal input
rlabel metal3 s 179200 111664 180000 111784 6 adc2_dat_i[29]
port 86 nsew signal input
rlabel metal3 s 179200 22312 180000 22432 6 adc2_dat_i[2]
port 87 nsew signal input
rlabel metal3 s 179200 114928 180000 115048 6 adc2_dat_i[30]
port 88 nsew signal input
rlabel metal3 s 179200 118192 180000 118312 6 adc2_dat_i[31]
port 89 nsew signal input
rlabel metal3 s 179200 26664 180000 26784 6 adc2_dat_i[3]
port 90 nsew signal input
rlabel metal3 s 179200 29928 180000 30048 6 adc2_dat_i[4]
port 91 nsew signal input
rlabel metal3 s 179200 33192 180000 33312 6 adc2_dat_i[5]
port 92 nsew signal input
rlabel metal3 s 179200 36456 180000 36576 6 adc2_dat_i[6]
port 93 nsew signal input
rlabel metal3 s 179200 39720 180000 39840 6 adc2_dat_i[7]
port 94 nsew signal input
rlabel metal3 s 179200 42984 180000 43104 6 adc2_dat_i[8]
port 95 nsew signal input
rlabel metal3 s 179200 46248 180000 46368 6 adc2_dat_i[9]
port 96 nsew signal input
rlabel metal3 s 179200 14696 180000 14816 6 adc_dvalid_i[0]
port 97 nsew signal input
rlabel metal3 s 179200 19048 180000 19168 6 adc_dvalid_i[1]
port 98 nsew signal input
rlabel metal3 s 179200 23400 180000 23520 6 adc_dvalid_i[2]
port 99 nsew signal input
rlabel metal2 s 754 119200 810 120000 6 io_in[0]
port 100 nsew signal input
rlabel metal2 s 45006 119200 45062 120000 6 io_in[10]
port 101 nsew signal input
rlabel metal2 s 49422 119200 49478 120000 6 io_in[11]
port 102 nsew signal input
rlabel metal2 s 53838 119200 53894 120000 6 io_in[12]
port 103 nsew signal input
rlabel metal2 s 58254 119200 58310 120000 6 io_in[13]
port 104 nsew signal input
rlabel metal2 s 62670 119200 62726 120000 6 io_in[14]
port 105 nsew signal input
rlabel metal2 s 67086 119200 67142 120000 6 io_in[15]
port 106 nsew signal input
rlabel metal2 s 71502 119200 71558 120000 6 io_in[16]
port 107 nsew signal input
rlabel metal2 s 76010 119200 76066 120000 6 io_in[17]
port 108 nsew signal input
rlabel metal2 s 80426 119200 80482 120000 6 io_in[18]
port 109 nsew signal input
rlabel metal2 s 84842 119200 84898 120000 6 io_in[19]
port 110 nsew signal input
rlabel metal2 s 5170 119200 5226 120000 6 io_in[1]
port 111 nsew signal input
rlabel metal2 s 89258 119200 89314 120000 6 io_in[20]
port 112 nsew signal input
rlabel metal2 s 93674 119200 93730 120000 6 io_in[21]
port 113 nsew signal input
rlabel metal2 s 98090 119200 98146 120000 6 io_in[22]
port 114 nsew signal input
rlabel metal2 s 102506 119200 102562 120000 6 io_in[23]
port 115 nsew signal input
rlabel metal2 s 106922 119200 106978 120000 6 io_in[24]
port 116 nsew signal input
rlabel metal2 s 111430 119200 111486 120000 6 io_in[25]
port 117 nsew signal input
rlabel metal2 s 115846 119200 115902 120000 6 io_in[26]
port 118 nsew signal input
rlabel metal2 s 120262 119200 120318 120000 6 io_in[27]
port 119 nsew signal input
rlabel metal2 s 124678 119200 124734 120000 6 io_in[28]
port 120 nsew signal input
rlabel metal2 s 129094 119200 129150 120000 6 io_in[29]
port 121 nsew signal input
rlabel metal2 s 9586 119200 9642 120000 6 io_in[2]
port 122 nsew signal input
rlabel metal2 s 133510 119200 133566 120000 6 io_in[30]
port 123 nsew signal input
rlabel metal2 s 137926 119200 137982 120000 6 io_in[31]
port 124 nsew signal input
rlabel metal2 s 142342 119200 142398 120000 6 io_in[32]
port 125 nsew signal input
rlabel metal2 s 146850 119200 146906 120000 6 io_in[33]
port 126 nsew signal input
rlabel metal2 s 151266 119200 151322 120000 6 io_in[34]
port 127 nsew signal input
rlabel metal2 s 155682 119200 155738 120000 6 io_in[35]
port 128 nsew signal input
rlabel metal2 s 160098 119200 160154 120000 6 io_in[36]
port 129 nsew signal input
rlabel metal2 s 164514 119200 164570 120000 6 io_in[37]
port 130 nsew signal input
rlabel metal2 s 14002 119200 14058 120000 6 io_in[3]
port 131 nsew signal input
rlabel metal2 s 18418 119200 18474 120000 6 io_in[4]
port 132 nsew signal input
rlabel metal2 s 22834 119200 22890 120000 6 io_in[5]
port 133 nsew signal input
rlabel metal2 s 27250 119200 27306 120000 6 io_in[6]
port 134 nsew signal input
rlabel metal2 s 31666 119200 31722 120000 6 io_in[7]
port 135 nsew signal input
rlabel metal2 s 36082 119200 36138 120000 6 io_in[8]
port 136 nsew signal input
rlabel metal2 s 40590 119200 40646 120000 6 io_in[9]
port 137 nsew signal input
rlabel metal2 s 2226 119200 2282 120000 6 io_oeb[0]
port 138 nsew signal output
rlabel metal2 s 46478 119200 46534 120000 6 io_oeb[10]
port 139 nsew signal output
rlabel metal2 s 50894 119200 50950 120000 6 io_oeb[11]
port 140 nsew signal output
rlabel metal2 s 55310 119200 55366 120000 6 io_oeb[12]
port 141 nsew signal output
rlabel metal2 s 59726 119200 59782 120000 6 io_oeb[13]
port 142 nsew signal output
rlabel metal2 s 64142 119200 64198 120000 6 io_oeb[14]
port 143 nsew signal output
rlabel metal2 s 68558 119200 68614 120000 6 io_oeb[15]
port 144 nsew signal output
rlabel metal2 s 73066 119200 73122 120000 6 io_oeb[16]
port 145 nsew signal output
rlabel metal2 s 77482 119200 77538 120000 6 io_oeb[17]
port 146 nsew signal output
rlabel metal2 s 81898 119200 81954 120000 6 io_oeb[18]
port 147 nsew signal output
rlabel metal2 s 86314 119200 86370 120000 6 io_oeb[19]
port 148 nsew signal output
rlabel metal2 s 6642 119200 6698 120000 6 io_oeb[1]
port 149 nsew signal output
rlabel metal2 s 90730 119200 90786 120000 6 io_oeb[20]
port 150 nsew signal output
rlabel metal2 s 95146 119200 95202 120000 6 io_oeb[21]
port 151 nsew signal output
rlabel metal2 s 99562 119200 99618 120000 6 io_oeb[22]
port 152 nsew signal output
rlabel metal2 s 103978 119200 104034 120000 6 io_oeb[23]
port 153 nsew signal output
rlabel metal2 s 108394 119200 108450 120000 6 io_oeb[24]
port 154 nsew signal output
rlabel metal2 s 112902 119200 112958 120000 6 io_oeb[25]
port 155 nsew signal output
rlabel metal2 s 117318 119200 117374 120000 6 io_oeb[26]
port 156 nsew signal output
rlabel metal2 s 121734 119200 121790 120000 6 io_oeb[27]
port 157 nsew signal output
rlabel metal2 s 126150 119200 126206 120000 6 io_oeb[28]
port 158 nsew signal output
rlabel metal2 s 130566 119200 130622 120000 6 io_oeb[29]
port 159 nsew signal output
rlabel metal2 s 11058 119200 11114 120000 6 io_oeb[2]
port 160 nsew signal output
rlabel metal2 s 134982 119200 135038 120000 6 io_oeb[30]
port 161 nsew signal output
rlabel metal2 s 139398 119200 139454 120000 6 io_oeb[31]
port 162 nsew signal output
rlabel metal2 s 143814 119200 143870 120000 6 io_oeb[32]
port 163 nsew signal output
rlabel metal2 s 148322 119200 148378 120000 6 io_oeb[33]
port 164 nsew signal output
rlabel metal2 s 152738 119200 152794 120000 6 io_oeb[34]
port 165 nsew signal output
rlabel metal2 s 157154 119200 157210 120000 6 io_oeb[35]
port 166 nsew signal output
rlabel metal2 s 161570 119200 161626 120000 6 io_oeb[36]
port 167 nsew signal output
rlabel metal2 s 165986 119200 166042 120000 6 io_oeb[37]
port 168 nsew signal output
rlabel metal2 s 15474 119200 15530 120000 6 io_oeb[3]
port 169 nsew signal output
rlabel metal2 s 19890 119200 19946 120000 6 io_oeb[4]
port 170 nsew signal output
rlabel metal2 s 24306 119200 24362 120000 6 io_oeb[5]
port 171 nsew signal output
rlabel metal2 s 28722 119200 28778 120000 6 io_oeb[6]
port 172 nsew signal output
rlabel metal2 s 33138 119200 33194 120000 6 io_oeb[7]
port 173 nsew signal output
rlabel metal2 s 37646 119200 37702 120000 6 io_oeb[8]
port 174 nsew signal output
rlabel metal2 s 42062 119200 42118 120000 6 io_oeb[9]
port 175 nsew signal output
rlabel metal2 s 3698 119200 3754 120000 6 io_out[0]
port 176 nsew signal output
rlabel metal2 s 47950 119200 48006 120000 6 io_out[10]
port 177 nsew signal output
rlabel metal2 s 52366 119200 52422 120000 6 io_out[11]
port 178 nsew signal output
rlabel metal2 s 56782 119200 56838 120000 6 io_out[12]
port 179 nsew signal output
rlabel metal2 s 61198 119200 61254 120000 6 io_out[13]
port 180 nsew signal output
rlabel metal2 s 65614 119200 65670 120000 6 io_out[14]
port 181 nsew signal output
rlabel metal2 s 70030 119200 70086 120000 6 io_out[15]
port 182 nsew signal output
rlabel metal2 s 74538 119200 74594 120000 6 io_out[16]
port 183 nsew signal output
rlabel metal2 s 78954 119200 79010 120000 6 io_out[17]
port 184 nsew signal output
rlabel metal2 s 83370 119200 83426 120000 6 io_out[18]
port 185 nsew signal output
rlabel metal2 s 87786 119200 87842 120000 6 io_out[19]
port 186 nsew signal output
rlabel metal2 s 8114 119200 8170 120000 6 io_out[1]
port 187 nsew signal output
rlabel metal2 s 92202 119200 92258 120000 6 io_out[20]
port 188 nsew signal output
rlabel metal2 s 96618 119200 96674 120000 6 io_out[21]
port 189 nsew signal output
rlabel metal2 s 101034 119200 101090 120000 6 io_out[22]
port 190 nsew signal output
rlabel metal2 s 105450 119200 105506 120000 6 io_out[23]
port 191 nsew signal output
rlabel metal2 s 109958 119200 110014 120000 6 io_out[24]
port 192 nsew signal output
rlabel metal2 s 114374 119200 114430 120000 6 io_out[25]
port 193 nsew signal output
rlabel metal2 s 118790 119200 118846 120000 6 io_out[26]
port 194 nsew signal output
rlabel metal2 s 123206 119200 123262 120000 6 io_out[27]
port 195 nsew signal output
rlabel metal2 s 127622 119200 127678 120000 6 io_out[28]
port 196 nsew signal output
rlabel metal2 s 132038 119200 132094 120000 6 io_out[29]
port 197 nsew signal output
rlabel metal2 s 12530 119200 12586 120000 6 io_out[2]
port 198 nsew signal output
rlabel metal2 s 136454 119200 136510 120000 6 io_out[30]
port 199 nsew signal output
rlabel metal2 s 140870 119200 140926 120000 6 io_out[31]
port 200 nsew signal output
rlabel metal2 s 145378 119200 145434 120000 6 io_out[32]
port 201 nsew signal output
rlabel metal2 s 149794 119200 149850 120000 6 io_out[33]
port 202 nsew signal output
rlabel metal2 s 154210 119200 154266 120000 6 io_out[34]
port 203 nsew signal output
rlabel metal2 s 158626 119200 158682 120000 6 io_out[35]
port 204 nsew signal output
rlabel metal2 s 163042 119200 163098 120000 6 io_out[36]
port 205 nsew signal output
rlabel metal2 s 167458 119200 167514 120000 6 io_out[37]
port 206 nsew signal output
rlabel metal2 s 16946 119200 17002 120000 6 io_out[3]
port 207 nsew signal output
rlabel metal2 s 21362 119200 21418 120000 6 io_out[4]
port 208 nsew signal output
rlabel metal2 s 25778 119200 25834 120000 6 io_out[5]
port 209 nsew signal output
rlabel metal2 s 30194 119200 30250 120000 6 io_out[6]
port 210 nsew signal output
rlabel metal2 s 34610 119200 34666 120000 6 io_out[7]
port 211 nsew signal output
rlabel metal2 s 39118 119200 39174 120000 6 io_out[8]
port 212 nsew signal output
rlabel metal2 s 43534 119200 43590 120000 6 io_out[9]
port 213 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 irq[0]
port 214 nsew signal output
rlabel metal2 s 177762 119200 177818 120000 6 irq[1]
port 215 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 irq[2]
port 216 nsew signal output
rlabel metal3 s 0 416 800 536 6 mem1_data_i[0]
port 217 nsew signal input
rlabel metal3 s 0 51416 800 51536 6 mem1_data_i[10]
port 218 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 mem1_data_i[11]
port 219 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 mem1_data_i[12]
port 220 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 mem1_data_i[13]
port 221 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 mem1_data_i[14]
port 222 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 mem1_data_i[15]
port 223 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 mem1_data_i[16]
port 224 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 mem1_data_i[17]
port 225 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 mem1_data_i[18]
port 226 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 mem1_data_i[19]
port 227 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 mem1_data_i[1]
port 228 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 mem1_data_i[20]
port 229 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 mem1_data_i[21]
port 230 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 mem1_data_i[22]
port 231 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 mem1_data_i[23]
port 232 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 mem1_data_i[24]
port 233 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 mem1_data_i[25]
port 234 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 mem1_data_i[26]
port 235 nsew signal input
rlabel metal3 s 0 101600 800 101720 6 mem1_data_i[27]
port 236 nsew signal input
rlabel metal3 s 0 104592 800 104712 6 mem1_data_i[28]
port 237 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 mem1_data_i[29]
port 238 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 mem1_data_i[2]
port 239 nsew signal input
rlabel metal3 s 0 110440 800 110560 6 mem1_data_i[30]
port 240 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 mem1_data_i[31]
port 241 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 mem1_data_i[3]
port 242 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 mem1_data_i[4]
port 243 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 mem1_data_i[5]
port 244 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 mem1_data_i[6]
port 245 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 mem1_data_i[7]
port 246 nsew signal input
rlabel metal3 s 0 43664 800 43784 6 mem1_data_i[8]
port 247 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 mem1_data_i[9]
port 248 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 mem_data_i[0]
port 249 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 mem_data_i[10]
port 250 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 mem_data_i[11]
port 251 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 mem_data_i[12]
port 252 nsew signal input
rlabel metal3 s 0 61344 800 61464 6 mem_data_i[13]
port 253 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 mem_data_i[14]
port 254 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 mem_data_i[15]
port 255 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 mem_data_i[16]
port 256 nsew signal input
rlabel metal3 s 0 73040 800 73160 6 mem_data_i[17]
port 257 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 mem_data_i[18]
port 258 nsew signal input
rlabel metal3 s 0 79024 800 79144 6 mem_data_i[19]
port 259 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 mem_data_i[1]
port 260 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 mem_data_i[20]
port 261 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 mem_data_i[21]
port 262 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 mem_data_i[22]
port 263 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 mem_data_i[23]
port 264 nsew signal input
rlabel metal3 s 0 93712 800 93832 6 mem_data_i[24]
port 265 nsew signal input
rlabel metal3 s 0 96704 800 96824 6 mem_data_i[25]
port 266 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 mem_data_i[26]
port 267 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 mem_data_i[27]
port 268 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 mem_data_i[28]
port 269 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 mem_data_i[29]
port 270 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 mem_data_i[2]
port 271 nsew signal input
rlabel metal3 s 0 111392 800 111512 6 mem_data_i[30]
port 272 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 mem_data_i[31]
port 273 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 mem_data_i[3]
port 274 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 mem_data_i[4]
port 275 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 mem_data_i[5]
port 276 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 mem_data_i[6]
port 277 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 mem_data_i[7]
port 278 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 mem_data_i[8]
port 279 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 mem_data_i[9]
port 280 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 mem_data_o[0]
port 281 nsew signal output
rlabel metal3 s 0 53456 800 53576 6 mem_data_o[10]
port 282 nsew signal output
rlabel metal3 s 0 56448 800 56568 6 mem_data_o[11]
port 283 nsew signal output
rlabel metal3 s 0 59304 800 59424 6 mem_data_o[12]
port 284 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 mem_data_o[13]
port 285 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 mem_data_o[14]
port 286 nsew signal output
rlabel metal3 s 0 68144 800 68264 6 mem_data_o[15]
port 287 nsew signal output
rlabel metal3 s 0 71136 800 71256 6 mem_data_o[16]
port 288 nsew signal output
rlabel metal3 s 0 74128 800 74248 6 mem_data_o[17]
port 289 nsew signal output
rlabel metal3 s 0 76984 800 77104 6 mem_data_o[18]
port 290 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 mem_data_o[19]
port 291 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 mem_data_o[1]
port 292 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 mem_data_o[20]
port 293 nsew signal output
rlabel metal3 s 0 85824 800 85944 6 mem_data_o[21]
port 294 nsew signal output
rlabel metal3 s 0 88816 800 88936 6 mem_data_o[22]
port 295 nsew signal output
rlabel metal3 s 0 91808 800 91928 6 mem_data_o[23]
port 296 nsew signal output
rlabel metal3 s 0 94800 800 94920 6 mem_data_o[24]
port 297 nsew signal output
rlabel metal3 s 0 97656 800 97776 6 mem_data_o[25]
port 298 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 mem_data_o[26]
port 299 nsew signal output
rlabel metal3 s 0 103640 800 103760 6 mem_data_o[27]
port 300 nsew signal output
rlabel metal3 s 0 106496 800 106616 6 mem_data_o[28]
port 301 nsew signal output
rlabel metal3 s 0 109488 800 109608 6 mem_data_o[29]
port 302 nsew signal output
rlabel metal3 s 0 16056 800 16176 6 mem_data_o[2]
port 303 nsew signal output
rlabel metal3 s 0 112480 800 112600 6 mem_data_o[30]
port 304 nsew signal output
rlabel metal3 s 0 115336 800 115456 6 mem_data_o[31]
port 305 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 mem_data_o[3]
port 306 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 mem_data_o[4]
port 307 nsew signal output
rlabel metal3 s 0 30880 800 31000 6 mem_data_o[5]
port 308 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 mem_data_o[6]
port 309 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 mem_data_o[7]
port 310 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 mem_data_o[8]
port 311 nsew signal output
rlabel metal3 s 0 50464 800 50584 6 mem_data_o[9]
port 312 nsew signal output
rlabel metal3 s 0 3272 800 3392 6 mem_raddr_o[0]
port 313 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 mem_raddr_o[1]
port 314 nsew signal output
rlabel metal3 s 0 17008 800 17128 6 mem_raddr_o[2]
port 315 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 mem_raddr_o[3]
port 316 nsew signal output
rlabel metal3 s 0 26936 800 27056 6 mem_raddr_o[4]
port 317 nsew signal output
rlabel metal3 s 0 31832 800 31952 6 mem_raddr_o[5]
port 318 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 mem_raddr_o[6]
port 319 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 mem_raddr_o[7]
port 320 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 mem_raddr_o[8]
port 321 nsew signal output
rlabel metal3 s 0 4224 800 4344 6 mem_renb_o[0]
port 322 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 mem_renb_o[1]
port 323 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 mem_waddr_o[0]
port 324 nsew signal output
rlabel metal3 s 0 12112 800 12232 6 mem_waddr_o[1]
port 325 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 mem_waddr_o[2]
port 326 nsew signal output
rlabel metal3 s 0 22992 800 23112 6 mem_waddr_o[3]
port 327 nsew signal output
rlabel metal3 s 0 27888 800 28008 6 mem_waddr_o[4]
port 328 nsew signal output
rlabel metal3 s 0 32784 800 32904 6 mem_waddr_o[5]
port 329 nsew signal output
rlabel metal3 s 0 37680 800 37800 6 mem_waddr_o[6]
port 330 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 mem_waddr_o[7]
port 331 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 mem_waddr_o[8]
port 332 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 mem_wenb_o[0]
port 333 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 mem_wenb_o[1]
port 334 nsew signal output
rlabel metal3 s 179200 552 180000 672 6 oversample_o[0]
port 335 nsew signal output
rlabel metal3 s 179200 1640 180000 1760 6 oversample_o[1]
port 336 nsew signal output
rlabel metal3 s 179200 2728 180000 2848 6 oversample_o[2]
port 337 nsew signal output
rlabel metal3 s 179200 3816 180000 3936 6 oversample_o[3]
port 338 nsew signal output
rlabel metal3 s 179200 4904 180000 5024 6 oversample_o[4]
port 339 nsew signal output
rlabel metal3 s 179200 5992 180000 6112 6 oversample_o[5]
port 340 nsew signal output
rlabel metal3 s 179200 7080 180000 7200 6 oversample_o[6]
port 341 nsew signal output
rlabel metal3 s 179200 8168 180000 8288 6 oversample_o[7]
port 342 nsew signal output
rlabel metal3 s 179200 9256 180000 9376 6 oversample_o[8]
port 343 nsew signal output
rlabel metal3 s 179200 10344 180000 10464 6 oversample_o[9]
port 344 nsew signal output
rlabel metal2 s 173346 119200 173402 120000 6 sinc3_en_o[0]
port 345 nsew signal output
rlabel metal2 s 174818 119200 174874 120000 6 sinc3_en_o[1]
port 346 nsew signal output
rlabel metal2 s 176290 119200 176346 120000 6 sinc3_en_o[2]
port 347 nsew signal output
rlabel metal2 s 168930 119200 168986 120000 6 vco_enb_o[0]
port 348 nsew signal output
rlabel metal2 s 170402 119200 170458 120000 6 vco_enb_o[1]
port 349 nsew signal output
rlabel metal2 s 171874 119200 171930 120000 6 vco_enb_o[2]
port 350 nsew signal output
rlabel metal2 s 846 0 902 800 6 wb_clk_i
port 351 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wb_rst_i
port 352 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_ack_o
port 353 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[0]
port 354 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 wbs_adr_i[10]
port 355 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 wbs_adr_i[11]
port 356 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_adr_i[12]
port 357 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_adr_i[13]
port 358 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[14]
port 359 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 wbs_adr_i[15]
port 360 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 wbs_adr_i[16]
port 361 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_adr_i[17]
port 362 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 wbs_adr_i[18]
port 363 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 wbs_adr_i[19]
port 364 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[1]
port 365 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 wbs_adr_i[20]
port 366 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 wbs_adr_i[21]
port 367 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 wbs_adr_i[22]
port 368 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 wbs_adr_i[23]
port 369 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 wbs_adr_i[24]
port 370 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 wbs_adr_i[25]
port 371 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 wbs_adr_i[26]
port 372 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 wbs_adr_i[27]
port 373 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 wbs_adr_i[28]
port 374 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 wbs_adr_i[29]
port 375 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[2]
port 376 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 wbs_adr_i[30]
port 377 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 wbs_adr_i[31]
port 378 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[3]
port 379 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[4]
port 380 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_adr_i[5]
port 381 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[6]
port 382 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_adr_i[7]
port 383 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_adr_i[8]
port 384 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 wbs_adr_i[9]
port 385 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_cyc_i
port 386 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[0]
port 387 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wbs_dat_i[10]
port 388 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_i[11]
port 389 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_i[12]
port 390 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_i[13]
port 391 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_i[14]
port 392 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 wbs_dat_i[15]
port 393 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 wbs_dat_i[16]
port 394 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 wbs_dat_i[17]
port 395 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 wbs_dat_i[18]
port 396 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 wbs_dat_i[19]
port 397 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[1]
port 398 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 wbs_dat_i[20]
port 399 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_i[21]
port 400 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 wbs_dat_i[22]
port 401 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 wbs_dat_i[23]
port 402 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 wbs_dat_i[24]
port 403 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 wbs_dat_i[25]
port 404 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 wbs_dat_i[26]
port 405 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 wbs_dat_i[27]
port 406 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 wbs_dat_i[28]
port 407 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 wbs_dat_i[29]
port 408 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[2]
port 409 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 wbs_dat_i[30]
port 410 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 wbs_dat_i[31]
port 411 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[3]
port 412 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_i[4]
port 413 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_i[5]
port 414 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_i[6]
port 415 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[7]
port 416 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 wbs_dat_i[8]
port 417 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[9]
port 418 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[0]
port 419 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[10]
port 420 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 wbs_dat_o[11]
port 421 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_o[12]
port 422 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_o[13]
port 423 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_o[14]
port 424 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 wbs_dat_o[15]
port 425 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 wbs_dat_o[16]
port 426 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 wbs_dat_o[17]
port 427 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 wbs_dat_o[18]
port 428 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 wbs_dat_o[19]
port 429 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[1]
port 430 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 wbs_dat_o[20]
port 431 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 wbs_dat_o[21]
port 432 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 wbs_dat_o[22]
port 433 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 wbs_dat_o[23]
port 434 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 wbs_dat_o[24]
port 435 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 wbs_dat_o[25]
port 436 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 wbs_dat_o[26]
port 437 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 wbs_dat_o[27]
port 438 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 wbs_dat_o[28]
port 439 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 wbs_dat_o[29]
port 440 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[2]
port 441 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 wbs_dat_o[30]
port 442 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 wbs_dat_o[31]
port 443 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_o[3]
port 444 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[4]
port 445 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[5]
port 446 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[6]
port 447 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[7]
port 448 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_o[8]
port 449 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 wbs_dat_o[9]
port 450 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_sel_i[0]
port 451 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_sel_i[1]
port 452 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_sel_i[2]
port 453 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_sel_i[3]
port 454 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_stb_i
port 455 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_we_i
port 456 nsew signal input
rlabel metal3 s 0 117376 800 117496 6 wmask_o[0]
port 457 nsew signal output
rlabel metal2 s 179234 119200 179290 120000 6 wmask_o[1]
port 458 nsew signal output
rlabel metal3 s 0 119280 800 119400 6 wmask_o[2]
port 459 nsew signal output
rlabel metal3 s 179200 119280 180000 119400 6 wmask_o[3]
port 460 nsew signal output
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 461 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 462 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 463 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 464 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 465 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 466 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 467 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 468 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 469 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 470 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 471 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 472 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 473 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 474 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 475 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 476 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 477 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 478 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 479 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 480 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 481 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 482 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 483 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 484 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 485 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 486 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 487 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 488 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 489 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 490 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 491 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 492 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 493 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 494 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 495 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 496 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 497 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 498 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 499 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 500 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 501 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 502 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 503 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 504 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 505 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 506 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 507 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 508 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 8644214
string GDS_START 671862
<< end >>

