VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_adc
  CLASS BLOCK ;
  FOREIGN vco_adc ;
  ORIGIN 0.000 0.000 ;
  SIZE 270.000 BY 270.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END clk
  PIN data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END data_out[0]
  PIN data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END data_out[10]
  PIN data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END data_out[11]
  PIN data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 0.000 110.310 4.000 ;
    END
  END data_out[12]
  PIN data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 118.310 0.000 118.590 4.000 ;
    END
  END data_out[13]
  PIN data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.130 0.000 126.410 4.000 ;
    END
  END data_out[14]
  PIN data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 0.000 134.690 4.000 ;
    END
  END data_out[15]
  PIN data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END data_out[16]
  PIN data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END data_out[17]
  PIN data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 4.000 ;
    END
  END data_out[18]
  PIN data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 4.000 ;
    END
  END data_out[19]
  PIN data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.870 0.000 20.150 4.000 ;
    END
  END data_out[1]
  PIN data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 4.000 ;
    END
  END data_out[20]
  PIN data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END data_out[21]
  PIN data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 4.000 ;
    END
  END data_out[22]
  PIN data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 0.000 200.010 4.000 ;
    END
  END data_out[23]
  PIN data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END data_out[24]
  PIN data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END data_out[25]
  PIN data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END data_out[26]
  PIN data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 0.000 233.130 4.000 ;
    END
  END data_out[27]
  PIN data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 240.670 0.000 240.950 4.000 ;
    END
  END data_out[28]
  PIN data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 0.000 249.230 4.000 ;
    END
  END data_out[29]
  PIN data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 0.000 28.430 4.000 ;
    END
  END data_out[2]
  PIN data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 0.000 257.510 4.000 ;
    END
  END data_out[30]
  PIN data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END data_out[31]
  PIN data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 0.000 36.710 4.000 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 4.000 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 4.000 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END data_out[7]
  PIN data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END data_out[8]
  PIN data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END data_out[9]
  PIN data_valid_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 0.000 4.050 4.000 ;
    END
  END data_valid_out
  PIN enable_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.720 4.000 52.320 ;
    END
  END enable_in
  PIN oversample_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.120 4.000 72.720 ;
    END
  END oversample_in[0]
  PIN oversample_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.200 4.000 93.800 ;
    END
  END oversample_in[1]
  PIN oversample_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END oversample_in[2]
  PIN oversample_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.680 4.000 135.280 ;
    END
  END oversample_in[3]
  PIN oversample_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 155.080 4.000 155.680 ;
    END
  END oversample_in[4]
  PIN oversample_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.160 4.000 176.760 ;
    END
  END oversample_in[5]
  PIN oversample_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END oversample_in[6]
  PIN oversample_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END oversample_in[7]
  PIN oversample_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END oversample_in[8]
  PIN oversample_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.120 4.000 259.720 ;
    END
  END oversample_in[9]
  PIN phase_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 266.000 12.330 270.000 ;
    END
  END phase_in[0]
  PIN phase_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 266.000 257.510 270.000 ;
    END
  END phase_in[10]
  PIN phase_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 36.430 266.000 36.710 270.000 ;
    END
  END phase_in[1]
  PIN phase_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.810 266.000 61.090 270.000 ;
    END
  END phase_in[2]
  PIN phase_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 266.000 85.930 270.000 ;
    END
  END phase_in[3]
  PIN phase_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 266.000 110.310 270.000 ;
    END
  END phase_in[4]
  PIN phase_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 266.000 134.690 270.000 ;
    END
  END phase_in[5]
  PIN phase_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 266.000 159.530 270.000 ;
    END
  END phase_in[6]
  PIN phase_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 266.000 183.910 270.000 ;
    END
  END phase_in[7]
  PIN phase_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 266.000 208.290 270.000 ;
    END
  END phase_in[8]
  PIN phase_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 266.000 233.130 270.000 ;
    END
  END phase_in[9]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END rst
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 258.640 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 258.640 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 258.640 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 258.640 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 3.145 264.040 258.485 ;
      LAYER met1 ;
        RECT 0.070 2.140 265.810 259.380 ;
      LAYER met2 ;
        RECT 0.090 265.720 11.770 266.000 ;
        RECT 12.610 265.720 36.150 266.000 ;
        RECT 36.990 265.720 60.530 266.000 ;
        RECT 61.370 265.720 85.370 266.000 ;
        RECT 86.210 265.720 109.750 266.000 ;
        RECT 110.590 265.720 134.130 266.000 ;
        RECT 134.970 265.720 158.970 266.000 ;
        RECT 159.810 265.720 183.350 266.000 ;
        RECT 184.190 265.720 207.730 266.000 ;
        RECT 208.570 265.720 232.570 266.000 ;
        RECT 233.410 265.720 256.950 266.000 ;
        RECT 257.790 265.720 265.780 266.000 ;
        RECT 0.090 4.280 265.780 265.720 ;
        RECT 0.090 2.390 3.490 4.280 ;
        RECT 4.330 2.390 11.310 4.280 ;
        RECT 12.150 2.390 19.590 4.280 ;
        RECT 20.430 2.390 27.870 4.280 ;
        RECT 28.710 2.390 36.150 4.280 ;
        RECT 36.990 2.390 43.970 4.280 ;
        RECT 44.810 2.390 52.250 4.280 ;
        RECT 53.090 2.390 60.530 4.280 ;
        RECT 61.370 2.390 68.810 4.280 ;
        RECT 69.650 2.390 77.090 4.280 ;
        RECT 77.930 2.390 84.910 4.280 ;
        RECT 85.750 2.390 93.190 4.280 ;
        RECT 94.030 2.390 101.470 4.280 ;
        RECT 102.310 2.390 109.750 4.280 ;
        RECT 110.590 2.390 118.030 4.280 ;
        RECT 118.870 2.390 125.850 4.280 ;
        RECT 126.690 2.390 134.130 4.280 ;
        RECT 134.970 2.390 142.410 4.280 ;
        RECT 143.250 2.390 150.690 4.280 ;
        RECT 151.530 2.390 158.510 4.280 ;
        RECT 159.350 2.390 166.790 4.280 ;
        RECT 167.630 2.390 175.070 4.280 ;
        RECT 175.910 2.390 183.350 4.280 ;
        RECT 184.190 2.390 191.630 4.280 ;
        RECT 192.470 2.390 199.450 4.280 ;
        RECT 200.290 2.390 207.730 4.280 ;
        RECT 208.570 2.390 216.010 4.280 ;
        RECT 216.850 2.390 224.290 4.280 ;
        RECT 225.130 2.390 232.570 4.280 ;
        RECT 233.410 2.390 240.390 4.280 ;
        RECT 241.230 2.390 248.670 4.280 ;
        RECT 249.510 2.390 256.950 4.280 ;
        RECT 257.790 2.390 265.230 4.280 ;
      LAYER met3 ;
        RECT 4.400 258.720 260.295 259.585 ;
        RECT 0.065 239.040 260.295 258.720 ;
        RECT 4.400 237.640 260.295 239.040 ;
        RECT 0.065 218.640 260.295 237.640 ;
        RECT 4.400 217.240 260.295 218.640 ;
        RECT 0.065 197.560 260.295 217.240 ;
        RECT 4.400 196.160 260.295 197.560 ;
        RECT 0.065 177.160 260.295 196.160 ;
        RECT 4.400 175.760 260.295 177.160 ;
        RECT 0.065 156.080 260.295 175.760 ;
        RECT 4.400 154.680 260.295 156.080 ;
        RECT 0.065 135.680 260.295 154.680 ;
        RECT 4.400 134.280 260.295 135.680 ;
        RECT 0.065 114.600 260.295 134.280 ;
        RECT 4.400 113.200 260.295 114.600 ;
        RECT 0.065 94.200 260.295 113.200 ;
        RECT 4.400 92.800 260.295 94.200 ;
        RECT 0.065 73.120 260.295 92.800 ;
        RECT 4.400 71.720 260.295 73.120 ;
        RECT 0.065 52.720 260.295 71.720 ;
        RECT 4.400 51.320 260.295 52.720 ;
        RECT 0.065 31.640 260.295 51.320 ;
        RECT 4.400 30.240 260.295 31.640 ;
        RECT 0.065 11.240 260.295 30.240 ;
        RECT 4.400 9.840 260.295 11.240 ;
        RECT 0.065 6.975 260.295 9.840 ;
      LAYER met4 ;
        RECT 0.295 11.055 20.640 231.705 ;
        RECT 23.040 11.055 97.440 231.705 ;
        RECT 99.840 11.055 174.240 231.705 ;
        RECT 176.640 11.055 251.040 231.705 ;
        RECT 253.440 11.055 258.650 231.705 ;
      LAYER met5 ;
        RECT 18.980 11.100 258.860 12.700 ;
  END
END vco_adc
END LIBRARY

