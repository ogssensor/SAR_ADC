magic
tech sky130A
magscale 1 2
timestamp 1623830371
<< obsli1 >>
rect 1104 1377 178848 117521
<< obsm1 >>
rect 474 1368 179570 118244
<< metal2 >>
rect 478 119200 534 120000
rect 1398 119200 1454 120000
rect 2410 119200 2466 120000
rect 3330 119200 3386 120000
rect 4342 119200 4398 120000
rect 5262 119200 5318 120000
rect 6274 119200 6330 120000
rect 7286 119200 7342 120000
rect 8206 119200 8262 120000
rect 9218 119200 9274 120000
rect 10138 119200 10194 120000
rect 11150 119200 11206 120000
rect 12070 119200 12126 120000
rect 13082 119200 13138 120000
rect 14094 119200 14150 120000
rect 15014 119200 15070 120000
rect 16026 119200 16082 120000
rect 16946 119200 17002 120000
rect 17958 119200 18014 120000
rect 18878 119200 18934 120000
rect 19890 119200 19946 120000
rect 20902 119200 20958 120000
rect 21822 119200 21878 120000
rect 22834 119200 22890 120000
rect 23754 119200 23810 120000
rect 24766 119200 24822 120000
rect 25778 119200 25834 120000
rect 26698 119200 26754 120000
rect 27710 119200 27766 120000
rect 28630 119200 28686 120000
rect 29642 119200 29698 120000
rect 30562 119200 30618 120000
rect 31574 119200 31630 120000
rect 32586 119200 32642 120000
rect 33506 119200 33562 120000
rect 34518 119200 34574 120000
rect 35438 119200 35494 120000
rect 36450 119200 36506 120000
rect 37370 119200 37426 120000
rect 38382 119200 38438 120000
rect 39394 119200 39450 120000
rect 40314 119200 40370 120000
rect 41326 119200 41382 120000
rect 42246 119200 42302 120000
rect 43258 119200 43314 120000
rect 44270 119200 44326 120000
rect 45190 119200 45246 120000
rect 46202 119200 46258 120000
rect 47122 119200 47178 120000
rect 48134 119200 48190 120000
rect 49054 119200 49110 120000
rect 50066 119200 50122 120000
rect 51078 119200 51134 120000
rect 51998 119200 52054 120000
rect 53010 119200 53066 120000
rect 53930 119200 53986 120000
rect 54942 119200 54998 120000
rect 55862 119200 55918 120000
rect 56874 119200 56930 120000
rect 57886 119200 57942 120000
rect 58806 119200 58862 120000
rect 59818 119200 59874 120000
rect 60738 119200 60794 120000
rect 61750 119200 61806 120000
rect 62762 119200 62818 120000
rect 63682 119200 63738 120000
rect 64694 119200 64750 120000
rect 65614 119200 65670 120000
rect 66626 119200 66682 120000
rect 67546 119200 67602 120000
rect 68558 119200 68614 120000
rect 69570 119200 69626 120000
rect 70490 119200 70546 120000
rect 71502 119200 71558 120000
rect 72422 119200 72478 120000
rect 73434 119200 73490 120000
rect 74354 119200 74410 120000
rect 75366 119200 75422 120000
rect 76378 119200 76434 120000
rect 77298 119200 77354 120000
rect 78310 119200 78366 120000
rect 79230 119200 79286 120000
rect 80242 119200 80298 120000
rect 81254 119200 81310 120000
rect 82174 119200 82230 120000
rect 83186 119200 83242 120000
rect 84106 119200 84162 120000
rect 85118 119200 85174 120000
rect 86038 119200 86094 120000
rect 87050 119200 87106 120000
rect 88062 119200 88118 120000
rect 88982 119200 89038 120000
rect 89994 119200 90050 120000
rect 90914 119200 90970 120000
rect 91926 119200 91982 120000
rect 92846 119200 92902 120000
rect 93858 119200 93914 120000
rect 94870 119200 94926 120000
rect 95790 119200 95846 120000
rect 96802 119200 96858 120000
rect 97722 119200 97778 120000
rect 98734 119200 98790 120000
rect 99654 119200 99710 120000
rect 100666 119200 100722 120000
rect 101678 119200 101734 120000
rect 102598 119200 102654 120000
rect 103610 119200 103666 120000
rect 104530 119200 104586 120000
rect 105542 119200 105598 120000
rect 106554 119200 106610 120000
rect 107474 119200 107530 120000
rect 108486 119200 108542 120000
rect 109406 119200 109462 120000
rect 110418 119200 110474 120000
rect 111338 119200 111394 120000
rect 112350 119200 112406 120000
rect 113362 119200 113418 120000
rect 114282 119200 114338 120000
rect 115294 119200 115350 120000
rect 116214 119200 116270 120000
rect 117226 119200 117282 120000
rect 118146 119200 118202 120000
rect 119158 119200 119214 120000
rect 120170 119200 120226 120000
rect 121090 119200 121146 120000
rect 122102 119200 122158 120000
rect 123022 119200 123078 120000
rect 124034 119200 124090 120000
rect 125046 119200 125102 120000
rect 125966 119200 126022 120000
rect 126978 119200 127034 120000
rect 127898 119200 127954 120000
rect 128910 119200 128966 120000
rect 129830 119200 129886 120000
rect 130842 119200 130898 120000
rect 131854 119200 131910 120000
rect 132774 119200 132830 120000
rect 133786 119200 133842 120000
rect 134706 119200 134762 120000
rect 135718 119200 135774 120000
rect 136638 119200 136694 120000
rect 137650 119200 137706 120000
rect 138662 119200 138718 120000
rect 139582 119200 139638 120000
rect 140594 119200 140650 120000
rect 141514 119200 141570 120000
rect 142526 119200 142582 120000
rect 143538 119200 143594 120000
rect 144458 119200 144514 120000
rect 145470 119200 145526 120000
rect 146390 119200 146446 120000
rect 147402 119200 147458 120000
rect 148322 119200 148378 120000
rect 149334 119200 149390 120000
rect 150346 119200 150402 120000
rect 151266 119200 151322 120000
rect 152278 119200 152334 120000
rect 153198 119200 153254 120000
rect 154210 119200 154266 120000
rect 155130 119200 155186 120000
rect 156142 119200 156198 120000
rect 157154 119200 157210 120000
rect 158074 119200 158130 120000
rect 159086 119200 159142 120000
rect 160006 119200 160062 120000
rect 161018 119200 161074 120000
rect 162030 119200 162086 120000
rect 162950 119200 163006 120000
rect 163962 119200 164018 120000
rect 164882 119200 164938 120000
rect 165894 119200 165950 120000
rect 166814 119200 166870 120000
rect 167826 119200 167882 120000
rect 168838 119200 168894 120000
rect 169758 119200 169814 120000
rect 170770 119200 170826 120000
rect 171690 119200 171746 120000
rect 172702 119200 172758 120000
rect 173622 119200 173678 120000
rect 174634 119200 174690 120000
rect 175646 119200 175702 120000
rect 176566 119200 176622 120000
rect 177578 119200 177634 120000
rect 178498 119200 178554 120000
rect 179510 119200 179566 120000
rect 570 0 626 800
rect 1766 0 1822 800
rect 3054 0 3110 800
rect 4250 0 4306 800
rect 5538 0 5594 800
rect 6734 0 6790 800
rect 8022 0 8078 800
rect 9310 0 9366 800
rect 10506 0 10562 800
rect 11794 0 11850 800
rect 12990 0 13046 800
rect 14278 0 14334 800
rect 15566 0 15622 800
rect 16762 0 16818 800
rect 18050 0 18106 800
rect 19246 0 19302 800
rect 20534 0 20590 800
rect 21822 0 21878 800
rect 23018 0 23074 800
rect 24306 0 24362 800
rect 25502 0 25558 800
rect 26790 0 26846 800
rect 27986 0 28042 800
rect 29274 0 29330 800
rect 30562 0 30618 800
rect 31758 0 31814 800
rect 33046 0 33102 800
rect 34242 0 34298 800
rect 35530 0 35586 800
rect 36818 0 36874 800
rect 38014 0 38070 800
rect 39302 0 39358 800
rect 40498 0 40554 800
rect 41786 0 41842 800
rect 43074 0 43130 800
rect 44270 0 44326 800
rect 45558 0 45614 800
rect 46754 0 46810 800
rect 48042 0 48098 800
rect 49330 0 49386 800
rect 50526 0 50582 800
rect 51814 0 51870 800
rect 53010 0 53066 800
rect 54298 0 54354 800
rect 55494 0 55550 800
rect 56782 0 56838 800
rect 58070 0 58126 800
rect 59266 0 59322 800
rect 60554 0 60610 800
rect 61750 0 61806 800
rect 63038 0 63094 800
rect 64326 0 64382 800
rect 65522 0 65578 800
rect 66810 0 66866 800
rect 68006 0 68062 800
rect 69294 0 69350 800
rect 70582 0 70638 800
rect 71778 0 71834 800
rect 73066 0 73122 800
rect 74262 0 74318 800
rect 75550 0 75606 800
rect 76838 0 76894 800
rect 78034 0 78090 800
rect 79322 0 79378 800
rect 80518 0 80574 800
rect 81806 0 81862 800
rect 83002 0 83058 800
rect 84290 0 84346 800
rect 85578 0 85634 800
rect 86774 0 86830 800
rect 88062 0 88118 800
rect 89258 0 89314 800
rect 90546 0 90602 800
rect 91834 0 91890 800
rect 93030 0 93086 800
rect 94318 0 94374 800
rect 95514 0 95570 800
rect 96802 0 96858 800
rect 98090 0 98146 800
rect 99286 0 99342 800
rect 100574 0 100630 800
rect 101770 0 101826 800
rect 103058 0 103114 800
rect 104254 0 104310 800
rect 105542 0 105598 800
rect 106830 0 106886 800
rect 108026 0 108082 800
rect 109314 0 109370 800
rect 110510 0 110566 800
rect 111798 0 111854 800
rect 113086 0 113142 800
rect 114282 0 114338 800
rect 115570 0 115626 800
rect 116766 0 116822 800
rect 118054 0 118110 800
rect 119342 0 119398 800
rect 120538 0 120594 800
rect 121826 0 121882 800
rect 123022 0 123078 800
rect 124310 0 124366 800
rect 125598 0 125654 800
rect 126794 0 126850 800
rect 128082 0 128138 800
rect 129278 0 129334 800
rect 130566 0 130622 800
rect 131762 0 131818 800
rect 133050 0 133106 800
rect 134338 0 134394 800
rect 135534 0 135590 800
rect 136822 0 136878 800
rect 138018 0 138074 800
rect 139306 0 139362 800
rect 140594 0 140650 800
rect 141790 0 141846 800
rect 143078 0 143134 800
rect 144274 0 144330 800
rect 145562 0 145618 800
rect 146850 0 146906 800
rect 148046 0 148102 800
rect 149334 0 149390 800
rect 150530 0 150586 800
rect 151818 0 151874 800
rect 153106 0 153162 800
rect 154302 0 154358 800
rect 155590 0 155646 800
rect 156786 0 156842 800
rect 158074 0 158130 800
rect 159270 0 159326 800
rect 160558 0 160614 800
rect 161846 0 161902 800
rect 163042 0 163098 800
rect 164330 0 164386 800
rect 165526 0 165582 800
rect 166814 0 166870 800
rect 168102 0 168158 800
rect 169298 0 169354 800
rect 170586 0 170642 800
rect 171782 0 171838 800
rect 173070 0 173126 800
rect 174358 0 174414 800
rect 175554 0 175610 800
rect 176842 0 176898 800
rect 178038 0 178094 800
rect 179326 0 179382 800
<< obsm2 >>
rect 590 119144 1342 119785
rect 1510 119144 2354 119785
rect 2522 119144 3274 119785
rect 3442 119144 4286 119785
rect 4454 119144 5206 119785
rect 5374 119144 6218 119785
rect 6386 119144 7230 119785
rect 7398 119144 8150 119785
rect 8318 119144 9162 119785
rect 9330 119144 10082 119785
rect 10250 119144 11094 119785
rect 11262 119144 12014 119785
rect 12182 119144 13026 119785
rect 13194 119144 14038 119785
rect 14206 119144 14958 119785
rect 15126 119144 15970 119785
rect 16138 119144 16890 119785
rect 17058 119144 17902 119785
rect 18070 119144 18822 119785
rect 18990 119144 19834 119785
rect 20002 119144 20846 119785
rect 21014 119144 21766 119785
rect 21934 119144 22778 119785
rect 22946 119144 23698 119785
rect 23866 119144 24710 119785
rect 24878 119144 25722 119785
rect 25890 119144 26642 119785
rect 26810 119144 27654 119785
rect 27822 119144 28574 119785
rect 28742 119144 29586 119785
rect 29754 119144 30506 119785
rect 30674 119144 31518 119785
rect 31686 119144 32530 119785
rect 32698 119144 33450 119785
rect 33618 119144 34462 119785
rect 34630 119144 35382 119785
rect 35550 119144 36394 119785
rect 36562 119144 37314 119785
rect 37482 119144 38326 119785
rect 38494 119144 39338 119785
rect 39506 119144 40258 119785
rect 40426 119144 41270 119785
rect 41438 119144 42190 119785
rect 42358 119144 43202 119785
rect 43370 119144 44214 119785
rect 44382 119144 45134 119785
rect 45302 119144 46146 119785
rect 46314 119144 47066 119785
rect 47234 119144 48078 119785
rect 48246 119144 48998 119785
rect 49166 119144 50010 119785
rect 50178 119144 51022 119785
rect 51190 119144 51942 119785
rect 52110 119144 52954 119785
rect 53122 119144 53874 119785
rect 54042 119144 54886 119785
rect 55054 119144 55806 119785
rect 55974 119144 56818 119785
rect 56986 119144 57830 119785
rect 57998 119144 58750 119785
rect 58918 119144 59762 119785
rect 59930 119144 60682 119785
rect 60850 119144 61694 119785
rect 61862 119144 62706 119785
rect 62874 119144 63626 119785
rect 63794 119144 64638 119785
rect 64806 119144 65558 119785
rect 65726 119144 66570 119785
rect 66738 119144 67490 119785
rect 67658 119144 68502 119785
rect 68670 119144 69514 119785
rect 69682 119144 70434 119785
rect 70602 119144 71446 119785
rect 71614 119144 72366 119785
rect 72534 119144 73378 119785
rect 73546 119144 74298 119785
rect 74466 119144 75310 119785
rect 75478 119144 76322 119785
rect 76490 119144 77242 119785
rect 77410 119144 78254 119785
rect 78422 119144 79174 119785
rect 79342 119144 80186 119785
rect 80354 119144 81198 119785
rect 81366 119144 82118 119785
rect 82286 119144 83130 119785
rect 83298 119144 84050 119785
rect 84218 119144 85062 119785
rect 85230 119144 85982 119785
rect 86150 119144 86994 119785
rect 87162 119144 88006 119785
rect 88174 119144 88926 119785
rect 89094 119144 89938 119785
rect 90106 119144 90858 119785
rect 91026 119144 91870 119785
rect 92038 119144 92790 119785
rect 92958 119144 93802 119785
rect 93970 119144 94814 119785
rect 94982 119144 95734 119785
rect 95902 119144 96746 119785
rect 96914 119144 97666 119785
rect 97834 119144 98678 119785
rect 98846 119144 99598 119785
rect 99766 119144 100610 119785
rect 100778 119144 101622 119785
rect 101790 119144 102542 119785
rect 102710 119144 103554 119785
rect 103722 119144 104474 119785
rect 104642 119144 105486 119785
rect 105654 119144 106498 119785
rect 106666 119144 107418 119785
rect 107586 119144 108430 119785
rect 108598 119144 109350 119785
rect 109518 119144 110362 119785
rect 110530 119144 111282 119785
rect 111450 119144 112294 119785
rect 112462 119144 113306 119785
rect 113474 119144 114226 119785
rect 114394 119144 115238 119785
rect 115406 119144 116158 119785
rect 116326 119144 117170 119785
rect 117338 119144 118090 119785
rect 118258 119144 119102 119785
rect 119270 119144 120114 119785
rect 120282 119144 121034 119785
rect 121202 119144 122046 119785
rect 122214 119144 122966 119785
rect 123134 119144 123978 119785
rect 124146 119144 124990 119785
rect 125158 119144 125910 119785
rect 126078 119144 126922 119785
rect 127090 119144 127842 119785
rect 128010 119144 128854 119785
rect 129022 119144 129774 119785
rect 129942 119144 130786 119785
rect 130954 119144 131798 119785
rect 131966 119144 132718 119785
rect 132886 119144 133730 119785
rect 133898 119144 134650 119785
rect 134818 119144 135662 119785
rect 135830 119144 136582 119785
rect 136750 119144 137594 119785
rect 137762 119144 138606 119785
rect 138774 119144 139526 119785
rect 139694 119144 140538 119785
rect 140706 119144 141458 119785
rect 141626 119144 142470 119785
rect 142638 119144 143482 119785
rect 143650 119144 144402 119785
rect 144570 119144 145414 119785
rect 145582 119144 146334 119785
rect 146502 119144 147346 119785
rect 147514 119144 148266 119785
rect 148434 119144 149278 119785
rect 149446 119144 150290 119785
rect 150458 119144 151210 119785
rect 151378 119144 152222 119785
rect 152390 119144 153142 119785
rect 153310 119144 154154 119785
rect 154322 119144 155074 119785
rect 155242 119144 156086 119785
rect 156254 119144 157098 119785
rect 157266 119144 158018 119785
rect 158186 119144 159030 119785
rect 159198 119144 159950 119785
rect 160118 119144 160962 119785
rect 161130 119144 161974 119785
rect 162142 119144 162894 119785
rect 163062 119144 163906 119785
rect 164074 119144 164826 119785
rect 164994 119144 165838 119785
rect 166006 119144 166758 119785
rect 166926 119144 167770 119785
rect 167938 119144 168782 119785
rect 168950 119144 169702 119785
rect 169870 119144 170714 119785
rect 170882 119144 171634 119785
rect 171802 119144 172646 119785
rect 172814 119144 173566 119785
rect 173734 119144 174578 119785
rect 174746 119144 175590 119785
rect 175758 119144 176510 119785
rect 176678 119144 177522 119785
rect 177690 119144 178442 119785
rect 178610 119144 179454 119785
rect 480 856 179564 119144
rect 480 167 514 856
rect 682 167 1710 856
rect 1878 167 2998 856
rect 3166 167 4194 856
rect 4362 167 5482 856
rect 5650 167 6678 856
rect 6846 167 7966 856
rect 8134 167 9254 856
rect 9422 167 10450 856
rect 10618 167 11738 856
rect 11906 167 12934 856
rect 13102 167 14222 856
rect 14390 167 15510 856
rect 15678 167 16706 856
rect 16874 167 17994 856
rect 18162 167 19190 856
rect 19358 167 20478 856
rect 20646 167 21766 856
rect 21934 167 22962 856
rect 23130 167 24250 856
rect 24418 167 25446 856
rect 25614 167 26734 856
rect 26902 167 27930 856
rect 28098 167 29218 856
rect 29386 167 30506 856
rect 30674 167 31702 856
rect 31870 167 32990 856
rect 33158 167 34186 856
rect 34354 167 35474 856
rect 35642 167 36762 856
rect 36930 167 37958 856
rect 38126 167 39246 856
rect 39414 167 40442 856
rect 40610 167 41730 856
rect 41898 167 43018 856
rect 43186 167 44214 856
rect 44382 167 45502 856
rect 45670 167 46698 856
rect 46866 167 47986 856
rect 48154 167 49274 856
rect 49442 167 50470 856
rect 50638 167 51758 856
rect 51926 167 52954 856
rect 53122 167 54242 856
rect 54410 167 55438 856
rect 55606 167 56726 856
rect 56894 167 58014 856
rect 58182 167 59210 856
rect 59378 167 60498 856
rect 60666 167 61694 856
rect 61862 167 62982 856
rect 63150 167 64270 856
rect 64438 167 65466 856
rect 65634 167 66754 856
rect 66922 167 67950 856
rect 68118 167 69238 856
rect 69406 167 70526 856
rect 70694 167 71722 856
rect 71890 167 73010 856
rect 73178 167 74206 856
rect 74374 167 75494 856
rect 75662 167 76782 856
rect 76950 167 77978 856
rect 78146 167 79266 856
rect 79434 167 80462 856
rect 80630 167 81750 856
rect 81918 167 82946 856
rect 83114 167 84234 856
rect 84402 167 85522 856
rect 85690 167 86718 856
rect 86886 167 88006 856
rect 88174 167 89202 856
rect 89370 167 90490 856
rect 90658 167 91778 856
rect 91946 167 92974 856
rect 93142 167 94262 856
rect 94430 167 95458 856
rect 95626 167 96746 856
rect 96914 167 98034 856
rect 98202 167 99230 856
rect 99398 167 100518 856
rect 100686 167 101714 856
rect 101882 167 103002 856
rect 103170 167 104198 856
rect 104366 167 105486 856
rect 105654 167 106774 856
rect 106942 167 107970 856
rect 108138 167 109258 856
rect 109426 167 110454 856
rect 110622 167 111742 856
rect 111910 167 113030 856
rect 113198 167 114226 856
rect 114394 167 115514 856
rect 115682 167 116710 856
rect 116878 167 117998 856
rect 118166 167 119286 856
rect 119454 167 120482 856
rect 120650 167 121770 856
rect 121938 167 122966 856
rect 123134 167 124254 856
rect 124422 167 125542 856
rect 125710 167 126738 856
rect 126906 167 128026 856
rect 128194 167 129222 856
rect 129390 167 130510 856
rect 130678 167 131706 856
rect 131874 167 132994 856
rect 133162 167 134282 856
rect 134450 167 135478 856
rect 135646 167 136766 856
rect 136934 167 137962 856
rect 138130 167 139250 856
rect 139418 167 140538 856
rect 140706 167 141734 856
rect 141902 167 143022 856
rect 143190 167 144218 856
rect 144386 167 145506 856
rect 145674 167 146794 856
rect 146962 167 147990 856
rect 148158 167 149278 856
rect 149446 167 150474 856
rect 150642 167 151762 856
rect 151930 167 153050 856
rect 153218 167 154246 856
rect 154414 167 155534 856
rect 155702 167 156730 856
rect 156898 167 158018 856
rect 158186 167 159214 856
rect 159382 167 160502 856
rect 160670 167 161790 856
rect 161958 167 162986 856
rect 163154 167 164274 856
rect 164442 167 165470 856
rect 165638 167 166758 856
rect 166926 167 168046 856
rect 168214 167 169242 856
rect 169410 167 170530 856
rect 170698 167 171726 856
rect 171894 167 173014 856
rect 173182 167 174302 856
rect 174470 167 175498 856
rect 175666 167 176786 856
rect 176954 167 177982 856
rect 178150 167 179270 856
rect 179438 167 179564 856
<< metal3 >>
rect 0 119688 800 119808
rect 0 119416 800 119536
rect 0 119144 800 119264
rect 0 118872 800 118992
rect 0 118600 800 118720
rect 0 118328 800 118448
rect 179200 118464 180000 118584
rect 0 118056 800 118176
rect 0 117784 800 117904
rect 0 117512 800 117632
rect 0 117240 800 117360
rect 0 116968 800 117088
rect 0 116696 800 116816
rect 0 116424 800 116544
rect 0 116152 800 116272
rect 0 115744 800 115864
rect 179200 115744 180000 115864
rect 0 115472 800 115592
rect 0 115200 800 115320
rect 0 114928 800 115048
rect 0 114656 800 114776
rect 0 114384 800 114504
rect 0 114112 800 114232
rect 0 113840 800 113960
rect 0 113568 800 113688
rect 0 113296 800 113416
rect 0 113024 800 113144
rect 179200 113024 180000 113144
rect 0 112752 800 112872
rect 0 112480 800 112600
rect 0 112208 800 112328
rect 0 111800 800 111920
rect 0 111528 800 111648
rect 0 111256 800 111376
rect 0 110984 800 111104
rect 0 110712 800 110832
rect 0 110440 800 110560
rect 0 110168 800 110288
rect 179200 110304 180000 110424
rect 0 109896 800 110016
rect 0 109624 800 109744
rect 0 109352 800 109472
rect 0 109080 800 109200
rect 0 108808 800 108928
rect 0 108536 800 108656
rect 0 108264 800 108384
rect 0 107856 800 107976
rect 0 107584 800 107704
rect 179200 107584 180000 107704
rect 0 107312 800 107432
rect 0 107040 800 107160
rect 0 106768 800 106888
rect 0 106496 800 106616
rect 0 106224 800 106344
rect 0 105952 800 106072
rect 0 105680 800 105800
rect 0 105408 800 105528
rect 0 105136 800 105256
rect 0 104864 800 104984
rect 179200 104864 180000 104984
rect 0 104592 800 104712
rect 0 104320 800 104440
rect 0 103912 800 104032
rect 0 103640 800 103760
rect 0 103368 800 103488
rect 0 103096 800 103216
rect 0 102824 800 102944
rect 0 102552 800 102672
rect 0 102280 800 102400
rect 0 102008 800 102128
rect 179200 102144 180000 102264
rect 0 101736 800 101856
rect 0 101464 800 101584
rect 0 101192 800 101312
rect 0 100920 800 101040
rect 0 100648 800 100768
rect 0 100376 800 100496
rect 0 100104 800 100224
rect 0 99696 800 99816
rect 0 99424 800 99544
rect 179200 99424 180000 99544
rect 0 99152 800 99272
rect 0 98880 800 99000
rect 0 98608 800 98728
rect 0 98336 800 98456
rect 0 98064 800 98184
rect 0 97792 800 97912
rect 0 97520 800 97640
rect 0 97248 800 97368
rect 0 96976 800 97096
rect 0 96704 800 96824
rect 179200 96704 180000 96824
rect 0 96432 800 96552
rect 0 96160 800 96280
rect 0 95752 800 95872
rect 0 95480 800 95600
rect 0 95208 800 95328
rect 0 94936 800 95056
rect 0 94664 800 94784
rect 0 94392 800 94512
rect 0 94120 800 94240
rect 0 93848 800 93968
rect 179200 93984 180000 94104
rect 0 93576 800 93696
rect 0 93304 800 93424
rect 0 93032 800 93152
rect 0 92760 800 92880
rect 0 92488 800 92608
rect 0 92216 800 92336
rect 0 91808 800 91928
rect 0 91536 800 91656
rect 0 91264 800 91384
rect 179200 91264 180000 91384
rect 0 90992 800 91112
rect 0 90720 800 90840
rect 0 90448 800 90568
rect 0 90176 800 90296
rect 0 89904 800 90024
rect 0 89632 800 89752
rect 0 89360 800 89480
rect 0 89088 800 89208
rect 0 88816 800 88936
rect 0 88544 800 88664
rect 179200 88544 180000 88664
rect 0 88272 800 88392
rect 0 87864 800 87984
rect 0 87592 800 87712
rect 0 87320 800 87440
rect 0 87048 800 87168
rect 0 86776 800 86896
rect 0 86504 800 86624
rect 0 86232 800 86352
rect 0 85960 800 86080
rect 0 85688 800 85808
rect 179200 85824 180000 85944
rect 0 85416 800 85536
rect 0 85144 800 85264
rect 0 84872 800 84992
rect 0 84600 800 84720
rect 0 84328 800 84448
rect 0 83920 800 84040
rect 0 83648 800 83768
rect 0 83376 800 83496
rect 0 83104 800 83224
rect 179200 83104 180000 83224
rect 0 82832 800 82952
rect 0 82560 800 82680
rect 0 82288 800 82408
rect 0 82016 800 82136
rect 0 81744 800 81864
rect 0 81472 800 81592
rect 0 81200 800 81320
rect 0 80928 800 81048
rect 0 80656 800 80776
rect 0 80384 800 80504
rect 179200 80384 180000 80504
rect 0 80112 800 80232
rect 0 79704 800 79824
rect 0 79432 800 79552
rect 0 79160 800 79280
rect 0 78888 800 79008
rect 0 78616 800 78736
rect 0 78344 800 78464
rect 0 78072 800 78192
rect 0 77800 800 77920
rect 0 77528 800 77648
rect 179200 77664 180000 77784
rect 0 77256 800 77376
rect 0 76984 800 77104
rect 0 76712 800 76832
rect 0 76440 800 76560
rect 0 76168 800 76288
rect 0 75760 800 75880
rect 0 75488 800 75608
rect 0 75216 800 75336
rect 0 74944 800 75064
rect 179200 74944 180000 75064
rect 0 74672 800 74792
rect 0 74400 800 74520
rect 0 74128 800 74248
rect 0 73856 800 73976
rect 0 73584 800 73704
rect 0 73312 800 73432
rect 0 73040 800 73160
rect 0 72768 800 72888
rect 0 72496 800 72616
rect 0 72224 800 72344
rect 179200 72224 180000 72344
rect 0 71816 800 71936
rect 0 71544 800 71664
rect 0 71272 800 71392
rect 0 71000 800 71120
rect 0 70728 800 70848
rect 0 70456 800 70576
rect 0 70184 800 70304
rect 0 69912 800 70032
rect 0 69640 800 69760
rect 0 69368 800 69488
rect 179200 69504 180000 69624
rect 0 69096 800 69216
rect 0 68824 800 68944
rect 0 68552 800 68672
rect 0 68280 800 68400
rect 0 67872 800 67992
rect 0 67600 800 67720
rect 0 67328 800 67448
rect 0 67056 800 67176
rect 0 66784 800 66904
rect 179200 66784 180000 66904
rect 0 66512 800 66632
rect 0 66240 800 66360
rect 0 65968 800 66088
rect 0 65696 800 65816
rect 0 65424 800 65544
rect 0 65152 800 65272
rect 0 64880 800 65000
rect 0 64608 800 64728
rect 0 64336 800 64456
rect 0 63928 800 64048
rect 179200 64064 180000 64184
rect 0 63656 800 63776
rect 0 63384 800 63504
rect 0 63112 800 63232
rect 0 62840 800 62960
rect 0 62568 800 62688
rect 0 62296 800 62416
rect 0 62024 800 62144
rect 0 61752 800 61872
rect 0 61480 800 61600
rect 0 61208 800 61328
rect 179200 61344 180000 61464
rect 0 60936 800 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 0 59712 800 59832
rect 0 59440 800 59560
rect 0 59168 800 59288
rect 0 58896 800 59016
rect 0 58624 800 58744
rect 0 58352 800 58472
rect 179200 58488 180000 58608
rect 0 58080 800 58200
rect 0 57808 800 57928
rect 0 57536 800 57656
rect 0 57264 800 57384
rect 0 56992 800 57112
rect 0 56720 800 56840
rect 0 56448 800 56568
rect 0 56176 800 56296
rect 0 55768 800 55888
rect 179200 55768 180000 55888
rect 0 55496 800 55616
rect 0 55224 800 55344
rect 0 54952 800 55072
rect 0 54680 800 54800
rect 0 54408 800 54528
rect 0 54136 800 54256
rect 0 53864 800 53984
rect 0 53592 800 53712
rect 0 53320 800 53440
rect 0 53048 800 53168
rect 179200 53048 180000 53168
rect 0 52776 800 52896
rect 0 52504 800 52624
rect 0 52232 800 52352
rect 0 51824 800 51944
rect 0 51552 800 51672
rect 0 51280 800 51400
rect 0 51008 800 51128
rect 0 50736 800 50856
rect 0 50464 800 50584
rect 0 50192 800 50312
rect 179200 50328 180000 50448
rect 0 49920 800 50040
rect 0 49648 800 49768
rect 0 49376 800 49496
rect 0 49104 800 49224
rect 0 48832 800 48952
rect 0 48560 800 48680
rect 0 48288 800 48408
rect 0 47880 800 48000
rect 0 47608 800 47728
rect 179200 47608 180000 47728
rect 0 47336 800 47456
rect 0 47064 800 47184
rect 0 46792 800 46912
rect 0 46520 800 46640
rect 0 46248 800 46368
rect 0 45976 800 46096
rect 0 45704 800 45824
rect 0 45432 800 45552
rect 0 45160 800 45280
rect 0 44888 800 45008
rect 179200 44888 180000 45008
rect 0 44616 800 44736
rect 0 44344 800 44464
rect 0 43936 800 44056
rect 0 43664 800 43784
rect 0 43392 800 43512
rect 0 43120 800 43240
rect 0 42848 800 42968
rect 0 42576 800 42696
rect 0 42304 800 42424
rect 0 42032 800 42152
rect 179200 42168 180000 42288
rect 0 41760 800 41880
rect 0 41488 800 41608
rect 0 41216 800 41336
rect 0 40944 800 41064
rect 0 40672 800 40792
rect 0 40400 800 40520
rect 0 40128 800 40248
rect 0 39720 800 39840
rect 0 39448 800 39568
rect 179200 39448 180000 39568
rect 0 39176 800 39296
rect 0 38904 800 39024
rect 0 38632 800 38752
rect 0 38360 800 38480
rect 0 38088 800 38208
rect 0 37816 800 37936
rect 0 37544 800 37664
rect 0 37272 800 37392
rect 0 37000 800 37120
rect 0 36728 800 36848
rect 179200 36728 180000 36848
rect 0 36456 800 36576
rect 0 36184 800 36304
rect 0 35776 800 35896
rect 0 35504 800 35624
rect 0 35232 800 35352
rect 0 34960 800 35080
rect 0 34688 800 34808
rect 0 34416 800 34536
rect 0 34144 800 34264
rect 0 33872 800 33992
rect 179200 34008 180000 34128
rect 0 33600 800 33720
rect 0 33328 800 33448
rect 0 33056 800 33176
rect 0 32784 800 32904
rect 0 32512 800 32632
rect 0 32240 800 32360
rect 0 31832 800 31952
rect 0 31560 800 31680
rect 0 31288 800 31408
rect 179200 31288 180000 31408
rect 0 31016 800 31136
rect 0 30744 800 30864
rect 0 30472 800 30592
rect 0 30200 800 30320
rect 0 29928 800 30048
rect 0 29656 800 29776
rect 0 29384 800 29504
rect 0 29112 800 29232
rect 0 28840 800 28960
rect 0 28568 800 28688
rect 179200 28568 180000 28688
rect 0 28296 800 28416
rect 0 27888 800 28008
rect 0 27616 800 27736
rect 0 27344 800 27464
rect 0 27072 800 27192
rect 0 26800 800 26920
rect 0 26528 800 26648
rect 0 26256 800 26376
rect 0 25984 800 26104
rect 0 25712 800 25832
rect 179200 25848 180000 25968
rect 0 25440 800 25560
rect 0 25168 800 25288
rect 0 24896 800 25016
rect 0 24624 800 24744
rect 0 24352 800 24472
rect 0 23944 800 24064
rect 0 23672 800 23792
rect 0 23400 800 23520
rect 0 23128 800 23248
rect 179200 23128 180000 23248
rect 0 22856 800 22976
rect 0 22584 800 22704
rect 0 22312 800 22432
rect 0 22040 800 22160
rect 0 21768 800 21888
rect 0 21496 800 21616
rect 0 21224 800 21344
rect 0 20952 800 21072
rect 0 20680 800 20800
rect 0 20408 800 20528
rect 179200 20408 180000 20528
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19456 800 19576
rect 0 19184 800 19304
rect 0 18912 800 19032
rect 0 18640 800 18760
rect 0 18368 800 18488
rect 0 18096 800 18216
rect 0 17824 800 17944
rect 0 17552 800 17672
rect 179200 17688 180000 17808
rect 0 17280 800 17400
rect 0 17008 800 17128
rect 0 16736 800 16856
rect 0 16464 800 16584
rect 0 16192 800 16312
rect 0 15784 800 15904
rect 0 15512 800 15632
rect 0 15240 800 15360
rect 0 14968 800 15088
rect 179200 14968 180000 15088
rect 0 14696 800 14816
rect 0 14424 800 14544
rect 0 14152 800 14272
rect 0 13880 800 14000
rect 0 13608 800 13728
rect 0 13336 800 13456
rect 0 13064 800 13184
rect 0 12792 800 12912
rect 0 12520 800 12640
rect 0 12248 800 12368
rect 179200 12248 180000 12368
rect 0 11840 800 11960
rect 0 11568 800 11688
rect 0 11296 800 11416
rect 0 11024 800 11144
rect 0 10752 800 10872
rect 0 10480 800 10600
rect 0 10208 800 10328
rect 0 9936 800 10056
rect 0 9664 800 9784
rect 0 9392 800 9512
rect 179200 9528 180000 9648
rect 0 9120 800 9240
rect 0 8848 800 8968
rect 0 8576 800 8696
rect 0 8304 800 8424
rect 0 7896 800 8016
rect 0 7624 800 7744
rect 0 7352 800 7472
rect 0 7080 800 7200
rect 0 6808 800 6928
rect 179200 6808 180000 6928
rect 0 6536 800 6656
rect 0 6264 800 6384
rect 0 5992 800 6112
rect 0 5720 800 5840
rect 0 5448 800 5568
rect 0 5176 800 5296
rect 0 4904 800 5024
rect 0 4632 800 4752
rect 0 4360 800 4480
rect 0 3952 800 4072
rect 179200 4088 180000 4208
rect 0 3680 800 3800
rect 0 3408 800 3528
rect 0 3136 800 3256
rect 0 2864 800 2984
rect 0 2592 800 2712
rect 0 2320 800 2440
rect 0 2048 800 2168
rect 0 1776 800 1896
rect 0 1504 800 1624
rect 0 1232 800 1352
rect 179200 1368 180000 1488
rect 0 960 800 1080
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
<< obsm3 >>
rect 880 118664 179200 119781
rect 880 118384 179120 118664
rect 880 116072 179200 118384
rect 800 115944 179200 116072
rect 880 115664 179120 115944
rect 880 113224 179200 115664
rect 880 112944 179120 113224
rect 880 112128 179200 112944
rect 800 112000 179200 112128
rect 880 110504 179200 112000
rect 880 110224 179120 110504
rect 880 108184 179200 110224
rect 800 108056 179200 108184
rect 880 107784 179200 108056
rect 880 107504 179120 107784
rect 880 105064 179200 107504
rect 880 104784 179120 105064
rect 880 104240 179200 104784
rect 800 104112 179200 104240
rect 880 102344 179200 104112
rect 880 102064 179120 102344
rect 880 100024 179200 102064
rect 800 99896 179200 100024
rect 880 99624 179200 99896
rect 880 99344 179120 99624
rect 880 96904 179200 99344
rect 880 96624 179120 96904
rect 880 96080 179200 96624
rect 800 95952 179200 96080
rect 880 94184 179200 95952
rect 880 93904 179120 94184
rect 880 92136 179200 93904
rect 800 92008 179200 92136
rect 880 91464 179200 92008
rect 880 91184 179120 91464
rect 880 88744 179200 91184
rect 880 88464 179120 88744
rect 880 88192 179200 88464
rect 800 88064 179200 88192
rect 880 86024 179200 88064
rect 880 85744 179120 86024
rect 880 84248 179200 85744
rect 800 84120 179200 84248
rect 880 83304 179200 84120
rect 880 83024 179120 83304
rect 880 80584 179200 83024
rect 880 80304 179120 80584
rect 880 80032 179200 80304
rect 800 79904 179200 80032
rect 880 77864 179200 79904
rect 880 77584 179120 77864
rect 880 76088 179200 77584
rect 800 75960 179200 76088
rect 880 75144 179200 75960
rect 880 74864 179120 75144
rect 880 72424 179200 74864
rect 880 72144 179120 72424
rect 800 72016 179200 72144
rect 880 69704 179200 72016
rect 880 69424 179120 69704
rect 880 68200 179200 69424
rect 800 68072 179200 68200
rect 880 66984 179200 68072
rect 880 66704 179120 66984
rect 880 64264 179200 66704
rect 880 64256 179120 64264
rect 800 64128 179120 64256
rect 880 63984 179120 64128
rect 880 61544 179200 63984
rect 880 61264 179120 61544
rect 880 60040 179200 61264
rect 800 59912 179200 60040
rect 880 58688 179200 59912
rect 880 58408 179120 58688
rect 880 56096 179200 58408
rect 800 55968 179200 56096
rect 880 55688 179120 55968
rect 880 53248 179200 55688
rect 880 52968 179120 53248
rect 880 52152 179200 52968
rect 800 52024 179200 52152
rect 880 50528 179200 52024
rect 880 50248 179120 50528
rect 880 48208 179200 50248
rect 800 48080 179200 48208
rect 880 47808 179200 48080
rect 880 47528 179120 47808
rect 880 45088 179200 47528
rect 880 44808 179120 45088
rect 880 44264 179200 44808
rect 800 44136 179200 44264
rect 880 42368 179200 44136
rect 880 42088 179120 42368
rect 880 40048 179200 42088
rect 800 39920 179200 40048
rect 880 39648 179200 39920
rect 880 39368 179120 39648
rect 880 36928 179200 39368
rect 880 36648 179120 36928
rect 880 36104 179200 36648
rect 800 35976 179200 36104
rect 880 34208 179200 35976
rect 880 33928 179120 34208
rect 880 32160 179200 33928
rect 800 32032 179200 32160
rect 880 31488 179200 32032
rect 880 31208 179120 31488
rect 880 28768 179200 31208
rect 880 28488 179120 28768
rect 880 28216 179200 28488
rect 800 28088 179200 28216
rect 880 26048 179200 28088
rect 880 25768 179120 26048
rect 880 24272 179200 25768
rect 800 24144 179200 24272
rect 880 23328 179200 24144
rect 880 23048 179120 23328
rect 880 20608 179200 23048
rect 880 20328 179120 20608
rect 880 20056 179200 20328
rect 800 19928 179200 20056
rect 880 17888 179200 19928
rect 880 17608 179120 17888
rect 880 16112 179200 17608
rect 800 15984 179200 16112
rect 880 15168 179200 15984
rect 880 14888 179120 15168
rect 880 12448 179200 14888
rect 880 12168 179120 12448
rect 800 12040 179200 12168
rect 880 9728 179200 12040
rect 880 9448 179120 9728
rect 880 8224 179200 9448
rect 800 8096 179200 8224
rect 880 7008 179200 8096
rect 880 6728 179120 7008
rect 880 4288 179200 6728
rect 880 4280 179120 4288
rect 800 4152 179120 4280
rect 880 4008 179120 4152
rect 880 1568 179200 4008
rect 880 1288 179120 1568
rect 880 171 179200 1288
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< labels >>
rlabel metal2 s 478 119200 534 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 29642 119200 29698 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 32586 119200 32642 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 35438 119200 35494 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 38382 119200 38438 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 41326 119200 41382 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 44270 119200 44326 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 47122 119200 47178 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 50066 119200 50122 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 53010 119200 53066 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 55862 119200 55918 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3330 119200 3386 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 58806 119200 58862 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 61750 119200 61806 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 64694 119200 64750 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 67546 119200 67602 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 70490 119200 70546 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 73434 119200 73490 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 76378 119200 76434 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 79230 119200 79286 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 82174 119200 82230 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 85118 119200 85174 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6274 119200 6330 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 88062 119200 88118 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 90914 119200 90970 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 93858 119200 93914 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 96802 119200 96858 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 99654 119200 99710 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 102598 119200 102654 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 105542 119200 105598 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 108486 119200 108542 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9218 119200 9274 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 12070 119200 12126 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 15014 119200 15070 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 17958 119200 18014 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 20902 119200 20958 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 23754 119200 23810 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 26698 119200 26754 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1398 119200 1454 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 30562 119200 30618 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 33506 119200 33562 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 36450 119200 36506 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 39394 119200 39450 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 42246 119200 42302 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 45190 119200 45246 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 48134 119200 48190 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 51078 119200 51134 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 53930 119200 53986 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 56874 119200 56930 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4342 119200 4398 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 59818 119200 59874 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 62762 119200 62818 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 65614 119200 65670 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 68558 119200 68614 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 71502 119200 71558 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 74354 119200 74410 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 77298 119200 77354 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 80242 119200 80298 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 83186 119200 83242 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 86038 119200 86094 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7286 119200 7342 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 88982 119200 89038 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 91926 119200 91982 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 94870 119200 94926 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 97722 119200 97778 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 100666 119200 100722 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 103610 119200 103666 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 106554 119200 106610 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 109406 119200 109462 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10138 119200 10194 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 13082 119200 13138 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 16026 119200 16082 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 18878 119200 18934 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 21822 119200 21878 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 24766 119200 24822 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 27710 119200 27766 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2410 119200 2466 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 31574 119200 31630 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 34518 119200 34574 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 37370 119200 37426 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 40314 119200 40370 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 43258 119200 43314 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 46202 119200 46258 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 49054 119200 49110 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 51998 119200 52054 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 54942 119200 54998 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 57886 119200 57942 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5262 119200 5318 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 60738 119200 60794 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 63682 119200 63738 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 66626 119200 66682 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 69570 119200 69626 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 72422 119200 72478 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 75366 119200 75422 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 78310 119200 78366 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 81254 119200 81310 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 84106 119200 84162 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8206 119200 8262 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 89994 119200 90050 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 92846 119200 92902 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 95790 119200 95846 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 98734 119200 98790 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 101678 119200 101734 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 104530 119200 104586 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 107474 119200 107530 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 110418 119200 110474 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11150 119200 11206 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 14094 119200 14150 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 16946 119200 17002 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 19890 119200 19946 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 22834 119200 22890 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 25778 119200 25834 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 28630 119200 28686 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 179200 1368 180000 1488 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 134338 0 134394 800 6 irq[1]
port 116 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 0 144 800 264 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 la_data_in[100]
port 119 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 la_data_in[101]
port 120 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 la_data_in[106]
port 125 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 la_data_in[108]
port 127 nsew signal input
rlabel metal3 s 0 92216 800 92336 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 la_data_in[10]
port 129 nsew signal input
rlabel metal3 s 0 93032 800 93152 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 0 95480 800 95600 6 la_data_in[113]
port 133 nsew signal input
rlabel metal3 s 0 96432 800 96552 6 la_data_in[114]
port 134 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 la_data_in[115]
port 135 nsew signal input
rlabel metal3 s 0 98064 800 98184 6 la_data_in[116]
port 136 nsew signal input
rlabel metal3 s 0 98880 800 99000 6 la_data_in[117]
port 137 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 la_data_in[11]
port 140 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 la_data_in[120]
port 141 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 la_data_in[121]
port 142 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 la_data_in[122]
port 143 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 la_data_in[123]
port 144 nsew signal input
rlabel metal3 s 0 104864 800 104984 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal3 s 0 106496 800 106616 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_data_in[12]
port 149 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 0 15240 800 15360 6 la_data_in[18]
port 155 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 la_data_in[19]
port 156 nsew signal input
rlabel metal3 s 0 960 800 1080 6 la_data_in[1]
port 157 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 la_data_in[21]
port 159 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 la_data_in[28]
port 166 nsew signal input
rlabel metal3 s 0 24624 800 24744 6 la_data_in[29]
port 167 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 la_data_in[2]
port 168 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 la_data_in[30]
port 169 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 la_data_in[31]
port 170 nsew signal input
rlabel metal3 s 0 27072 800 27192 6 la_data_in[32]
port 171 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 la_data_in[33]
port 172 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 la_data_in[35]
port 174 nsew signal input
rlabel metal3 s 0 30472 800 30592 6 la_data_in[36]
port 175 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 0 32240 800 32360 6 la_data_in[38]
port 177 nsew signal input
rlabel metal3 s 0 33056 800 33176 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 la_data_in[3]
port 179 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 la_data_in[40]
port 180 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 la_data_in[43]
port 183 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 la_data_in[46]
port 186 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 la_data_in[47]
port 187 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 la_data_in[48]
port 188 nsew signal input
rlabel metal3 s 0 41488 800 41608 6 la_data_in[49]
port 189 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 la_data_in[50]
port 191 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 la_data_in[51]
port 192 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 0 44888 800 45008 6 la_data_in[53]
port 194 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 la_data_in[54]
port 195 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 la_data_in[55]
port 196 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 la_data_in[56]
port 197 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 la_data_in[57]
port 198 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 la_data_in[58]
port 199 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 la_data_in[5]
port 201 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 la_data_in[60]
port 202 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 53320 800 53440 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 la_data_in[64]
port 206 nsew signal input
rlabel metal3 s 0 54952 800 55072 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 la_data_in[66]
port 208 nsew signal input
rlabel metal3 s 0 56720 800 56840 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 57536 800 57656 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 0 58352 800 58472 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 0 5176 800 5296 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 la_data_in[71]
port 214 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 la_data_in[72]
port 215 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 la_data_in[73]
port 216 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_data_in[74]
port 217 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 la_data_in[75]
port 218 nsew signal input
rlabel metal3 s 0 64336 800 64456 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 0 65152 800 65272 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 0 66784 800 66904 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 0 5992 800 6112 6 la_data_in[7]
port 223 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 la_data_in[82]
port 226 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 la_data_in[84]
port 228 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 74400 800 74520 6 la_data_in[88]
port 232 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 la_data_in[89]
port 233 nsew signal input
rlabel metal3 s 0 6808 800 6928 6 la_data_in[8]
port 234 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 la_data_in[90]
port 235 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 la_data_in[92]
port 237 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 la_data_in[93]
port 238 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 la_data_in[99]
port 244 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 416 800 536 6 la_data_out[0]
port 246 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 86504 800 86624 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 0 88272 800 88392 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 89088 800 89208 6 la_data_out[105]
port 252 nsew signal output
rlabel metal3 s 0 89904 800 90024 6 la_data_out[106]
port 253 nsew signal output
rlabel metal3 s 0 90720 800 90840 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 0 91536 800 91656 6 la_data_out[108]
port 255 nsew signal output
rlabel metal3 s 0 92488 800 92608 6 la_data_out[109]
port 256 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 la_data_out[10]
port 257 nsew signal output
rlabel metal3 s 0 93304 800 93424 6 la_data_out[110]
port 258 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 la_data_out[111]
port 259 nsew signal output
rlabel metal3 s 0 94936 800 95056 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 95752 800 95872 6 la_data_out[113]
port 261 nsew signal output
rlabel metal3 s 0 96704 800 96824 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 0 97520 800 97640 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 0 98336 800 98456 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 99152 800 99272 6 la_data_out[117]
port 265 nsew signal output
rlabel metal3 s 0 100104 800 100224 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 100920 800 101040 6 la_data_out[119]
port 267 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 0 101736 800 101856 6 la_data_out[120]
port 269 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 la_data_out[121]
port 270 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 0 104320 800 104440 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 105136 800 105256 6 la_data_out[124]
port 273 nsew signal output
rlabel metal3 s 0 105952 800 106072 6 la_data_out[125]
port 274 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 107584 800 107704 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 0 11296 800 11416 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 la_data_out[15]
port 280 nsew signal output
rlabel metal3 s 0 13880 800 14000 6 la_data_out[16]
port 281 nsew signal output
rlabel metal3 s 0 14696 800 14816 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 0 15512 800 15632 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 16464 800 16584 6 la_data_out[19]
port 284 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 18096 800 18216 6 la_data_out[21]
port 287 nsew signal output
rlabel metal3 s 0 18912 800 19032 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 la_data_out[23]
port 289 nsew signal output
rlabel metal3 s 0 20680 800 20800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 22312 800 22432 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 la_data_out[27]
port 293 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 0 24896 800 25016 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 la_data_out[2]
port 296 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 la_data_out[31]
port 298 nsew signal output
rlabel metal3 s 0 27344 800 27464 6 la_data_out[32]
port 299 nsew signal output
rlabel metal3 s 0 28296 800 28416 6 la_data_out[33]
port 300 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 la_data_out[34]
port 301 nsew signal output
rlabel metal3 s 0 29928 800 30048 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 30744 800 30864 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 la_data_out[37]
port 304 nsew signal output
rlabel metal3 s 0 32512 800 32632 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 0 33328 800 33448 6 la_data_out[39]
port 306 nsew signal output
rlabel metal3 s 0 2864 800 2984 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 la_data_out[40]
port 308 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 la_data_out[41]
port 309 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 la_data_out[42]
port 310 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 la_data_out[43]
port 311 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 la_data_out[45]
port 313 nsew signal output
rlabel metal3 s 0 39176 800 39296 6 la_data_out[46]
port 314 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 40944 800 41064 6 la_data_out[48]
port 316 nsew signal output
rlabel metal3 s 0 41760 800 41880 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 3680 800 3800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 la_data_out[50]
port 319 nsew signal output
rlabel metal3 s 0 43392 800 43512 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 la_data_out[56]
port 325 nsew signal output
rlabel metal3 s 0 48560 800 48680 6 la_data_out[57]
port 326 nsew signal output
rlabel metal3 s 0 49376 800 49496 6 la_data_out[58]
port 327 nsew signal output
rlabel metal3 s 0 50192 800 50312 6 la_data_out[59]
port 328 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 la_data_out[5]
port 329 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 la_data_out[60]
port 330 nsew signal output
rlabel metal3 s 0 51824 800 51944 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 0 52776 800 52896 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 0 53592 800 53712 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 0 54408 800 54528 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 0 55224 800 55344 6 la_data_out[65]
port 335 nsew signal output
rlabel metal3 s 0 56176 800 56296 6 la_data_out[66]
port 336 nsew signal output
rlabel metal3 s 0 56992 800 57112 6 la_data_out[67]
port 337 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 la_data_out[68]
port 338 nsew signal output
rlabel metal3 s 0 58624 800 58744 6 la_data_out[69]
port 339 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 la_data_out[6]
port 340 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 la_data_out[71]
port 342 nsew signal output
rlabel metal3 s 0 61208 800 61328 6 la_data_out[72]
port 343 nsew signal output
rlabel metal3 s 0 62024 800 62144 6 la_data_out[73]
port 344 nsew signal output
rlabel metal3 s 0 62840 800 62960 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 0 63656 800 63776 6 la_data_out[75]
port 346 nsew signal output
rlabel metal3 s 0 64608 800 64728 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 0 65424 800 65544 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 la_data_out[78]
port 349 nsew signal output
rlabel metal3 s 0 67056 800 67176 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 0 6264 800 6384 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 la_data_out[80]
port 352 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 la_data_out[81]
port 353 nsew signal output
rlabel metal3 s 0 69640 800 69760 6 la_data_out[82]
port 354 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 71272 800 71392 6 la_data_out[84]
port 356 nsew signal output
rlabel metal3 s 0 72224 800 72344 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 0 73040 800 73160 6 la_data_out[86]
port 358 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 la_data_out[87]
port 359 nsew signal output
rlabel metal3 s 0 74672 800 74792 6 la_data_out[88]
port 360 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 la_data_out[89]
port 361 nsew signal output
rlabel metal3 s 0 7080 800 7200 6 la_data_out[8]
port 362 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 la_data_out[90]
port 363 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 la_data_out[91]
port 364 nsew signal output
rlabel metal3 s 0 78072 800 78192 6 la_data_out[92]
port 365 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 la_data_out[93]
port 366 nsew signal output
rlabel metal3 s 0 79704 800 79824 6 la_data_out[94]
port 367 nsew signal output
rlabel metal3 s 0 80656 800 80776 6 la_data_out[95]
port 368 nsew signal output
rlabel metal3 s 0 81472 800 81592 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 82288 800 82408 6 la_data_out[97]
port 370 nsew signal output
rlabel metal3 s 0 83104 800 83224 6 la_data_out[98]
port 371 nsew signal output
rlabel metal3 s 0 83920 800 84040 6 la_data_out[99]
port 372 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 la_data_out[9]
port 373 nsew signal output
rlabel metal3 s 0 688 800 808 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 0 85144 800 85264 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 la_oenb[101]
port 376 nsew signal input
rlabel metal3 s 0 86776 800 86896 6 la_oenb[102]
port 377 nsew signal input
rlabel metal3 s 0 87592 800 87712 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 0 88544 800 88664 6 la_oenb[104]
port 379 nsew signal input
rlabel metal3 s 0 89360 800 89480 6 la_oenb[105]
port 380 nsew signal input
rlabel metal3 s 0 90176 800 90296 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 0 90992 800 91112 6 la_oenb[107]
port 382 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 la_oenb[108]
port 383 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 la_oenb[109]
port 384 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 la_oenb[110]
port 386 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 la_oenb[112]
port 388 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 la_oenb[113]
port 389 nsew signal input
rlabel metal3 s 0 96976 800 97096 6 la_oenb[114]
port 390 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 la_oenb[115]
port 391 nsew signal input
rlabel metal3 s 0 98608 800 98728 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 0 9936 800 10056 6 la_oenb[11]
port 396 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 la_oenb[120]
port 397 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 0 104592 800 104712 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 106224 800 106344 6 la_oenb[125]
port 402 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 0 107856 800 107976 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 0 10752 800 10872 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 12520 800 12640 6 la_oenb[14]
port 407 nsew signal input
rlabel metal3 s 0 13336 800 13456 6 la_oenb[15]
port 408 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 la_oenb[17]
port 410 nsew signal input
rlabel metal3 s 0 15784 800 15904 6 la_oenb[18]
port 411 nsew signal input
rlabel metal3 s 0 16736 800 16856 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 la_oenb[21]
port 415 nsew signal input
rlabel metal3 s 0 19184 800 19304 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 la_oenb[23]
port 417 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 la_oenb[24]
port 418 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 la_oenb[25]
port 419 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 la_oenb[27]
port 421 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 la_oenb[28]
port 422 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 la_oenb[30]
port 425 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 la_oenb[31]
port 426 nsew signal input
rlabel metal3 s 0 27616 800 27736 6 la_oenb[32]
port 427 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 0 29384 800 29504 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 la_oenb[36]
port 431 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 0 32784 800 32904 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 la_oenb[39]
port 434 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 la_oenb[40]
port 436 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 la_oenb[41]
port 437 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 la_oenb[44]
port 440 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 la_oenb[45]
port 441 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_oenb[46]
port 442 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 0 41216 800 41336 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 0 42032 800 42152 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 la_oenb[4]
port 446 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_oenb[50]
port 447 nsew signal input
rlabel metal3 s 0 43664 800 43784 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 44616 800 44736 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 0 45432 800 45552 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 la_oenb[54]
port 451 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 la_oenb[57]
port 454 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 0 50464 800 50584 6 la_oenb[59]
port 456 nsew signal input
rlabel metal3 s 0 4904 800 5024 6 la_oenb[5]
port 457 nsew signal input
rlabel metal3 s 0 51280 800 51400 6 la_oenb[60]
port 458 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 la_oenb[61]
port 459 nsew signal input
rlabel metal3 s 0 53048 800 53168 6 la_oenb[62]
port 460 nsew signal input
rlabel metal3 s 0 53864 800 53984 6 la_oenb[63]
port 461 nsew signal input
rlabel metal3 s 0 54680 800 54800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 la_oenb[65]
port 463 nsew signal input
rlabel metal3 s 0 56448 800 56568 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 0 58080 800 58200 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 58896 800 59016 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 la_oenb[73]
port 472 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 la_oenb[74]
port 473 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 la_oenb[75]
port 474 nsew signal input
rlabel metal3 s 0 64880 800 65000 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 0 66512 800 66632 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 6536 800 6656 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 la_oenb[82]
port 482 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 la_oenb[84]
port 484 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_oenb[87]
port 487 nsew signal input
rlabel metal3 s 0 74944 800 75064 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 0 75760 800 75880 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 0 7352 800 7472 6 la_oenb[8]
port 490 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 la_oenb[91]
port 492 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 la_oenb[93]
port 494 nsew signal input
rlabel metal3 s 0 80112 800 80232 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 la_oenb[95]
port 496 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 la_oenb[96]
port 497 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 la_oenb[99]
port 500 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 mem1_data_i[0]
port 502 nsew signal input
rlabel metal3 s 0 113568 800 113688 6 mem1_data_i[10]
port 503 nsew signal input
rlabel metal2 s 153106 0 153162 800 6 mem1_data_i[11]
port 504 nsew signal input
rlabel metal3 s 179200 64064 180000 64184 6 mem1_data_i[12]
port 505 nsew signal input
rlabel metal3 s 179200 72224 180000 72344 6 mem1_data_i[13]
port 506 nsew signal input
rlabel metal2 s 163962 119200 164018 120000 6 mem1_data_i[14]
port 507 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 mem1_data_i[15]
port 508 nsew signal input
rlabel metal2 s 165894 119200 165950 120000 6 mem1_data_i[16]
port 509 nsew signal input
rlabel metal3 s 0 114928 800 115048 6 mem1_data_i[17]
port 510 nsew signal input
rlabel metal3 s 0 115200 800 115320 6 mem1_data_i[18]
port 511 nsew signal input
rlabel metal2 s 163042 0 163098 800 6 mem1_data_i[19]
port 512 nsew signal input
rlabel metal3 s 179200 14968 180000 15088 6 mem1_data_i[1]
port 513 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 mem1_data_i[20]
port 514 nsew signal input
rlabel metal3 s 179200 93984 180000 94104 6 mem1_data_i[21]
port 515 nsew signal input
rlabel metal3 s 179200 96704 180000 96824 6 mem1_data_i[22]
port 516 nsew signal input
rlabel metal3 s 0 117512 800 117632 6 mem1_data_i[23]
port 517 nsew signal input
rlabel metal2 s 169298 0 169354 800 6 mem1_data_i[24]
port 518 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 mem1_data_i[25]
port 519 nsew signal input
rlabel metal3 s 179200 104864 180000 104984 6 mem1_data_i[26]
port 520 nsew signal input
rlabel metal2 s 173070 0 173126 800 6 mem1_data_i[27]
port 521 nsew signal input
rlabel metal2 s 174358 0 174414 800 6 mem1_data_i[28]
port 522 nsew signal input
rlabel metal3 s 179200 113024 180000 113144 6 mem1_data_i[29]
port 523 nsew signal input
rlabel metal2 s 151266 119200 151322 120000 6 mem1_data_i[2]
port 524 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 mem1_data_i[30]
port 525 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 mem1_data_i[31]
port 526 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 mem1_data_i[3]
port 527 nsew signal input
rlabel metal2 s 155130 119200 155186 120000 6 mem1_data_i[4]
port 528 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 mem1_data_i[5]
port 529 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 mem1_data_i[6]
port 530 nsew signal input
rlabel metal3 s 179200 44888 180000 45008 6 mem1_data_i[7]
port 531 nsew signal input
rlabel metal3 s 0 113024 800 113144 6 mem1_data_i[8]
port 532 nsew signal input
rlabel metal2 s 160006 119200 160062 120000 6 mem1_data_i[9]
port 533 nsew signal input
rlabel metal3 s 179200 4088 180000 4208 6 mem_data2_i[0]
port 534 nsew signal input
rlabel metal2 s 150530 0 150586 800 6 mem_data2_i[10]
port 535 nsew signal input
rlabel metal3 s 179200 61344 180000 61464 6 mem_data2_i[11]
port 536 nsew signal input
rlabel metal3 s 0 113840 800 113960 6 mem_data2_i[12]
port 537 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 mem_data2_i[13]
port 538 nsew signal input
rlabel metal2 s 164882 119200 164938 120000 6 mem_data2_i[14]
port 539 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 mem_data2_i[15]
port 540 nsew signal input
rlabel metal2 s 160558 0 160614 800 6 mem_data2_i[16]
port 541 nsew signal input
rlabel metal3 s 179200 83104 180000 83224 6 mem_data2_i[17]
port 542 nsew signal input
rlabel metal3 s 0 115472 800 115592 6 mem_data2_i[18]
port 543 nsew signal input
rlabel metal3 s 0 116152 800 116272 6 mem_data2_i[19]
port 544 nsew signal input
rlabel metal2 s 146390 119200 146446 120000 6 mem_data2_i[1]
port 545 nsew signal input
rlabel metal3 s 179200 91264 180000 91384 6 mem_data2_i[20]
port 546 nsew signal input
rlabel metal2 s 167826 119200 167882 120000 6 mem_data2_i[21]
port 547 nsew signal input
rlabel metal3 s 179200 99424 180000 99544 6 mem_data2_i[22]
port 548 nsew signal input
rlabel metal3 s 179200 102144 180000 102264 6 mem_data2_i[23]
port 549 nsew signal input
rlabel metal2 s 171690 119200 171746 120000 6 mem_data2_i[24]
port 550 nsew signal input
rlabel metal2 s 174634 119200 174690 120000 6 mem_data2_i[25]
port 551 nsew signal input
rlabel metal2 s 170586 0 170642 800 6 mem_data2_i[26]
port 552 nsew signal input
rlabel metal3 s 179200 107584 180000 107704 6 mem_data2_i[27]
port 553 nsew signal input
rlabel metal2 s 175646 119200 175702 120000 6 mem_data2_i[28]
port 554 nsew signal input
rlabel metal2 s 175554 0 175610 800 6 mem_data2_i[29]
port 555 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 mem_data2_i[2]
port 556 nsew signal input
rlabel metal3 s 179200 115744 180000 115864 6 mem_data2_i[30]
port 557 nsew signal input
rlabel metal2 s 179510 119200 179566 120000 6 mem_data2_i[31]
port 558 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 mem_data2_i[3]
port 559 nsew signal input
rlabel metal3 s 179200 31288 180000 31408 6 mem_data2_i[4]
port 560 nsew signal input
rlabel metal3 s 179200 36728 180000 36848 6 mem_data2_i[5]
port 561 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 mem_data2_i[6]
port 562 nsew signal input
rlabel metal2 s 159086 119200 159142 120000 6 mem_data2_i[7]
port 563 nsew signal input
rlabel metal3 s 179200 50328 180000 50448 6 mem_data2_i[8]
port 564 nsew signal input
rlabel metal2 s 161018 119200 161074 120000 6 mem_data2_i[9]
port 565 nsew signal input
rlabel metal3 s 179200 6808 180000 6928 6 mem_data_i[0]
port 566 nsew signal input
rlabel metal2 s 151818 0 151874 800 6 mem_data_i[10]
port 567 nsew signal input
rlabel metal2 s 162950 119200 163006 120000 6 mem_data_i[11]
port 568 nsew signal input
rlabel metal3 s 179200 66784 180000 66904 6 mem_data_i[12]
port 569 nsew signal input
rlabel metal3 s 179200 74944 180000 75064 6 mem_data_i[13]
port 570 nsew signal input
rlabel metal3 s 179200 80384 180000 80504 6 mem_data_i[14]
port 571 nsew signal input
rlabel metal2 s 158074 0 158130 800 6 mem_data_i[15]
port 572 nsew signal input
rlabel metal3 s 0 114656 800 114776 6 mem_data_i[16]
port 573 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 mem_data_i[17]
port 574 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 mem_data_i[18]
port 575 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 mem_data_i[19]
port 576 nsew signal input
rlabel metal2 s 147402 119200 147458 120000 6 mem_data_i[1]
port 577 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 mem_data_i[20]
port 578 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 mem_data_i[21]
port 579 nsew signal input
rlabel metal2 s 168102 0 168158 800 6 mem_data_i[22]
port 580 nsew signal input
rlabel metal2 s 169758 119200 169814 120000 6 mem_data_i[23]
port 581 nsew signal input
rlabel metal2 s 172702 119200 172758 120000 6 mem_data_i[24]
port 582 nsew signal input
rlabel metal3 s 0 118056 800 118176 6 mem_data_i[25]
port 583 nsew signal input
rlabel metal2 s 171782 0 171838 800 6 mem_data_i[26]
port 584 nsew signal input
rlabel metal3 s 0 118872 800 118992 6 mem_data_i[27]
port 585 nsew signal input
rlabel metal2 s 176566 119200 176622 120000 6 mem_data_i[28]
port 586 nsew signal input
rlabel metal2 s 176842 0 176898 800 6 mem_data_i[29]
port 587 nsew signal input
rlabel metal2 s 152278 119200 152334 120000 6 mem_data_i[2]
port 588 nsew signal input
rlabel metal3 s 179200 118464 180000 118584 6 mem_data_i[30]
port 589 nsew signal input
rlabel metal2 s 179326 0 179382 800 6 mem_data_i[31]
port 590 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 mem_data_i[3]
port 591 nsew signal input
rlabel metal3 s 179200 34008 180000 34128 6 mem_data_i[4]
port 592 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 mem_data_i[5]
port 593 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 mem_data_i[6]
port 594 nsew signal input
rlabel metal2 s 143078 0 143134 800 6 mem_data_i[7]
port 595 nsew signal input
rlabel metal2 s 145562 0 145618 800 6 mem_data_i[8]
port 596 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 mem_data_i[9]
port 597 nsew signal input
rlabel metal2 s 143538 119200 143594 120000 6 mem_data_o[0]
port 598 nsew signal output
rlabel metal3 s 179200 58488 180000 58608 6 mem_data_o[10]
port 599 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 mem_data_o[11]
port 600 nsew signal output
rlabel metal3 s 179200 69504 180000 69624 6 mem_data_o[12]
port 601 nsew signal output
rlabel metal3 s 179200 77664 180000 77784 6 mem_data_o[13]
port 602 nsew signal output
rlabel metal2 s 156786 0 156842 800 6 mem_data_o[14]
port 603 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 mem_data_o[15]
port 604 nsew signal output
rlabel metal2 s 166814 119200 166870 120000 6 mem_data_o[16]
port 605 nsew signal output
rlabel metal3 s 179200 85824 180000 85944 6 mem_data_o[17]
port 606 nsew signal output
rlabel metal3 s 179200 88544 180000 88664 6 mem_data_o[18]
port 607 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 mem_data_o[19]
port 608 nsew signal output
rlabel metal2 s 148322 119200 148378 120000 6 mem_data_o[1]
port 609 nsew signal output
rlabel metal2 s 165526 0 165582 800 6 mem_data_o[20]
port 610 nsew signal output
rlabel metal2 s 166814 0 166870 800 6 mem_data_o[21]
port 611 nsew signal output
rlabel metal2 s 168838 119200 168894 120000 6 mem_data_o[22]
port 612 nsew signal output
rlabel metal2 s 170770 119200 170826 120000 6 mem_data_o[23]
port 613 nsew signal output
rlabel metal2 s 173622 119200 173678 120000 6 mem_data_o[24]
port 614 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 mem_data_o[25]
port 615 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 mem_data_o[26]
port 616 nsew signal output
rlabel metal3 s 179200 110304 180000 110424 6 mem_data_o[27]
port 617 nsew signal output
rlabel metal2 s 177578 119200 177634 120000 6 mem_data_o[28]
port 618 nsew signal output
rlabel metal2 s 178038 0 178094 800 6 mem_data_o[29]
port 619 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 mem_data_o[2]
port 620 nsew signal output
rlabel metal2 s 178498 119200 178554 120000 6 mem_data_o[30]
port 621 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 mem_data_o[31]
port 622 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 mem_data_o[3]
port 623 nsew signal output
rlabel metal2 s 156142 119200 156198 120000 6 mem_data_o[4]
port 624 nsew signal output
rlabel metal3 s 179200 39448 180000 39568 6 mem_data_o[5]
port 625 nsew signal output
rlabel metal2 s 158074 119200 158130 120000 6 mem_data_o[6]
port 626 nsew signal output
rlabel metal3 s 0 112752 800 112872 6 mem_data_o[7]
port 627 nsew signal output
rlabel metal3 s 0 113296 800 113416 6 mem_data_o[8]
port 628 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 mem_data_o[9]
port 629 nsew signal output
rlabel metal2 s 144458 119200 144514 120000 6 mem_raddr_o[0]
port 630 nsew signal output
rlabel metal3 s 179200 17688 180000 17808 6 mem_raddr_o[1]
port 631 nsew signal output
rlabel metal3 s 179200 23128 180000 23248 6 mem_raddr_o[2]
port 632 nsew signal output
rlabel metal2 s 154210 119200 154266 120000 6 mem_raddr_o[3]
port 633 nsew signal output
rlabel metal2 s 157154 119200 157210 120000 6 mem_raddr_o[4]
port 634 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 mem_raddr_o[5]
port 635 nsew signal output
rlabel metal3 s 0 112480 800 112600 6 mem_raddr_o[6]
port 636 nsew signal output
rlabel metal3 s 179200 47608 180000 47728 6 mem_raddr_o[7]
port 637 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 mem_raddr_o[8]
port 638 nsew signal output
rlabel metal2 s 162030 119200 162086 120000 6 mem_raddr_o[9]
port 639 nsew signal output
rlabel metal3 s 179200 9528 180000 9648 6 mem_renb_o[0]
port 640 nsew signal output
rlabel metal2 s 149334 119200 149390 120000 6 mem_renb_o[1]
port 641 nsew signal output
rlabel metal3 s 0 108264 800 108384 6 mem_waddr_o[0]
port 642 nsew signal output
rlabel metal3 s 179200 20408 180000 20528 6 mem_waddr_o[1]
port 643 nsew signal output
rlabel metal2 s 153198 119200 153254 120000 6 mem_waddr_o[2]
port 644 nsew signal output
rlabel metal2 s 138018 0 138074 800 6 mem_waddr_o[3]
port 645 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 mem_waddr_o[4]
port 646 nsew signal output
rlabel metal3 s 0 111256 800 111376 6 mem_waddr_o[5]
port 647 nsew signal output
rlabel metal3 s 179200 42168 180000 42288 6 mem_waddr_o[6]
port 648 nsew signal output
rlabel metal2 s 144274 0 144330 800 6 mem_waddr_o[7]
port 649 nsew signal output
rlabel metal3 s 179200 53048 180000 53168 6 mem_waddr_o[8]
port 650 nsew signal output
rlabel metal3 s 179200 55768 180000 55888 6 mem_waddr_o[9]
port 651 nsew signal output
rlabel metal3 s 179200 12248 180000 12368 6 mem_wenb_o[0]
port 652 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 mem_wenb_o[1]
port 653 nsew signal output
rlabel metal2 s 111338 119200 111394 120000 6 phase0_in[0]
port 654 nsew signal input
rlabel metal2 s 140594 119200 140650 120000 6 phase0_in[10]
port 655 nsew signal input
rlabel metal2 s 114282 119200 114338 120000 6 phase0_in[1]
port 656 nsew signal input
rlabel metal2 s 117226 119200 117282 120000 6 phase0_in[2]
port 657 nsew signal input
rlabel metal2 s 120170 119200 120226 120000 6 phase0_in[3]
port 658 nsew signal input
rlabel metal2 s 123022 119200 123078 120000 6 phase0_in[4]
port 659 nsew signal input
rlabel metal2 s 125966 119200 126022 120000 6 phase0_in[5]
port 660 nsew signal input
rlabel metal2 s 128910 119200 128966 120000 6 phase0_in[6]
port 661 nsew signal input
rlabel metal2 s 131854 119200 131910 120000 6 phase0_in[7]
port 662 nsew signal input
rlabel metal2 s 134706 119200 134762 120000 6 phase0_in[8]
port 663 nsew signal input
rlabel metal2 s 137650 119200 137706 120000 6 phase0_in[9]
port 664 nsew signal input
rlabel metal2 s 112350 119200 112406 120000 6 phase1_in[0]
port 665 nsew signal input
rlabel metal2 s 141514 119200 141570 120000 6 phase1_in[10]
port 666 nsew signal input
rlabel metal2 s 115294 119200 115350 120000 6 phase1_in[1]
port 667 nsew signal input
rlabel metal2 s 118146 119200 118202 120000 6 phase1_in[2]
port 668 nsew signal input
rlabel metal2 s 121090 119200 121146 120000 6 phase1_in[3]
port 669 nsew signal input
rlabel metal2 s 124034 119200 124090 120000 6 phase1_in[4]
port 670 nsew signal input
rlabel metal2 s 126978 119200 127034 120000 6 phase1_in[5]
port 671 nsew signal input
rlabel metal2 s 129830 119200 129886 120000 6 phase1_in[6]
port 672 nsew signal input
rlabel metal2 s 132774 119200 132830 120000 6 phase1_in[7]
port 673 nsew signal input
rlabel metal2 s 135718 119200 135774 120000 6 phase1_in[8]
port 674 nsew signal input
rlabel metal2 s 138662 119200 138718 120000 6 phase1_in[9]
port 675 nsew signal input
rlabel metal2 s 113362 119200 113418 120000 6 phase2_in[0]
port 676 nsew signal input
rlabel metal2 s 142526 119200 142582 120000 6 phase2_in[10]
port 677 nsew signal input
rlabel metal2 s 116214 119200 116270 120000 6 phase2_in[1]
port 678 nsew signal input
rlabel metal2 s 119158 119200 119214 120000 6 phase2_in[2]
port 679 nsew signal input
rlabel metal2 s 122102 119200 122158 120000 6 phase2_in[3]
port 680 nsew signal input
rlabel metal2 s 125046 119200 125102 120000 6 phase2_in[4]
port 681 nsew signal input
rlabel metal2 s 127898 119200 127954 120000 6 phase2_in[5]
port 682 nsew signal input
rlabel metal2 s 130842 119200 130898 120000 6 phase2_in[6]
port 683 nsew signal input
rlabel metal2 s 133786 119200 133842 120000 6 phase2_in[7]
port 684 nsew signal input
rlabel metal2 s 136638 119200 136694 120000 6 phase2_in[8]
port 685 nsew signal input
rlabel metal2 s 139582 119200 139638 120000 6 phase2_in[9]
port 686 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 vco_enb_o[0]
port 687 nsew signal output
rlabel metal2 s 135534 0 135590 800 6 vco_enb_o[1]
port 688 nsew signal output
rlabel metal3 s 179200 25848 180000 25968 6 vco_enb_o[2]
port 689 nsew signal output
rlabel metal2 s 570 0 626 800 6 wb_clk_i
port 690 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 wb_rst_i
port 691 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_ack_o
port 692 nsew signal output
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[0]
port 693 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 wbs_adr_i[10]
port 694 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 wbs_adr_i[11]
port 695 nsew signal input
rlabel metal2 s 58070 0 58126 800 6 wbs_adr_i[12]
port 696 nsew signal input
rlabel metal2 s 61750 0 61806 800 6 wbs_adr_i[13]
port 697 nsew signal input
rlabel metal2 s 65522 0 65578 800 6 wbs_adr_i[14]
port 698 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_adr_i[15]
port 699 nsew signal input
rlabel metal2 s 73066 0 73122 800 6 wbs_adr_i[16]
port 700 nsew signal input
rlabel metal2 s 76838 0 76894 800 6 wbs_adr_i[17]
port 701 nsew signal input
rlabel metal2 s 80518 0 80574 800 6 wbs_adr_i[18]
port 702 nsew signal input
rlabel metal2 s 84290 0 84346 800 6 wbs_adr_i[19]
port 703 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[1]
port 704 nsew signal input
rlabel metal2 s 88062 0 88118 800 6 wbs_adr_i[20]
port 705 nsew signal input
rlabel metal2 s 91834 0 91890 800 6 wbs_adr_i[21]
port 706 nsew signal input
rlabel metal2 s 95514 0 95570 800 6 wbs_adr_i[22]
port 707 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 wbs_adr_i[23]
port 708 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 wbs_adr_i[24]
port 709 nsew signal input
rlabel metal2 s 106830 0 106886 800 6 wbs_adr_i[25]
port 710 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 wbs_adr_i[26]
port 711 nsew signal input
rlabel metal2 s 114282 0 114338 800 6 wbs_adr_i[27]
port 712 nsew signal input
rlabel metal2 s 118054 0 118110 800 6 wbs_adr_i[28]
port 713 nsew signal input
rlabel metal2 s 121826 0 121882 800 6 wbs_adr_i[29]
port 714 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 wbs_adr_i[2]
port 715 nsew signal input
rlabel metal2 s 125598 0 125654 800 6 wbs_adr_i[30]
port 716 nsew signal input
rlabel metal2 s 129278 0 129334 800 6 wbs_adr_i[31]
port 717 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 wbs_adr_i[3]
port 718 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 wbs_adr_i[4]
port 719 nsew signal input
rlabel metal2 s 31758 0 31814 800 6 wbs_adr_i[5]
port 720 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 wbs_adr_i[6]
port 721 nsew signal input
rlabel metal2 s 39302 0 39358 800 6 wbs_adr_i[7]
port 722 nsew signal input
rlabel metal2 s 43074 0 43130 800 6 wbs_adr_i[8]
port 723 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 wbs_adr_i[9]
port 724 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_cyc_i
port 725 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[0]
port 726 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 wbs_dat_i[10]
port 727 nsew signal input
rlabel metal2 s 55494 0 55550 800 6 wbs_dat_i[11]
port 728 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_dat_i[12]
port 729 nsew signal input
rlabel metal2 s 63038 0 63094 800 6 wbs_dat_i[13]
port 730 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_dat_i[14]
port 731 nsew signal input
rlabel metal2 s 70582 0 70638 800 6 wbs_dat_i[15]
port 732 nsew signal input
rlabel metal2 s 74262 0 74318 800 6 wbs_dat_i[16]
port 733 nsew signal input
rlabel metal2 s 78034 0 78090 800 6 wbs_dat_i[17]
port 734 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 wbs_dat_i[18]
port 735 nsew signal input
rlabel metal2 s 85578 0 85634 800 6 wbs_dat_i[19]
port 736 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_dat_i[1]
port 737 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 wbs_dat_i[20]
port 738 nsew signal input
rlabel metal2 s 93030 0 93086 800 6 wbs_dat_i[21]
port 739 nsew signal input
rlabel metal2 s 96802 0 96858 800 6 wbs_dat_i[22]
port 740 nsew signal input
rlabel metal2 s 100574 0 100630 800 6 wbs_dat_i[23]
port 741 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 wbs_dat_i[24]
port 742 nsew signal input
rlabel metal2 s 108026 0 108082 800 6 wbs_dat_i[25]
port 743 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 wbs_dat_i[26]
port 744 nsew signal input
rlabel metal2 s 115570 0 115626 800 6 wbs_dat_i[27]
port 745 nsew signal input
rlabel metal2 s 119342 0 119398 800 6 wbs_dat_i[28]
port 746 nsew signal input
rlabel metal2 s 123022 0 123078 800 6 wbs_dat_i[29]
port 747 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_i[2]
port 748 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 wbs_dat_i[30]
port 749 nsew signal input
rlabel metal2 s 130566 0 130622 800 6 wbs_dat_i[31]
port 750 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_i[3]
port 751 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_dat_i[4]
port 752 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[5]
port 753 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 wbs_dat_i[6]
port 754 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 wbs_dat_i[7]
port 755 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_i[8]
port 756 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 wbs_dat_i[9]
port 757 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_o[0]
port 758 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 wbs_dat_o[10]
port 759 nsew signal output
rlabel metal2 s 56782 0 56838 800 6 wbs_dat_o[11]
port 760 nsew signal output
rlabel metal2 s 60554 0 60610 800 6 wbs_dat_o[12]
port 761 nsew signal output
rlabel metal2 s 64326 0 64382 800 6 wbs_dat_o[13]
port 762 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 wbs_dat_o[14]
port 763 nsew signal output
rlabel metal2 s 71778 0 71834 800 6 wbs_dat_o[15]
port 764 nsew signal output
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_o[16]
port 765 nsew signal output
rlabel metal2 s 79322 0 79378 800 6 wbs_dat_o[17]
port 766 nsew signal output
rlabel metal2 s 83002 0 83058 800 6 wbs_dat_o[18]
port 767 nsew signal output
rlabel metal2 s 86774 0 86830 800 6 wbs_dat_o[19]
port 768 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_dat_o[1]
port 769 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 wbs_dat_o[20]
port 770 nsew signal output
rlabel metal2 s 94318 0 94374 800 6 wbs_dat_o[21]
port 771 nsew signal output
rlabel metal2 s 98090 0 98146 800 6 wbs_dat_o[22]
port 772 nsew signal output
rlabel metal2 s 101770 0 101826 800 6 wbs_dat_o[23]
port 773 nsew signal output
rlabel metal2 s 105542 0 105598 800 6 wbs_dat_o[24]
port 774 nsew signal output
rlabel metal2 s 109314 0 109370 800 6 wbs_dat_o[25]
port 775 nsew signal output
rlabel metal2 s 113086 0 113142 800 6 wbs_dat_o[26]
port 776 nsew signal output
rlabel metal2 s 116766 0 116822 800 6 wbs_dat_o[27]
port 777 nsew signal output
rlabel metal2 s 120538 0 120594 800 6 wbs_dat_o[28]
port 778 nsew signal output
rlabel metal2 s 124310 0 124366 800 6 wbs_dat_o[29]
port 779 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[2]
port 780 nsew signal output
rlabel metal2 s 128082 0 128138 800 6 wbs_dat_o[30]
port 781 nsew signal output
rlabel metal2 s 131762 0 131818 800 6 wbs_dat_o[31]
port 782 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_o[3]
port 783 nsew signal output
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_o[4]
port 784 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 wbs_dat_o[5]
port 785 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[6]
port 786 nsew signal output
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_o[7]
port 787 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_o[8]
port 788 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 wbs_dat_o[9]
port 789 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_sel_i[0]
port 790 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 wbs_sel_i[1]
port 791 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 wbs_sel_i[2]
port 792 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_sel_i[3]
port 793 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 wbs_stb_i
port 794 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wbs_we_i
port 795 nsew signal input
rlabel metal2 s 145470 119200 145526 120000 6 wmask_o[0]
port 796 nsew signal output
rlabel metal2 s 150346 119200 150402 120000 6 wmask_o[1]
port 797 nsew signal output
rlabel metal3 s 179200 28568 180000 28688 6 wmask_o[2]
port 798 nsew signal output
rlabel metal2 s 139306 0 139362 800 6 wmask_o[3]
port 799 nsew signal output
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 800 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 801 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 802 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 803 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 804 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 805 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 806 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 807 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 808 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 809 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 810 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 811 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 812 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 813 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 814 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 815 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 816 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 817 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 818 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 819 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 820 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 821 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 822 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 823 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 824 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 825 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 826 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 827 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 828 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 829 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 830 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 831 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 832 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 833 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 834 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 835 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 836 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 837 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 838 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 839 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 840 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 841 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 842 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 843 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 844 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 845 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 846 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 847 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 14935224
string GDS_START 972144
<< end >>

