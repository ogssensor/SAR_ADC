magic
tech sky130A
magscale 1 2
timestamp 1625589648
<< obsli1 >>
rect 1104 2159 138828 137649
<< obsm1 >>
rect 474 1844 139458 137680
<< metal2 >>
rect 478 139200 534 140000
rect 1490 139200 1546 140000
rect 2502 139200 2558 140000
rect 3606 139200 3662 140000
rect 4618 139200 4674 140000
rect 5722 139200 5778 140000
rect 6734 139200 6790 140000
rect 7838 139200 7894 140000
rect 8850 139200 8906 140000
rect 9862 139200 9918 140000
rect 10966 139200 11022 140000
rect 11978 139200 12034 140000
rect 13082 139200 13138 140000
rect 14094 139200 14150 140000
rect 15198 139200 15254 140000
rect 16210 139200 16266 140000
rect 17314 139200 17370 140000
rect 18326 139200 18382 140000
rect 19338 139200 19394 140000
rect 20442 139200 20498 140000
rect 21454 139200 21510 140000
rect 22558 139200 22614 140000
rect 23570 139200 23626 140000
rect 24674 139200 24730 140000
rect 25686 139200 25742 140000
rect 26790 139200 26846 140000
rect 27802 139200 27858 140000
rect 28814 139200 28870 140000
rect 29918 139200 29974 140000
rect 30930 139200 30986 140000
rect 32034 139200 32090 140000
rect 33046 139200 33102 140000
rect 34150 139200 34206 140000
rect 35162 139200 35218 140000
rect 36266 139200 36322 140000
rect 37278 139200 37334 140000
rect 38290 139200 38346 140000
rect 39394 139200 39450 140000
rect 40406 139200 40462 140000
rect 41510 139200 41566 140000
rect 42522 139200 42578 140000
rect 43626 139200 43682 140000
rect 44638 139200 44694 140000
rect 45742 139200 45798 140000
rect 46754 139200 46810 140000
rect 47766 139200 47822 140000
rect 48870 139200 48926 140000
rect 49882 139200 49938 140000
rect 50986 139200 51042 140000
rect 51998 139200 52054 140000
rect 53102 139200 53158 140000
rect 54114 139200 54170 140000
rect 55218 139200 55274 140000
rect 56230 139200 56286 140000
rect 57242 139200 57298 140000
rect 58346 139200 58402 140000
rect 59358 139200 59414 140000
rect 60462 139200 60518 140000
rect 61474 139200 61530 140000
rect 62578 139200 62634 140000
rect 63590 139200 63646 140000
rect 64694 139200 64750 140000
rect 65706 139200 65762 140000
rect 66718 139200 66774 140000
rect 67822 139200 67878 140000
rect 68834 139200 68890 140000
rect 69938 139200 69994 140000
rect 70950 139200 71006 140000
rect 72054 139200 72110 140000
rect 73066 139200 73122 140000
rect 74170 139200 74226 140000
rect 75182 139200 75238 140000
rect 76194 139200 76250 140000
rect 77298 139200 77354 140000
rect 78310 139200 78366 140000
rect 79414 139200 79470 140000
rect 80426 139200 80482 140000
rect 81530 139200 81586 140000
rect 82542 139200 82598 140000
rect 83646 139200 83702 140000
rect 84658 139200 84714 140000
rect 85670 139200 85726 140000
rect 86774 139200 86830 140000
rect 87786 139200 87842 140000
rect 88890 139200 88946 140000
rect 89902 139200 89958 140000
rect 91006 139200 91062 140000
rect 92018 139200 92074 140000
rect 93122 139200 93178 140000
rect 94134 139200 94190 140000
rect 95146 139200 95202 140000
rect 96250 139200 96306 140000
rect 97262 139200 97318 140000
rect 98366 139200 98422 140000
rect 99378 139200 99434 140000
rect 100482 139200 100538 140000
rect 101494 139200 101550 140000
rect 102598 139200 102654 140000
rect 103610 139200 103666 140000
rect 104622 139200 104678 140000
rect 105726 139200 105782 140000
rect 106738 139200 106794 140000
rect 107842 139200 107898 140000
rect 108854 139200 108910 140000
rect 109958 139200 110014 140000
rect 110970 139200 111026 140000
rect 112074 139200 112130 140000
rect 113086 139200 113142 140000
rect 114098 139200 114154 140000
rect 115202 139200 115258 140000
rect 116214 139200 116270 140000
rect 117318 139200 117374 140000
rect 118330 139200 118386 140000
rect 119434 139200 119490 140000
rect 120446 139200 120502 140000
rect 121550 139200 121606 140000
rect 122562 139200 122618 140000
rect 123574 139200 123630 140000
rect 124678 139200 124734 140000
rect 125690 139200 125746 140000
rect 126794 139200 126850 140000
rect 127806 139200 127862 140000
rect 128910 139200 128966 140000
rect 129922 139200 129978 140000
rect 131026 139200 131082 140000
rect 132038 139200 132094 140000
rect 133050 139200 133106 140000
rect 134154 139200 134210 140000
rect 135166 139200 135222 140000
rect 136270 139200 136326 140000
rect 137282 139200 137338 140000
rect 138386 139200 138442 140000
rect 139398 139200 139454 140000
rect 662 0 718 800
rect 1950 0 2006 800
rect 3238 0 3294 800
rect 4618 0 4674 800
rect 5906 0 5962 800
rect 7194 0 7250 800
rect 8574 0 8630 800
rect 9862 0 9918 800
rect 11150 0 11206 800
rect 12530 0 12586 800
rect 13818 0 13874 800
rect 15106 0 15162 800
rect 16486 0 16542 800
rect 17774 0 17830 800
rect 19154 0 19210 800
rect 20442 0 20498 800
rect 21730 0 21786 800
rect 23110 0 23166 800
rect 24398 0 24454 800
rect 25686 0 25742 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 31022 0 31078 800
rect 32310 0 32366 800
rect 33598 0 33654 800
rect 34978 0 35034 800
rect 36266 0 36322 800
rect 37646 0 37702 800
rect 38934 0 38990 800
rect 40222 0 40278 800
rect 41602 0 41658 800
rect 42890 0 42946 800
rect 44178 0 44234 800
rect 45558 0 45614 800
rect 46846 0 46902 800
rect 48134 0 48190 800
rect 49514 0 49570 800
rect 50802 0 50858 800
rect 52090 0 52146 800
rect 53470 0 53526 800
rect 54758 0 54814 800
rect 56138 0 56194 800
rect 57426 0 57482 800
rect 58714 0 58770 800
rect 60094 0 60150 800
rect 61382 0 61438 800
rect 62670 0 62726 800
rect 64050 0 64106 800
rect 65338 0 65394 800
rect 66626 0 66682 800
rect 68006 0 68062 800
rect 69294 0 69350 800
rect 70674 0 70730 800
rect 71962 0 72018 800
rect 73250 0 73306 800
rect 74630 0 74686 800
rect 75918 0 75974 800
rect 77206 0 77262 800
rect 78586 0 78642 800
rect 79874 0 79930 800
rect 81162 0 81218 800
rect 82542 0 82598 800
rect 83830 0 83886 800
rect 85118 0 85174 800
rect 86498 0 86554 800
rect 87786 0 87842 800
rect 89166 0 89222 800
rect 90454 0 90510 800
rect 91742 0 91798 800
rect 93122 0 93178 800
rect 94410 0 94466 800
rect 95698 0 95754 800
rect 97078 0 97134 800
rect 98366 0 98422 800
rect 99654 0 99710 800
rect 101034 0 101090 800
rect 102322 0 102378 800
rect 103610 0 103666 800
rect 104990 0 105046 800
rect 106278 0 106334 800
rect 107658 0 107714 800
rect 108946 0 109002 800
rect 110234 0 110290 800
rect 111614 0 111670 800
rect 112902 0 112958 800
rect 114190 0 114246 800
rect 115570 0 115626 800
rect 116858 0 116914 800
rect 118146 0 118202 800
rect 119526 0 119582 800
rect 120814 0 120870 800
rect 122102 0 122158 800
rect 123482 0 123538 800
rect 124770 0 124826 800
rect 126150 0 126206 800
rect 127438 0 127494 800
rect 128726 0 128782 800
rect 130106 0 130162 800
rect 131394 0 131450 800
rect 132682 0 132738 800
rect 134062 0 134118 800
rect 135350 0 135406 800
rect 136638 0 136694 800
rect 138018 0 138074 800
rect 139306 0 139362 800
<< obsm2 >>
rect 590 139144 1434 139641
rect 1602 139144 2446 139641
rect 2614 139144 3550 139641
rect 3718 139144 4562 139641
rect 4730 139144 5666 139641
rect 5834 139144 6678 139641
rect 6846 139144 7782 139641
rect 7950 139144 8794 139641
rect 8962 139144 9806 139641
rect 9974 139144 10910 139641
rect 11078 139144 11922 139641
rect 12090 139144 13026 139641
rect 13194 139144 14038 139641
rect 14206 139144 15142 139641
rect 15310 139144 16154 139641
rect 16322 139144 17258 139641
rect 17426 139144 18270 139641
rect 18438 139144 19282 139641
rect 19450 139144 20386 139641
rect 20554 139144 21398 139641
rect 21566 139144 22502 139641
rect 22670 139144 23514 139641
rect 23682 139144 24618 139641
rect 24786 139144 25630 139641
rect 25798 139144 26734 139641
rect 26902 139144 27746 139641
rect 27914 139144 28758 139641
rect 28926 139144 29862 139641
rect 30030 139144 30874 139641
rect 31042 139144 31978 139641
rect 32146 139144 32990 139641
rect 33158 139144 34094 139641
rect 34262 139144 35106 139641
rect 35274 139144 36210 139641
rect 36378 139144 37222 139641
rect 37390 139144 38234 139641
rect 38402 139144 39338 139641
rect 39506 139144 40350 139641
rect 40518 139144 41454 139641
rect 41622 139144 42466 139641
rect 42634 139144 43570 139641
rect 43738 139144 44582 139641
rect 44750 139144 45686 139641
rect 45854 139144 46698 139641
rect 46866 139144 47710 139641
rect 47878 139144 48814 139641
rect 48982 139144 49826 139641
rect 49994 139144 50930 139641
rect 51098 139144 51942 139641
rect 52110 139144 53046 139641
rect 53214 139144 54058 139641
rect 54226 139144 55162 139641
rect 55330 139144 56174 139641
rect 56342 139144 57186 139641
rect 57354 139144 58290 139641
rect 58458 139144 59302 139641
rect 59470 139144 60406 139641
rect 60574 139144 61418 139641
rect 61586 139144 62522 139641
rect 62690 139144 63534 139641
rect 63702 139144 64638 139641
rect 64806 139144 65650 139641
rect 65818 139144 66662 139641
rect 66830 139144 67766 139641
rect 67934 139144 68778 139641
rect 68946 139144 69882 139641
rect 70050 139144 70894 139641
rect 71062 139144 71998 139641
rect 72166 139144 73010 139641
rect 73178 139144 74114 139641
rect 74282 139144 75126 139641
rect 75294 139144 76138 139641
rect 76306 139144 77242 139641
rect 77410 139144 78254 139641
rect 78422 139144 79358 139641
rect 79526 139144 80370 139641
rect 80538 139144 81474 139641
rect 81642 139144 82486 139641
rect 82654 139144 83590 139641
rect 83758 139144 84602 139641
rect 84770 139144 85614 139641
rect 85782 139144 86718 139641
rect 86886 139144 87730 139641
rect 87898 139144 88834 139641
rect 89002 139144 89846 139641
rect 90014 139144 90950 139641
rect 91118 139144 91962 139641
rect 92130 139144 93066 139641
rect 93234 139144 94078 139641
rect 94246 139144 95090 139641
rect 95258 139144 96194 139641
rect 96362 139144 97206 139641
rect 97374 139144 98310 139641
rect 98478 139144 99322 139641
rect 99490 139144 100426 139641
rect 100594 139144 101438 139641
rect 101606 139144 102542 139641
rect 102710 139144 103554 139641
rect 103722 139144 104566 139641
rect 104734 139144 105670 139641
rect 105838 139144 106682 139641
rect 106850 139144 107786 139641
rect 107954 139144 108798 139641
rect 108966 139144 109902 139641
rect 110070 139144 110914 139641
rect 111082 139144 112018 139641
rect 112186 139144 113030 139641
rect 113198 139144 114042 139641
rect 114210 139144 115146 139641
rect 115314 139144 116158 139641
rect 116326 139144 117262 139641
rect 117430 139144 118274 139641
rect 118442 139144 119378 139641
rect 119546 139144 120390 139641
rect 120558 139144 121494 139641
rect 121662 139144 122506 139641
rect 122674 139144 123518 139641
rect 123686 139144 124622 139641
rect 124790 139144 125634 139641
rect 125802 139144 126738 139641
rect 126906 139144 127750 139641
rect 127918 139144 128854 139641
rect 129022 139144 129866 139641
rect 130034 139144 130970 139641
rect 131138 139144 131982 139641
rect 132150 139144 132994 139641
rect 133162 139144 134098 139641
rect 134266 139144 135110 139641
rect 135278 139144 136214 139641
rect 136382 139144 137226 139641
rect 137394 139144 138330 139641
rect 138498 139144 139342 139641
rect 480 856 139452 139144
rect 480 303 606 856
rect 774 303 1894 856
rect 2062 303 3182 856
rect 3350 303 4562 856
rect 4730 303 5850 856
rect 6018 303 7138 856
rect 7306 303 8518 856
rect 8686 303 9806 856
rect 9974 303 11094 856
rect 11262 303 12474 856
rect 12642 303 13762 856
rect 13930 303 15050 856
rect 15218 303 16430 856
rect 16598 303 17718 856
rect 17886 303 19098 856
rect 19266 303 20386 856
rect 20554 303 21674 856
rect 21842 303 23054 856
rect 23222 303 24342 856
rect 24510 303 25630 856
rect 25798 303 27010 856
rect 27178 303 28298 856
rect 28466 303 29586 856
rect 29754 303 30966 856
rect 31134 303 32254 856
rect 32422 303 33542 856
rect 33710 303 34922 856
rect 35090 303 36210 856
rect 36378 303 37590 856
rect 37758 303 38878 856
rect 39046 303 40166 856
rect 40334 303 41546 856
rect 41714 303 42834 856
rect 43002 303 44122 856
rect 44290 303 45502 856
rect 45670 303 46790 856
rect 46958 303 48078 856
rect 48246 303 49458 856
rect 49626 303 50746 856
rect 50914 303 52034 856
rect 52202 303 53414 856
rect 53582 303 54702 856
rect 54870 303 56082 856
rect 56250 303 57370 856
rect 57538 303 58658 856
rect 58826 303 60038 856
rect 60206 303 61326 856
rect 61494 303 62614 856
rect 62782 303 63994 856
rect 64162 303 65282 856
rect 65450 303 66570 856
rect 66738 303 67950 856
rect 68118 303 69238 856
rect 69406 303 70618 856
rect 70786 303 71906 856
rect 72074 303 73194 856
rect 73362 303 74574 856
rect 74742 303 75862 856
rect 76030 303 77150 856
rect 77318 303 78530 856
rect 78698 303 79818 856
rect 79986 303 81106 856
rect 81274 303 82486 856
rect 82654 303 83774 856
rect 83942 303 85062 856
rect 85230 303 86442 856
rect 86610 303 87730 856
rect 87898 303 89110 856
rect 89278 303 90398 856
rect 90566 303 91686 856
rect 91854 303 93066 856
rect 93234 303 94354 856
rect 94522 303 95642 856
rect 95810 303 97022 856
rect 97190 303 98310 856
rect 98478 303 99598 856
rect 99766 303 100978 856
rect 101146 303 102266 856
rect 102434 303 103554 856
rect 103722 303 104934 856
rect 105102 303 106222 856
rect 106390 303 107602 856
rect 107770 303 108890 856
rect 109058 303 110178 856
rect 110346 303 111558 856
rect 111726 303 112846 856
rect 113014 303 114134 856
rect 114302 303 115514 856
rect 115682 303 116802 856
rect 116970 303 118090 856
rect 118258 303 119470 856
rect 119638 303 120758 856
rect 120926 303 122046 856
rect 122214 303 123426 856
rect 123594 303 124714 856
rect 124882 303 126094 856
rect 126262 303 127382 856
rect 127550 303 128670 856
rect 128838 303 130050 856
rect 130218 303 131338 856
rect 131506 303 132626 856
rect 132794 303 134006 856
rect 134174 303 135294 856
rect 135462 303 136582 856
rect 136750 303 137962 856
rect 138130 303 139250 856
rect 139418 303 139452 856
<< metal3 >>
rect 0 139544 800 139664
rect 0 138864 800 138984
rect 0 138184 800 138304
rect 0 137640 800 137760
rect 139200 137504 140000 137624
rect 0 136960 800 137080
rect 0 136280 800 136400
rect 0 135600 800 135720
rect 0 135056 800 135176
rect 0 134376 800 134496
rect 0 133696 800 133816
rect 0 133152 800 133272
rect 139200 132880 140000 133000
rect 0 132472 800 132592
rect 0 131792 800 131912
rect 0 131112 800 131232
rect 0 130568 800 130688
rect 0 129888 800 130008
rect 0 129208 800 129328
rect 0 128664 800 128784
rect 139200 128256 140000 128376
rect 0 127984 800 128104
rect 0 127304 800 127424
rect 0 126624 800 126744
rect 0 126080 800 126200
rect 0 125400 800 125520
rect 0 124720 800 124840
rect 0 124040 800 124160
rect 0 123496 800 123616
rect 139200 123496 140000 123616
rect 0 122816 800 122936
rect 0 122136 800 122256
rect 0 121592 800 121712
rect 0 120912 800 121032
rect 0 120232 800 120352
rect 0 119552 800 119672
rect 0 119008 800 119128
rect 139200 118872 140000 118992
rect 0 118328 800 118448
rect 0 117648 800 117768
rect 0 117104 800 117224
rect 0 116424 800 116544
rect 0 115744 800 115864
rect 0 115064 800 115184
rect 0 114520 800 114640
rect 139200 114248 140000 114368
rect 0 113840 800 113960
rect 0 113160 800 113280
rect 0 112616 800 112736
rect 0 111936 800 112056
rect 0 111256 800 111376
rect 0 110576 800 110696
rect 0 110032 800 110152
rect 0 109352 800 109472
rect 139200 109488 140000 109608
rect 0 108672 800 108792
rect 0 107992 800 108112
rect 0 107448 800 107568
rect 0 106768 800 106888
rect 0 106088 800 106208
rect 0 105544 800 105664
rect 0 104864 800 104984
rect 139200 104864 140000 104984
rect 0 104184 800 104304
rect 0 103504 800 103624
rect 0 102960 800 103080
rect 0 102280 800 102400
rect 0 101600 800 101720
rect 0 101056 800 101176
rect 0 100376 800 100496
rect 139200 100240 140000 100360
rect 0 99696 800 99816
rect 0 99016 800 99136
rect 0 98472 800 98592
rect 0 97792 800 97912
rect 0 97112 800 97232
rect 0 96568 800 96688
rect 0 95888 800 96008
rect 139200 95616 140000 95736
rect 0 95208 800 95328
rect 0 94528 800 94648
rect 0 93984 800 94104
rect 0 93304 800 93424
rect 0 92624 800 92744
rect 0 91944 800 92064
rect 0 91400 800 91520
rect 0 90720 800 90840
rect 139200 90856 140000 90976
rect 0 90040 800 90160
rect 0 89496 800 89616
rect 0 88816 800 88936
rect 0 88136 800 88256
rect 0 87456 800 87576
rect 0 86912 800 87032
rect 0 86232 800 86352
rect 139200 86232 140000 86352
rect 0 85552 800 85672
rect 0 85008 800 85128
rect 0 84328 800 84448
rect 0 83648 800 83768
rect 0 82968 800 83088
rect 0 82424 800 82544
rect 0 81744 800 81864
rect 139200 81608 140000 81728
rect 0 81064 800 81184
rect 0 80520 800 80640
rect 0 79840 800 79960
rect 0 79160 800 79280
rect 0 78480 800 78600
rect 0 77936 800 78056
rect 0 77256 800 77376
rect 139200 76848 140000 76968
rect 0 76576 800 76696
rect 0 75896 800 76016
rect 0 75352 800 75472
rect 0 74672 800 74792
rect 0 73992 800 74112
rect 0 73448 800 73568
rect 0 72768 800 72888
rect 0 72088 800 72208
rect 139200 72224 140000 72344
rect 0 71408 800 71528
rect 0 70864 800 70984
rect 0 70184 800 70304
rect 0 69504 800 69624
rect 0 68960 800 69080
rect 0 68280 800 68400
rect 0 67600 800 67720
rect 139200 67600 140000 67720
rect 0 66920 800 67040
rect 0 66376 800 66496
rect 0 65696 800 65816
rect 0 65016 800 65136
rect 0 64472 800 64592
rect 0 63792 800 63912
rect 0 63112 800 63232
rect 139200 62840 140000 62960
rect 0 62432 800 62552
rect 0 61888 800 62008
rect 0 61208 800 61328
rect 0 60528 800 60648
rect 0 59848 800 59968
rect 0 59304 800 59424
rect 0 58624 800 58744
rect 139200 58216 140000 58336
rect 0 57944 800 58064
rect 0 57400 800 57520
rect 0 56720 800 56840
rect 0 56040 800 56160
rect 0 55360 800 55480
rect 0 54816 800 54936
rect 0 54136 800 54256
rect 0 53456 800 53576
rect 139200 53592 140000 53712
rect 0 52912 800 53032
rect 0 52232 800 52352
rect 0 51552 800 51672
rect 0 50872 800 50992
rect 0 50328 800 50448
rect 0 49648 800 49768
rect 0 48968 800 49088
rect 139200 48968 140000 49088
rect 0 48424 800 48544
rect 0 47744 800 47864
rect 0 47064 800 47184
rect 0 46384 800 46504
rect 0 45840 800 45960
rect 0 45160 800 45280
rect 0 44480 800 44600
rect 139200 44208 140000 44328
rect 0 43800 800 43920
rect 0 43256 800 43376
rect 0 42576 800 42696
rect 0 41896 800 42016
rect 0 41352 800 41472
rect 0 40672 800 40792
rect 0 39992 800 40112
rect 139200 39584 140000 39704
rect 0 39312 800 39432
rect 0 38768 800 38888
rect 0 38088 800 38208
rect 0 37408 800 37528
rect 0 36864 800 36984
rect 0 36184 800 36304
rect 0 35504 800 35624
rect 0 34824 800 34944
rect 139200 34960 140000 35080
rect 0 34280 800 34400
rect 0 33600 800 33720
rect 0 32920 800 33040
rect 0 32376 800 32496
rect 0 31696 800 31816
rect 0 31016 800 31136
rect 0 30336 800 30456
rect 139200 30200 140000 30320
rect 0 29792 800 29912
rect 0 29112 800 29232
rect 0 28432 800 28552
rect 0 27752 800 27872
rect 0 27208 800 27328
rect 0 26528 800 26648
rect 0 25848 800 25968
rect 139200 25576 140000 25696
rect 0 25304 800 25424
rect 0 24624 800 24744
rect 0 23944 800 24064
rect 0 23264 800 23384
rect 0 22720 800 22840
rect 0 22040 800 22160
rect 0 21360 800 21480
rect 0 20816 800 20936
rect 139200 20952 140000 21072
rect 0 20136 800 20256
rect 0 19456 800 19576
rect 0 18776 800 18896
rect 0 18232 800 18352
rect 0 17552 800 17672
rect 0 16872 800 16992
rect 0 16328 800 16448
rect 139200 16192 140000 16312
rect 0 15648 800 15768
rect 0 14968 800 15088
rect 0 14288 800 14408
rect 0 13744 800 13864
rect 0 13064 800 13184
rect 0 12384 800 12504
rect 0 11704 800 11824
rect 139200 11568 140000 11688
rect 0 11160 800 11280
rect 0 10480 800 10600
rect 0 9800 800 9920
rect 0 9256 800 9376
rect 0 8576 800 8696
rect 0 7896 800 8016
rect 0 7216 800 7336
rect 139200 6944 140000 7064
rect 0 6672 800 6792
rect 0 5992 800 6112
rect 0 5312 800 5432
rect 0 4768 800 4888
rect 0 4088 800 4208
rect 0 3408 800 3528
rect 0 2728 800 2848
rect 0 2184 800 2304
rect 139200 2320 140000 2440
rect 0 1504 800 1624
rect 0 824 800 944
rect 0 280 800 400
<< obsm3 >>
rect 880 139464 139200 139637
rect 800 139064 139200 139464
rect 880 138784 139200 139064
rect 800 138384 139200 138784
rect 880 138104 139200 138384
rect 800 137840 139200 138104
rect 880 137704 139200 137840
rect 880 137560 139120 137704
rect 800 137424 139120 137560
rect 800 137160 139200 137424
rect 880 136880 139200 137160
rect 800 136480 139200 136880
rect 880 136200 139200 136480
rect 800 135800 139200 136200
rect 880 135520 139200 135800
rect 800 135256 139200 135520
rect 880 134976 139200 135256
rect 800 134576 139200 134976
rect 880 134296 139200 134576
rect 800 133896 139200 134296
rect 880 133616 139200 133896
rect 800 133352 139200 133616
rect 880 133080 139200 133352
rect 880 133072 139120 133080
rect 800 132800 139120 133072
rect 800 132672 139200 132800
rect 880 132392 139200 132672
rect 800 131992 139200 132392
rect 880 131712 139200 131992
rect 800 131312 139200 131712
rect 880 131032 139200 131312
rect 800 130768 139200 131032
rect 880 130488 139200 130768
rect 800 130088 139200 130488
rect 880 129808 139200 130088
rect 800 129408 139200 129808
rect 880 129128 139200 129408
rect 800 128864 139200 129128
rect 880 128584 139200 128864
rect 800 128456 139200 128584
rect 800 128184 139120 128456
rect 880 128176 139120 128184
rect 880 127904 139200 128176
rect 800 127504 139200 127904
rect 880 127224 139200 127504
rect 800 126824 139200 127224
rect 880 126544 139200 126824
rect 800 126280 139200 126544
rect 880 126000 139200 126280
rect 800 125600 139200 126000
rect 880 125320 139200 125600
rect 800 124920 139200 125320
rect 880 124640 139200 124920
rect 800 124240 139200 124640
rect 880 123960 139200 124240
rect 800 123696 139200 123960
rect 880 123416 139120 123696
rect 800 123016 139200 123416
rect 880 122736 139200 123016
rect 800 122336 139200 122736
rect 880 122056 139200 122336
rect 800 121792 139200 122056
rect 880 121512 139200 121792
rect 800 121112 139200 121512
rect 880 120832 139200 121112
rect 800 120432 139200 120832
rect 880 120152 139200 120432
rect 800 119752 139200 120152
rect 880 119472 139200 119752
rect 800 119208 139200 119472
rect 880 119072 139200 119208
rect 880 118928 139120 119072
rect 800 118792 139120 118928
rect 800 118528 139200 118792
rect 880 118248 139200 118528
rect 800 117848 139200 118248
rect 880 117568 139200 117848
rect 800 117304 139200 117568
rect 880 117024 139200 117304
rect 800 116624 139200 117024
rect 880 116344 139200 116624
rect 800 115944 139200 116344
rect 880 115664 139200 115944
rect 800 115264 139200 115664
rect 880 114984 139200 115264
rect 800 114720 139200 114984
rect 880 114448 139200 114720
rect 880 114440 139120 114448
rect 800 114168 139120 114440
rect 800 114040 139200 114168
rect 880 113760 139200 114040
rect 800 113360 139200 113760
rect 880 113080 139200 113360
rect 800 112816 139200 113080
rect 880 112536 139200 112816
rect 800 112136 139200 112536
rect 880 111856 139200 112136
rect 800 111456 139200 111856
rect 880 111176 139200 111456
rect 800 110776 139200 111176
rect 880 110496 139200 110776
rect 800 110232 139200 110496
rect 880 109952 139200 110232
rect 800 109688 139200 109952
rect 800 109552 139120 109688
rect 880 109408 139120 109552
rect 880 109272 139200 109408
rect 800 108872 139200 109272
rect 880 108592 139200 108872
rect 800 108192 139200 108592
rect 880 107912 139200 108192
rect 800 107648 139200 107912
rect 880 107368 139200 107648
rect 800 106968 139200 107368
rect 880 106688 139200 106968
rect 800 106288 139200 106688
rect 880 106008 139200 106288
rect 800 105744 139200 106008
rect 880 105464 139200 105744
rect 800 105064 139200 105464
rect 880 104784 139120 105064
rect 800 104384 139200 104784
rect 880 104104 139200 104384
rect 800 103704 139200 104104
rect 880 103424 139200 103704
rect 800 103160 139200 103424
rect 880 102880 139200 103160
rect 800 102480 139200 102880
rect 880 102200 139200 102480
rect 800 101800 139200 102200
rect 880 101520 139200 101800
rect 800 101256 139200 101520
rect 880 100976 139200 101256
rect 800 100576 139200 100976
rect 880 100440 139200 100576
rect 880 100296 139120 100440
rect 800 100160 139120 100296
rect 800 99896 139200 100160
rect 880 99616 139200 99896
rect 800 99216 139200 99616
rect 880 98936 139200 99216
rect 800 98672 139200 98936
rect 880 98392 139200 98672
rect 800 97992 139200 98392
rect 880 97712 139200 97992
rect 800 97312 139200 97712
rect 880 97032 139200 97312
rect 800 96768 139200 97032
rect 880 96488 139200 96768
rect 800 96088 139200 96488
rect 880 95816 139200 96088
rect 880 95808 139120 95816
rect 800 95536 139120 95808
rect 800 95408 139200 95536
rect 880 95128 139200 95408
rect 800 94728 139200 95128
rect 880 94448 139200 94728
rect 800 94184 139200 94448
rect 880 93904 139200 94184
rect 800 93504 139200 93904
rect 880 93224 139200 93504
rect 800 92824 139200 93224
rect 880 92544 139200 92824
rect 800 92144 139200 92544
rect 880 91864 139200 92144
rect 800 91600 139200 91864
rect 880 91320 139200 91600
rect 800 91056 139200 91320
rect 800 90920 139120 91056
rect 880 90776 139120 90920
rect 880 90640 139200 90776
rect 800 90240 139200 90640
rect 880 89960 139200 90240
rect 800 89696 139200 89960
rect 880 89416 139200 89696
rect 800 89016 139200 89416
rect 880 88736 139200 89016
rect 800 88336 139200 88736
rect 880 88056 139200 88336
rect 800 87656 139200 88056
rect 880 87376 139200 87656
rect 800 87112 139200 87376
rect 880 86832 139200 87112
rect 800 86432 139200 86832
rect 880 86152 139120 86432
rect 800 85752 139200 86152
rect 880 85472 139200 85752
rect 800 85208 139200 85472
rect 880 84928 139200 85208
rect 800 84528 139200 84928
rect 880 84248 139200 84528
rect 800 83848 139200 84248
rect 880 83568 139200 83848
rect 800 83168 139200 83568
rect 880 82888 139200 83168
rect 800 82624 139200 82888
rect 880 82344 139200 82624
rect 800 81944 139200 82344
rect 880 81808 139200 81944
rect 880 81664 139120 81808
rect 800 81528 139120 81664
rect 800 81264 139200 81528
rect 880 80984 139200 81264
rect 800 80720 139200 80984
rect 880 80440 139200 80720
rect 800 80040 139200 80440
rect 880 79760 139200 80040
rect 800 79360 139200 79760
rect 880 79080 139200 79360
rect 800 78680 139200 79080
rect 880 78400 139200 78680
rect 800 78136 139200 78400
rect 880 77856 139200 78136
rect 800 77456 139200 77856
rect 880 77176 139200 77456
rect 800 77048 139200 77176
rect 800 76776 139120 77048
rect 880 76768 139120 76776
rect 880 76496 139200 76768
rect 800 76096 139200 76496
rect 880 75816 139200 76096
rect 800 75552 139200 75816
rect 880 75272 139200 75552
rect 800 74872 139200 75272
rect 880 74592 139200 74872
rect 800 74192 139200 74592
rect 880 73912 139200 74192
rect 800 73648 139200 73912
rect 880 73368 139200 73648
rect 800 72968 139200 73368
rect 880 72688 139200 72968
rect 800 72424 139200 72688
rect 800 72288 139120 72424
rect 880 72144 139120 72288
rect 880 72008 139200 72144
rect 800 71608 139200 72008
rect 880 71328 139200 71608
rect 800 71064 139200 71328
rect 880 70784 139200 71064
rect 800 70384 139200 70784
rect 880 70104 139200 70384
rect 800 69704 139200 70104
rect 880 69424 139200 69704
rect 800 69160 139200 69424
rect 880 68880 139200 69160
rect 800 68480 139200 68880
rect 880 68200 139200 68480
rect 800 67800 139200 68200
rect 880 67520 139120 67800
rect 800 67120 139200 67520
rect 880 66840 139200 67120
rect 800 66576 139200 66840
rect 880 66296 139200 66576
rect 800 65896 139200 66296
rect 880 65616 139200 65896
rect 800 65216 139200 65616
rect 880 64936 139200 65216
rect 800 64672 139200 64936
rect 880 64392 139200 64672
rect 800 63992 139200 64392
rect 880 63712 139200 63992
rect 800 63312 139200 63712
rect 880 63040 139200 63312
rect 880 63032 139120 63040
rect 800 62760 139120 63032
rect 800 62632 139200 62760
rect 880 62352 139200 62632
rect 800 62088 139200 62352
rect 880 61808 139200 62088
rect 800 61408 139200 61808
rect 880 61128 139200 61408
rect 800 60728 139200 61128
rect 880 60448 139200 60728
rect 800 60048 139200 60448
rect 880 59768 139200 60048
rect 800 59504 139200 59768
rect 880 59224 139200 59504
rect 800 58824 139200 59224
rect 880 58544 139200 58824
rect 800 58416 139200 58544
rect 800 58144 139120 58416
rect 880 58136 139120 58144
rect 880 57864 139200 58136
rect 800 57600 139200 57864
rect 880 57320 139200 57600
rect 800 56920 139200 57320
rect 880 56640 139200 56920
rect 800 56240 139200 56640
rect 880 55960 139200 56240
rect 800 55560 139200 55960
rect 880 55280 139200 55560
rect 800 55016 139200 55280
rect 880 54736 139200 55016
rect 800 54336 139200 54736
rect 880 54056 139200 54336
rect 800 53792 139200 54056
rect 800 53656 139120 53792
rect 880 53512 139120 53656
rect 880 53376 139200 53512
rect 800 53112 139200 53376
rect 880 52832 139200 53112
rect 800 52432 139200 52832
rect 880 52152 139200 52432
rect 800 51752 139200 52152
rect 880 51472 139200 51752
rect 800 51072 139200 51472
rect 880 50792 139200 51072
rect 800 50528 139200 50792
rect 880 50248 139200 50528
rect 800 49848 139200 50248
rect 880 49568 139200 49848
rect 800 49168 139200 49568
rect 880 48888 139120 49168
rect 800 48624 139200 48888
rect 880 48344 139200 48624
rect 800 47944 139200 48344
rect 880 47664 139200 47944
rect 800 47264 139200 47664
rect 880 46984 139200 47264
rect 800 46584 139200 46984
rect 880 46304 139200 46584
rect 800 46040 139200 46304
rect 880 45760 139200 46040
rect 800 45360 139200 45760
rect 880 45080 139200 45360
rect 800 44680 139200 45080
rect 880 44408 139200 44680
rect 880 44400 139120 44408
rect 800 44128 139120 44400
rect 800 44000 139200 44128
rect 880 43720 139200 44000
rect 800 43456 139200 43720
rect 880 43176 139200 43456
rect 800 42776 139200 43176
rect 880 42496 139200 42776
rect 800 42096 139200 42496
rect 880 41816 139200 42096
rect 800 41552 139200 41816
rect 880 41272 139200 41552
rect 800 40872 139200 41272
rect 880 40592 139200 40872
rect 800 40192 139200 40592
rect 880 39912 139200 40192
rect 800 39784 139200 39912
rect 800 39512 139120 39784
rect 880 39504 139120 39512
rect 880 39232 139200 39504
rect 800 38968 139200 39232
rect 880 38688 139200 38968
rect 800 38288 139200 38688
rect 880 38008 139200 38288
rect 800 37608 139200 38008
rect 880 37328 139200 37608
rect 800 37064 139200 37328
rect 880 36784 139200 37064
rect 800 36384 139200 36784
rect 880 36104 139200 36384
rect 800 35704 139200 36104
rect 880 35424 139200 35704
rect 800 35160 139200 35424
rect 800 35024 139120 35160
rect 880 34880 139120 35024
rect 880 34744 139200 34880
rect 800 34480 139200 34744
rect 880 34200 139200 34480
rect 800 33800 139200 34200
rect 880 33520 139200 33800
rect 800 33120 139200 33520
rect 880 32840 139200 33120
rect 800 32576 139200 32840
rect 880 32296 139200 32576
rect 800 31896 139200 32296
rect 880 31616 139200 31896
rect 800 31216 139200 31616
rect 880 30936 139200 31216
rect 800 30536 139200 30936
rect 880 30400 139200 30536
rect 880 30256 139120 30400
rect 800 30120 139120 30256
rect 800 29992 139200 30120
rect 880 29712 139200 29992
rect 800 29312 139200 29712
rect 880 29032 139200 29312
rect 800 28632 139200 29032
rect 880 28352 139200 28632
rect 800 27952 139200 28352
rect 880 27672 139200 27952
rect 800 27408 139200 27672
rect 880 27128 139200 27408
rect 800 26728 139200 27128
rect 880 26448 139200 26728
rect 800 26048 139200 26448
rect 880 25776 139200 26048
rect 880 25768 139120 25776
rect 800 25504 139120 25768
rect 880 25496 139120 25504
rect 880 25224 139200 25496
rect 800 24824 139200 25224
rect 880 24544 139200 24824
rect 800 24144 139200 24544
rect 880 23864 139200 24144
rect 800 23464 139200 23864
rect 880 23184 139200 23464
rect 800 22920 139200 23184
rect 880 22640 139200 22920
rect 800 22240 139200 22640
rect 880 21960 139200 22240
rect 800 21560 139200 21960
rect 880 21280 139200 21560
rect 800 21152 139200 21280
rect 800 21016 139120 21152
rect 880 20872 139120 21016
rect 880 20736 139200 20872
rect 800 20336 139200 20736
rect 880 20056 139200 20336
rect 800 19656 139200 20056
rect 880 19376 139200 19656
rect 800 18976 139200 19376
rect 880 18696 139200 18976
rect 800 18432 139200 18696
rect 880 18152 139200 18432
rect 800 17752 139200 18152
rect 880 17472 139200 17752
rect 800 17072 139200 17472
rect 880 16792 139200 17072
rect 800 16528 139200 16792
rect 880 16392 139200 16528
rect 880 16248 139120 16392
rect 800 16112 139120 16248
rect 800 15848 139200 16112
rect 880 15568 139200 15848
rect 800 15168 139200 15568
rect 880 14888 139200 15168
rect 800 14488 139200 14888
rect 880 14208 139200 14488
rect 800 13944 139200 14208
rect 880 13664 139200 13944
rect 800 13264 139200 13664
rect 880 12984 139200 13264
rect 800 12584 139200 12984
rect 880 12304 139200 12584
rect 800 11904 139200 12304
rect 880 11768 139200 11904
rect 880 11624 139120 11768
rect 800 11488 139120 11624
rect 800 11360 139200 11488
rect 880 11080 139200 11360
rect 800 10680 139200 11080
rect 880 10400 139200 10680
rect 800 10000 139200 10400
rect 880 9720 139200 10000
rect 800 9456 139200 9720
rect 880 9176 139200 9456
rect 800 8776 139200 9176
rect 880 8496 139200 8776
rect 800 8096 139200 8496
rect 880 7816 139200 8096
rect 800 7416 139200 7816
rect 880 7144 139200 7416
rect 880 7136 139120 7144
rect 800 6872 139120 7136
rect 880 6864 139120 6872
rect 880 6592 139200 6864
rect 800 6192 139200 6592
rect 880 5912 139200 6192
rect 800 5512 139200 5912
rect 880 5232 139200 5512
rect 800 4968 139200 5232
rect 880 4688 139200 4968
rect 800 4288 139200 4688
rect 880 4008 139200 4288
rect 800 3608 139200 4008
rect 880 3328 139200 3608
rect 800 2928 139200 3328
rect 880 2648 139200 2928
rect 800 2520 139200 2648
rect 800 2384 139120 2520
rect 880 2240 139120 2384
rect 880 2104 139200 2240
rect 800 1704 139200 2104
rect 880 1424 139200 1704
rect 800 1024 139200 1424
rect 880 744 139200 1024
rect 800 480 139200 744
rect 880 307 139200 480
<< metal4 >>
rect 4208 2128 4528 137680
rect 19568 2128 19888 137680
rect 34928 2128 35248 137680
rect 50288 2128 50608 137680
rect 65648 2128 65968 137680
rect 81008 2128 81328 137680
rect 96368 2128 96688 137680
rect 111728 2128 112048 137680
rect 127088 2128 127408 137680
<< labels >>
rlabel metal2 s 478 139200 534 140000 6 adc0_dat_i[0]
port 1 nsew signal input
rlabel metal2 s 35162 139200 35218 140000 6 adc0_dat_i[10]
port 2 nsew signal input
rlabel metal2 s 38290 139200 38346 140000 6 adc0_dat_i[11]
port 3 nsew signal input
rlabel metal2 s 41510 139200 41566 140000 6 adc0_dat_i[12]
port 4 nsew signal input
rlabel metal2 s 44638 139200 44694 140000 6 adc0_dat_i[13]
port 5 nsew signal input
rlabel metal2 s 47766 139200 47822 140000 6 adc0_dat_i[14]
port 6 nsew signal input
rlabel metal2 s 50986 139200 51042 140000 6 adc0_dat_i[15]
port 7 nsew signal input
rlabel metal2 s 54114 139200 54170 140000 6 adc0_dat_i[16]
port 8 nsew signal input
rlabel metal2 s 57242 139200 57298 140000 6 adc0_dat_i[17]
port 9 nsew signal input
rlabel metal2 s 60462 139200 60518 140000 6 adc0_dat_i[18]
port 10 nsew signal input
rlabel metal2 s 63590 139200 63646 140000 6 adc0_dat_i[19]
port 11 nsew signal input
rlabel metal2 s 4618 139200 4674 140000 6 adc0_dat_i[1]
port 12 nsew signal input
rlabel metal2 s 66718 139200 66774 140000 6 adc0_dat_i[20]
port 13 nsew signal input
rlabel metal2 s 69938 139200 69994 140000 6 adc0_dat_i[21]
port 14 nsew signal input
rlabel metal2 s 73066 139200 73122 140000 6 adc0_dat_i[22]
port 15 nsew signal input
rlabel metal2 s 76194 139200 76250 140000 6 adc0_dat_i[23]
port 16 nsew signal input
rlabel metal2 s 79414 139200 79470 140000 6 adc0_dat_i[24]
port 17 nsew signal input
rlabel metal2 s 82542 139200 82598 140000 6 adc0_dat_i[25]
port 18 nsew signal input
rlabel metal2 s 85670 139200 85726 140000 6 adc0_dat_i[26]
port 19 nsew signal input
rlabel metal2 s 88890 139200 88946 140000 6 adc0_dat_i[27]
port 20 nsew signal input
rlabel metal2 s 92018 139200 92074 140000 6 adc0_dat_i[28]
port 21 nsew signal input
rlabel metal2 s 95146 139200 95202 140000 6 adc0_dat_i[29]
port 22 nsew signal input
rlabel metal2 s 8850 139200 8906 140000 6 adc0_dat_i[2]
port 23 nsew signal input
rlabel metal2 s 98366 139200 98422 140000 6 adc0_dat_i[30]
port 24 nsew signal input
rlabel metal2 s 101494 139200 101550 140000 6 adc0_dat_i[31]
port 25 nsew signal input
rlabel metal2 s 13082 139200 13138 140000 6 adc0_dat_i[3]
port 26 nsew signal input
rlabel metal2 s 16210 139200 16266 140000 6 adc0_dat_i[4]
port 27 nsew signal input
rlabel metal2 s 19338 139200 19394 140000 6 adc0_dat_i[5]
port 28 nsew signal input
rlabel metal2 s 22558 139200 22614 140000 6 adc0_dat_i[6]
port 29 nsew signal input
rlabel metal2 s 25686 139200 25742 140000 6 adc0_dat_i[7]
port 30 nsew signal input
rlabel metal2 s 28814 139200 28870 140000 6 adc0_dat_i[8]
port 31 nsew signal input
rlabel metal2 s 32034 139200 32090 140000 6 adc0_dat_i[9]
port 32 nsew signal input
rlabel metal2 s 1490 139200 1546 140000 6 adc1_dat_i[0]
port 33 nsew signal input
rlabel metal2 s 36266 139200 36322 140000 6 adc1_dat_i[10]
port 34 nsew signal input
rlabel metal2 s 39394 139200 39450 140000 6 adc1_dat_i[11]
port 35 nsew signal input
rlabel metal2 s 42522 139200 42578 140000 6 adc1_dat_i[12]
port 36 nsew signal input
rlabel metal2 s 45742 139200 45798 140000 6 adc1_dat_i[13]
port 37 nsew signal input
rlabel metal2 s 48870 139200 48926 140000 6 adc1_dat_i[14]
port 38 nsew signal input
rlabel metal2 s 51998 139200 52054 140000 6 adc1_dat_i[15]
port 39 nsew signal input
rlabel metal2 s 55218 139200 55274 140000 6 adc1_dat_i[16]
port 40 nsew signal input
rlabel metal2 s 58346 139200 58402 140000 6 adc1_dat_i[17]
port 41 nsew signal input
rlabel metal2 s 61474 139200 61530 140000 6 adc1_dat_i[18]
port 42 nsew signal input
rlabel metal2 s 64694 139200 64750 140000 6 adc1_dat_i[19]
port 43 nsew signal input
rlabel metal2 s 5722 139200 5778 140000 6 adc1_dat_i[1]
port 44 nsew signal input
rlabel metal2 s 67822 139200 67878 140000 6 adc1_dat_i[20]
port 45 nsew signal input
rlabel metal2 s 70950 139200 71006 140000 6 adc1_dat_i[21]
port 46 nsew signal input
rlabel metal2 s 74170 139200 74226 140000 6 adc1_dat_i[22]
port 47 nsew signal input
rlabel metal2 s 77298 139200 77354 140000 6 adc1_dat_i[23]
port 48 nsew signal input
rlabel metal2 s 80426 139200 80482 140000 6 adc1_dat_i[24]
port 49 nsew signal input
rlabel metal2 s 83646 139200 83702 140000 6 adc1_dat_i[25]
port 50 nsew signal input
rlabel metal2 s 86774 139200 86830 140000 6 adc1_dat_i[26]
port 51 nsew signal input
rlabel metal2 s 89902 139200 89958 140000 6 adc1_dat_i[27]
port 52 nsew signal input
rlabel metal2 s 93122 139200 93178 140000 6 adc1_dat_i[28]
port 53 nsew signal input
rlabel metal2 s 96250 139200 96306 140000 6 adc1_dat_i[29]
port 54 nsew signal input
rlabel metal2 s 9862 139200 9918 140000 6 adc1_dat_i[2]
port 55 nsew signal input
rlabel metal2 s 99378 139200 99434 140000 6 adc1_dat_i[30]
port 56 nsew signal input
rlabel metal2 s 102598 139200 102654 140000 6 adc1_dat_i[31]
port 57 nsew signal input
rlabel metal2 s 14094 139200 14150 140000 6 adc1_dat_i[3]
port 58 nsew signal input
rlabel metal2 s 17314 139200 17370 140000 6 adc1_dat_i[4]
port 59 nsew signal input
rlabel metal2 s 20442 139200 20498 140000 6 adc1_dat_i[5]
port 60 nsew signal input
rlabel metal2 s 23570 139200 23626 140000 6 adc1_dat_i[6]
port 61 nsew signal input
rlabel metal2 s 26790 139200 26846 140000 6 adc1_dat_i[7]
port 62 nsew signal input
rlabel metal2 s 29918 139200 29974 140000 6 adc1_dat_i[8]
port 63 nsew signal input
rlabel metal2 s 33046 139200 33102 140000 6 adc1_dat_i[9]
port 64 nsew signal input
rlabel metal2 s 2502 139200 2558 140000 6 adc2_dat_i[0]
port 65 nsew signal input
rlabel metal2 s 37278 139200 37334 140000 6 adc2_dat_i[10]
port 66 nsew signal input
rlabel metal2 s 40406 139200 40462 140000 6 adc2_dat_i[11]
port 67 nsew signal input
rlabel metal2 s 43626 139200 43682 140000 6 adc2_dat_i[12]
port 68 nsew signal input
rlabel metal2 s 46754 139200 46810 140000 6 adc2_dat_i[13]
port 69 nsew signal input
rlabel metal2 s 49882 139200 49938 140000 6 adc2_dat_i[14]
port 70 nsew signal input
rlabel metal2 s 53102 139200 53158 140000 6 adc2_dat_i[15]
port 71 nsew signal input
rlabel metal2 s 56230 139200 56286 140000 6 adc2_dat_i[16]
port 72 nsew signal input
rlabel metal2 s 59358 139200 59414 140000 6 adc2_dat_i[17]
port 73 nsew signal input
rlabel metal2 s 62578 139200 62634 140000 6 adc2_dat_i[18]
port 74 nsew signal input
rlabel metal2 s 65706 139200 65762 140000 6 adc2_dat_i[19]
port 75 nsew signal input
rlabel metal2 s 6734 139200 6790 140000 6 adc2_dat_i[1]
port 76 nsew signal input
rlabel metal2 s 68834 139200 68890 140000 6 adc2_dat_i[20]
port 77 nsew signal input
rlabel metal2 s 72054 139200 72110 140000 6 adc2_dat_i[21]
port 78 nsew signal input
rlabel metal2 s 75182 139200 75238 140000 6 adc2_dat_i[22]
port 79 nsew signal input
rlabel metal2 s 78310 139200 78366 140000 6 adc2_dat_i[23]
port 80 nsew signal input
rlabel metal2 s 81530 139200 81586 140000 6 adc2_dat_i[24]
port 81 nsew signal input
rlabel metal2 s 84658 139200 84714 140000 6 adc2_dat_i[25]
port 82 nsew signal input
rlabel metal2 s 87786 139200 87842 140000 6 adc2_dat_i[26]
port 83 nsew signal input
rlabel metal2 s 91006 139200 91062 140000 6 adc2_dat_i[27]
port 84 nsew signal input
rlabel metal2 s 94134 139200 94190 140000 6 adc2_dat_i[28]
port 85 nsew signal input
rlabel metal2 s 97262 139200 97318 140000 6 adc2_dat_i[29]
port 86 nsew signal input
rlabel metal2 s 10966 139200 11022 140000 6 adc2_dat_i[2]
port 87 nsew signal input
rlabel metal2 s 100482 139200 100538 140000 6 adc2_dat_i[30]
port 88 nsew signal input
rlabel metal2 s 103610 139200 103666 140000 6 adc2_dat_i[31]
port 89 nsew signal input
rlabel metal2 s 15198 139200 15254 140000 6 adc2_dat_i[3]
port 90 nsew signal input
rlabel metal2 s 18326 139200 18382 140000 6 adc2_dat_i[4]
port 91 nsew signal input
rlabel metal2 s 21454 139200 21510 140000 6 adc2_dat_i[5]
port 92 nsew signal input
rlabel metal2 s 24674 139200 24730 140000 6 adc2_dat_i[6]
port 93 nsew signal input
rlabel metal2 s 27802 139200 27858 140000 6 adc2_dat_i[7]
port 94 nsew signal input
rlabel metal2 s 30930 139200 30986 140000 6 adc2_dat_i[8]
port 95 nsew signal input
rlabel metal2 s 34150 139200 34206 140000 6 adc2_dat_i[9]
port 96 nsew signal input
rlabel metal2 s 3606 139200 3662 140000 6 adc_dvalid_i[0]
port 97 nsew signal input
rlabel metal2 s 7838 139200 7894 140000 6 adc_dvalid_i[1]
port 98 nsew signal input
rlabel metal2 s 11978 139200 12034 140000 6 adc_dvalid_i[2]
port 99 nsew signal input
rlabel metal3 s 139200 6944 140000 7064 6 io_oeb[0]
port 100 nsew signal output
rlabel metal3 s 139200 100240 140000 100360 6 io_oeb[10]
port 101 nsew signal output
rlabel metal3 s 139200 109488 140000 109608 6 io_oeb[11]
port 102 nsew signal output
rlabel metal3 s 139200 118872 140000 118992 6 io_oeb[12]
port 103 nsew signal output
rlabel metal3 s 139200 128256 140000 128376 6 io_oeb[13]
port 104 nsew signal output
rlabel metal3 s 139200 137504 140000 137624 6 io_oeb[14]
port 105 nsew signal output
rlabel metal2 s 139398 139200 139454 140000 6 io_oeb[15]
port 106 nsew signal output
rlabel metal2 s 137282 139200 137338 140000 6 io_oeb[16]
port 107 nsew signal output
rlabel metal2 s 135166 139200 135222 140000 6 io_oeb[17]
port 108 nsew signal output
rlabel metal2 s 133050 139200 133106 140000 6 io_oeb[18]
port 109 nsew signal output
rlabel metal2 s 131026 139200 131082 140000 6 io_oeb[19]
port 110 nsew signal output
rlabel metal3 s 139200 16192 140000 16312 6 io_oeb[1]
port 111 nsew signal output
rlabel metal2 s 128910 139200 128966 140000 6 io_oeb[20]
port 112 nsew signal output
rlabel metal2 s 126794 139200 126850 140000 6 io_oeb[21]
port 113 nsew signal output
rlabel metal2 s 124678 139200 124734 140000 6 io_oeb[22]
port 114 nsew signal output
rlabel metal2 s 122562 139200 122618 140000 6 io_oeb[23]
port 115 nsew signal output
rlabel metal3 s 0 122816 800 122936 6 io_oeb[24]
port 116 nsew signal output
rlabel metal3 s 0 124040 800 124160 6 io_oeb[25]
port 117 nsew signal output
rlabel metal3 s 0 125400 800 125520 6 io_oeb[26]
port 118 nsew signal output
rlabel metal3 s 0 126624 800 126744 6 io_oeb[27]
port 119 nsew signal output
rlabel metal3 s 0 127984 800 128104 6 io_oeb[28]
port 120 nsew signal output
rlabel metal3 s 0 129208 800 129328 6 io_oeb[29]
port 121 nsew signal output
rlabel metal3 s 139200 25576 140000 25696 6 io_oeb[2]
port 122 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 io_oeb[30]
port 123 nsew signal output
rlabel metal3 s 0 131792 800 131912 6 io_oeb[31]
port 124 nsew signal output
rlabel metal3 s 0 133152 800 133272 6 io_oeb[32]
port 125 nsew signal output
rlabel metal3 s 0 134376 800 134496 6 io_oeb[33]
port 126 nsew signal output
rlabel metal3 s 0 135600 800 135720 6 io_oeb[34]
port 127 nsew signal output
rlabel metal3 s 0 136960 800 137080 6 io_oeb[35]
port 128 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 io_oeb[36]
port 129 nsew signal output
rlabel metal3 s 0 139544 800 139664 6 io_oeb[37]
port 130 nsew signal output
rlabel metal3 s 139200 34960 140000 35080 6 io_oeb[3]
port 131 nsew signal output
rlabel metal3 s 139200 44208 140000 44328 6 io_oeb[4]
port 132 nsew signal output
rlabel metal3 s 139200 53592 140000 53712 6 io_oeb[5]
port 133 nsew signal output
rlabel metal3 s 139200 62840 140000 62960 6 io_oeb[6]
port 134 nsew signal output
rlabel metal3 s 139200 72224 140000 72344 6 io_oeb[7]
port 135 nsew signal output
rlabel metal3 s 139200 81608 140000 81728 6 io_oeb[8]
port 136 nsew signal output
rlabel metal3 s 139200 90856 140000 90976 6 io_oeb[9]
port 137 nsew signal output
rlabel metal3 s 139200 2320 140000 2440 6 io_out[0]
port 138 nsew signal output
rlabel metal3 s 139200 95616 140000 95736 6 io_out[10]
port 139 nsew signal output
rlabel metal3 s 139200 104864 140000 104984 6 io_out[11]
port 140 nsew signal output
rlabel metal3 s 139200 114248 140000 114368 6 io_out[12]
port 141 nsew signal output
rlabel metal3 s 139200 123496 140000 123616 6 io_out[13]
port 142 nsew signal output
rlabel metal3 s 139200 132880 140000 133000 6 io_out[14]
port 143 nsew signal output
rlabel metal2 s 138386 139200 138442 140000 6 io_out[15]
port 144 nsew signal output
rlabel metal2 s 136270 139200 136326 140000 6 io_out[16]
port 145 nsew signal output
rlabel metal2 s 134154 139200 134210 140000 6 io_out[17]
port 146 nsew signal output
rlabel metal2 s 132038 139200 132094 140000 6 io_out[18]
port 147 nsew signal output
rlabel metal2 s 129922 139200 129978 140000 6 io_out[19]
port 148 nsew signal output
rlabel metal3 s 139200 11568 140000 11688 6 io_out[1]
port 149 nsew signal output
rlabel metal2 s 127806 139200 127862 140000 6 io_out[20]
port 150 nsew signal output
rlabel metal2 s 125690 139200 125746 140000 6 io_out[21]
port 151 nsew signal output
rlabel metal2 s 123574 139200 123630 140000 6 io_out[22]
port 152 nsew signal output
rlabel metal2 s 121550 139200 121606 140000 6 io_out[23]
port 153 nsew signal output
rlabel metal3 s 0 122136 800 122256 6 io_out[24]
port 154 nsew signal output
rlabel metal3 s 0 123496 800 123616 6 io_out[25]
port 155 nsew signal output
rlabel metal3 s 0 124720 800 124840 6 io_out[26]
port 156 nsew signal output
rlabel metal3 s 0 126080 800 126200 6 io_out[27]
port 157 nsew signal output
rlabel metal3 s 0 127304 800 127424 6 io_out[28]
port 158 nsew signal output
rlabel metal3 s 0 128664 800 128784 6 io_out[29]
port 159 nsew signal output
rlabel metal3 s 139200 20952 140000 21072 6 io_out[2]
port 160 nsew signal output
rlabel metal3 s 0 129888 800 130008 6 io_out[30]
port 161 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 io_out[31]
port 162 nsew signal output
rlabel metal3 s 0 132472 800 132592 6 io_out[32]
port 163 nsew signal output
rlabel metal3 s 0 133696 800 133816 6 io_out[33]
port 164 nsew signal output
rlabel metal3 s 0 135056 800 135176 6 io_out[34]
port 165 nsew signal output
rlabel metal3 s 0 136280 800 136400 6 io_out[35]
port 166 nsew signal output
rlabel metal3 s 0 137640 800 137760 6 io_out[36]
port 167 nsew signal output
rlabel metal3 s 0 138864 800 138984 6 io_out[37]
port 168 nsew signal output
rlabel metal3 s 139200 30200 140000 30320 6 io_out[3]
port 169 nsew signal output
rlabel metal3 s 139200 39584 140000 39704 6 io_out[4]
port 170 nsew signal output
rlabel metal3 s 139200 48968 140000 49088 6 io_out[5]
port 171 nsew signal output
rlabel metal3 s 139200 58216 140000 58336 6 io_out[6]
port 172 nsew signal output
rlabel metal3 s 139200 67600 140000 67720 6 io_out[7]
port 173 nsew signal output
rlabel metal3 s 139200 76848 140000 76968 6 io_out[8]
port 174 nsew signal output
rlabel metal3 s 139200 86232 140000 86352 6 io_out[9]
port 175 nsew signal output
rlabel metal3 s 0 39992 800 40112 6 mem0_data_i[0]
port 176 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 mem0_data_i[10]
port 177 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 mem0_data_i[11]
port 178 nsew signal input
rlabel metal3 s 0 70864 800 70984 6 mem0_data_i[12]
port 179 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 mem0_data_i[13]
port 180 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 mem0_data_i[14]
port 181 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 mem0_data_i[15]
port 182 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 mem0_data_i[16]
port 183 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 mem0_data_i[17]
port 184 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 mem0_data_i[18]
port 185 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 mem0_data_i[19]
port 186 nsew signal input
rlabel metal3 s 0 42576 800 42696 6 mem0_data_i[1]
port 187 nsew signal input
rlabel metal3 s 0 91400 800 91520 6 mem0_data_i[20]
port 188 nsew signal input
rlabel metal3 s 0 93984 800 94104 6 mem0_data_i[21]
port 189 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 mem0_data_i[22]
port 190 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 mem0_data_i[23]
port 191 nsew signal input
rlabel metal3 s 0 101600 800 101720 6 mem0_data_i[24]
port 192 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 mem0_data_i[25]
port 193 nsew signal input
rlabel metal3 s 0 106768 800 106888 6 mem0_data_i[26]
port 194 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 mem0_data_i[27]
port 195 nsew signal input
rlabel metal3 s 0 111936 800 112056 6 mem0_data_i[28]
port 196 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 mem0_data_i[29]
port 197 nsew signal input
rlabel metal3 s 0 45160 800 45280 6 mem0_data_i[2]
port 198 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 mem0_data_i[30]
port 199 nsew signal input
rlabel metal3 s 0 119552 800 119672 6 mem0_data_i[31]
port 200 nsew signal input
rlabel metal3 s 0 47744 800 47864 6 mem0_data_i[3]
port 201 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 mem0_data_i[4]
port 202 nsew signal input
rlabel metal3 s 0 52912 800 53032 6 mem0_data_i[5]
port 203 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 mem0_data_i[6]
port 204 nsew signal input
rlabel metal3 s 0 57944 800 58064 6 mem0_data_i[7]
port 205 nsew signal input
rlabel metal3 s 0 60528 800 60648 6 mem0_data_i[8]
port 206 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 mem0_data_i[9]
port 207 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 mem1_data_i[0]
port 208 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 mem1_data_i[10]
port 209 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 mem1_data_i[11]
port 210 nsew signal input
rlabel metal3 s 0 71408 800 71528 6 mem1_data_i[12]
port 211 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 mem1_data_i[13]
port 212 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 mem1_data_i[14]
port 213 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 mem1_data_i[15]
port 214 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 mem1_data_i[16]
port 215 nsew signal input
rlabel metal3 s 0 84328 800 84448 6 mem1_data_i[17]
port 216 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 mem1_data_i[18]
port 217 nsew signal input
rlabel metal3 s 0 89496 800 89616 6 mem1_data_i[19]
port 218 nsew signal input
rlabel metal3 s 0 43256 800 43376 6 mem1_data_i[1]
port 219 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 mem1_data_i[20]
port 220 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 mem1_data_i[21]
port 221 nsew signal input
rlabel metal3 s 0 97112 800 97232 6 mem1_data_i[22]
port 222 nsew signal input
rlabel metal3 s 0 99696 800 99816 6 mem1_data_i[23]
port 223 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 mem1_data_i[24]
port 224 nsew signal input
rlabel metal3 s 0 104864 800 104984 6 mem1_data_i[25]
port 225 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 mem1_data_i[26]
port 226 nsew signal input
rlabel metal3 s 0 110032 800 110152 6 mem1_data_i[27]
port 227 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 mem1_data_i[28]
port 228 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 mem1_data_i[29]
port 229 nsew signal input
rlabel metal3 s 0 45840 800 45960 6 mem1_data_i[2]
port 230 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 mem1_data_i[30]
port 231 nsew signal input
rlabel metal3 s 0 120232 800 120352 6 mem1_data_i[31]
port 232 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 mem1_data_i[3]
port 233 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 mem1_data_i[4]
port 234 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 mem1_data_i[5]
port 235 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 mem1_data_i[6]
port 236 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 mem1_data_i[7]
port 237 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 mem1_data_i[8]
port 238 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 mem1_data_i[9]
port 239 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 mem2_data_i[0]
port 240 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 mem2_data_i[10]
port 241 nsew signal input
rlabel metal3 s 0 69504 800 69624 6 mem2_data_i[11]
port 242 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 mem2_data_i[12]
port 243 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 mem2_data_i[13]
port 244 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 mem2_data_i[14]
port 245 nsew signal input
rlabel metal3 s 0 79840 800 79960 6 mem2_data_i[15]
port 246 nsew signal input
rlabel metal3 s 0 82424 800 82544 6 mem2_data_i[16]
port 247 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 mem2_data_i[17]
port 248 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 mem2_data_i[18]
port 249 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 mem2_data_i[19]
port 250 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 mem2_data_i[1]
port 251 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 mem2_data_i[20]
port 252 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 mem2_data_i[21]
port 253 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 mem2_data_i[22]
port 254 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 mem2_data_i[23]
port 255 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 mem2_data_i[24]
port 256 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 mem2_data_i[25]
port 257 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 mem2_data_i[26]
port 258 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 mem2_data_i[27]
port 259 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 mem2_data_i[28]
port 260 nsew signal input
rlabel metal3 s 0 115744 800 115864 6 mem2_data_i[29]
port 261 nsew signal input
rlabel metal3 s 0 46384 800 46504 6 mem2_data_i[2]
port 262 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 mem2_data_i[30]
port 263 nsew signal input
rlabel metal3 s 0 120912 800 121032 6 mem2_data_i[31]
port 264 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 mem2_data_i[3]
port 265 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 mem2_data_i[4]
port 266 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 mem2_data_i[5]
port 267 nsew signal input
rlabel metal3 s 0 56720 800 56840 6 mem2_data_i[6]
port 268 nsew signal input
rlabel metal3 s 0 59304 800 59424 6 mem2_data_i[7]
port 269 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 mem2_data_i[8]
port 270 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 mem2_data_i[9]
port 271 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 mem3_data_i[0]
port 272 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 mem3_data_i[10]
port 273 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 mem3_data_i[11]
port 274 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 mem3_data_i[12]
port 275 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 mem3_data_i[13]
port 276 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 mem3_data_i[14]
port 277 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 mem3_data_i[15]
port 278 nsew signal input
rlabel metal3 s 0 82968 800 83088 6 mem3_data_i[16]
port 279 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 mem3_data_i[17]
port 280 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 mem3_data_i[18]
port 281 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 mem3_data_i[19]
port 282 nsew signal input
rlabel metal3 s 0 44480 800 44600 6 mem3_data_i[1]
port 283 nsew signal input
rlabel metal3 s 0 93304 800 93424 6 mem3_data_i[20]
port 284 nsew signal input
rlabel metal3 s 0 95888 800 96008 6 mem3_data_i[21]
port 285 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 mem3_data_i[22]
port 286 nsew signal input
rlabel metal3 s 0 101056 800 101176 6 mem3_data_i[23]
port 287 nsew signal input
rlabel metal3 s 0 103504 800 103624 6 mem3_data_i[24]
port 288 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 mem3_data_i[25]
port 289 nsew signal input
rlabel metal3 s 0 108672 800 108792 6 mem3_data_i[26]
port 290 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 mem3_data_i[27]
port 291 nsew signal input
rlabel metal3 s 0 113840 800 113960 6 mem3_data_i[28]
port 292 nsew signal input
rlabel metal3 s 0 116424 800 116544 6 mem3_data_i[29]
port 293 nsew signal input
rlabel metal3 s 0 47064 800 47184 6 mem3_data_i[2]
port 294 nsew signal input
rlabel metal3 s 0 119008 800 119128 6 mem3_data_i[30]
port 295 nsew signal input
rlabel metal3 s 0 121592 800 121712 6 mem3_data_i[31]
port 296 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 mem3_data_i[3]
port 297 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 mem3_data_i[4]
port 298 nsew signal input
rlabel metal3 s 0 54816 800 54936 6 mem3_data_i[5]
port 299 nsew signal input
rlabel metal3 s 0 57400 800 57520 6 mem3_data_i[6]
port 300 nsew signal input
rlabel metal3 s 0 59848 800 59968 6 mem3_data_i[7]
port 301 nsew signal input
rlabel metal3 s 0 62432 800 62552 6 mem3_data_i[8]
port 302 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 mem3_data_i[9]
port 303 nsew signal input
rlabel metal3 s 0 16872 800 16992 6 mem_data_o[0]
port 304 nsew signal output
rlabel metal3 s 0 23264 800 23384 6 mem_data_o[10]
port 305 nsew signal output
rlabel metal3 s 0 23944 800 24064 6 mem_data_o[11]
port 306 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 mem_data_o[12]
port 307 nsew signal output
rlabel metal3 s 0 25304 800 25424 6 mem_data_o[13]
port 308 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 mem_data_o[14]
port 309 nsew signal output
rlabel metal3 s 0 26528 800 26648 6 mem_data_o[15]
port 310 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 mem_data_o[16]
port 311 nsew signal output
rlabel metal3 s 0 27752 800 27872 6 mem_data_o[17]
port 312 nsew signal output
rlabel metal3 s 0 28432 800 28552 6 mem_data_o[18]
port 313 nsew signal output
rlabel metal3 s 0 29112 800 29232 6 mem_data_o[19]
port 314 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 mem_data_o[1]
port 315 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 mem_data_o[20]
port 316 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 mem_data_o[21]
port 317 nsew signal output
rlabel metal3 s 0 31016 800 31136 6 mem_data_o[22]
port 318 nsew signal output
rlabel metal3 s 0 31696 800 31816 6 mem_data_o[23]
port 319 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 mem_data_o[24]
port 320 nsew signal output
rlabel metal3 s 0 32920 800 33040 6 mem_data_o[25]
port 321 nsew signal output
rlabel metal3 s 0 33600 800 33720 6 mem_data_o[26]
port 322 nsew signal output
rlabel metal3 s 0 34280 800 34400 6 mem_data_o[27]
port 323 nsew signal output
rlabel metal3 s 0 34824 800 34944 6 mem_data_o[28]
port 324 nsew signal output
rlabel metal3 s 0 35504 800 35624 6 mem_data_o[29]
port 325 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 mem_data_o[2]
port 326 nsew signal output
rlabel metal3 s 0 36184 800 36304 6 mem_data_o[30]
port 327 nsew signal output
rlabel metal3 s 0 36864 800 36984 6 mem_data_o[31]
port 328 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 mem_data_o[3]
port 329 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 mem_data_o[4]
port 330 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 mem_data_o[5]
port 331 nsew signal output
rlabel metal3 s 0 20816 800 20936 6 mem_data_o[6]
port 332 nsew signal output
rlabel metal3 s 0 21360 800 21480 6 mem_data_o[7]
port 333 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 mem_data_o[8]
port 334 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 mem_data_o[9]
port 335 nsew signal output
rlabel metal3 s 0 280 800 400 6 mem_raddr_o[0]
port 336 nsew signal output
rlabel metal3 s 0 824 800 944 6 mem_raddr_o[1]
port 337 nsew signal output
rlabel metal3 s 0 1504 800 1624 6 mem_raddr_o[2]
port 338 nsew signal output
rlabel metal3 s 0 2184 800 2304 6 mem_raddr_o[3]
port 339 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 mem_raddr_o[4]
port 340 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 mem_raddr_o[5]
port 341 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 mem_raddr_o[6]
port 342 nsew signal output
rlabel metal3 s 0 4768 800 4888 6 mem_raddr_o[7]
port 343 nsew signal output
rlabel metal3 s 0 5312 800 5432 6 mem_raddr_o[8]
port 344 nsew signal output
rlabel metal3 s 0 11704 800 11824 6 mem_renb_o[0]
port 345 nsew signal output
rlabel metal3 s 0 12384 800 12504 6 mem_renb_o[1]
port 346 nsew signal output
rlabel metal3 s 0 13064 800 13184 6 mem_renb_o[2]
port 347 nsew signal output
rlabel metal3 s 0 13744 800 13864 6 mem_renb_o[3]
port 348 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 mem_waddr_o[0]
port 349 nsew signal output
rlabel metal3 s 0 6672 800 6792 6 mem_waddr_o[1]
port 350 nsew signal output
rlabel metal3 s 0 7216 800 7336 6 mem_waddr_o[2]
port 351 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 mem_waddr_o[3]
port 352 nsew signal output
rlabel metal3 s 0 8576 800 8696 6 mem_waddr_o[4]
port 353 nsew signal output
rlabel metal3 s 0 9256 800 9376 6 mem_waddr_o[5]
port 354 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 mem_waddr_o[6]
port 355 nsew signal output
rlabel metal3 s 0 10480 800 10600 6 mem_waddr_o[7]
port 356 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 mem_waddr_o[8]
port 357 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 mem_wenb_o[0]
port 358 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 mem_wenb_o[1]
port 359 nsew signal output
rlabel metal3 s 0 15648 800 15768 6 mem_wenb_o[2]
port 360 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 mem_wenb_o[3]
port 361 nsew signal output
rlabel metal2 s 104622 139200 104678 140000 6 oversample_o[0]
port 362 nsew signal output
rlabel metal2 s 105726 139200 105782 140000 6 oversample_o[1]
port 363 nsew signal output
rlabel metal2 s 106738 139200 106794 140000 6 oversample_o[2]
port 364 nsew signal output
rlabel metal2 s 107842 139200 107898 140000 6 oversample_o[3]
port 365 nsew signal output
rlabel metal2 s 108854 139200 108910 140000 6 oversample_o[4]
port 366 nsew signal output
rlabel metal2 s 109958 139200 110014 140000 6 oversample_o[5]
port 367 nsew signal output
rlabel metal2 s 110970 139200 111026 140000 6 oversample_o[6]
port 368 nsew signal output
rlabel metal2 s 112074 139200 112130 140000 6 oversample_o[7]
port 369 nsew signal output
rlabel metal2 s 113086 139200 113142 140000 6 oversample_o[8]
port 370 nsew signal output
rlabel metal2 s 114098 139200 114154 140000 6 oversample_o[9]
port 371 nsew signal output
rlabel metal2 s 118330 139200 118386 140000 6 sinc3_en_o[0]
port 372 nsew signal output
rlabel metal2 s 119434 139200 119490 140000 6 sinc3_en_o[1]
port 373 nsew signal output
rlabel metal2 s 120446 139200 120502 140000 6 sinc3_en_o[2]
port 374 nsew signal output
rlabel metal2 s 115202 139200 115258 140000 6 vco_enb_o[0]
port 375 nsew signal output
rlabel metal2 s 116214 139200 116270 140000 6 vco_enb_o[1]
port 376 nsew signal output
rlabel metal2 s 117318 139200 117374 140000 6 vco_enb_o[2]
port 377 nsew signal output
rlabel metal2 s 662 0 718 800 6 wb_clk_i
port 378 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wb_rst_i
port 379 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_ack_o
port 380 nsew signal output
rlabel metal2 s 8574 0 8630 800 6 wbs_adr_i[0]
port 381 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_adr_i[10]
port 382 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 wbs_adr_i[11]
port 383 nsew signal input
rlabel metal2 s 61382 0 61438 800 6 wbs_adr_i[12]
port 384 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_adr_i[13]
port 385 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 wbs_adr_i[14]
port 386 nsew signal input
rlabel metal2 s 73250 0 73306 800 6 wbs_adr_i[15]
port 387 nsew signal input
rlabel metal2 s 77206 0 77262 800 6 wbs_adr_i[16]
port 388 nsew signal input
rlabel metal2 s 81162 0 81218 800 6 wbs_adr_i[17]
port 389 nsew signal input
rlabel metal2 s 85118 0 85174 800 6 wbs_adr_i[18]
port 390 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[19]
port 391 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[1]
port 392 nsew signal input
rlabel metal2 s 93122 0 93178 800 6 wbs_adr_i[20]
port 393 nsew signal input
rlabel metal2 s 97078 0 97134 800 6 wbs_adr_i[21]
port 394 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 wbs_adr_i[22]
port 395 nsew signal input
rlabel metal2 s 104990 0 105046 800 6 wbs_adr_i[23]
port 396 nsew signal input
rlabel metal2 s 108946 0 109002 800 6 wbs_adr_i[24]
port 397 nsew signal input
rlabel metal2 s 112902 0 112958 800 6 wbs_adr_i[25]
port 398 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 wbs_adr_i[26]
port 399 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 wbs_adr_i[27]
port 400 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 wbs_adr_i[28]
port 401 nsew signal input
rlabel metal2 s 128726 0 128782 800 6 wbs_adr_i[29]
port 402 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_adr_i[2]
port 403 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 wbs_adr_i[30]
port 404 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 wbs_adr_i[31]
port 405 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 wbs_adr_i[3]
port 406 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_adr_i[4]
port 407 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 wbs_adr_i[5]
port 408 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wbs_adr_i[6]
port 409 nsew signal input
rlabel metal2 s 41602 0 41658 800 6 wbs_adr_i[7]
port 410 nsew signal input
rlabel metal2 s 45558 0 45614 800 6 wbs_adr_i[8]
port 411 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 wbs_adr_i[9]
port 412 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_cyc_i
port 413 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_i[0]
port 414 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 wbs_dat_i[10]
port 415 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_i[11]
port 416 nsew signal input
rlabel metal2 s 62670 0 62726 800 6 wbs_dat_i[12]
port 417 nsew signal input
rlabel metal2 s 66626 0 66682 800 6 wbs_dat_i[13]
port 418 nsew signal input
rlabel metal2 s 70674 0 70730 800 6 wbs_dat_i[14]
port 419 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 wbs_dat_i[15]
port 420 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 wbs_dat_i[16]
port 421 nsew signal input
rlabel metal2 s 82542 0 82598 800 6 wbs_dat_i[17]
port 422 nsew signal input
rlabel metal2 s 86498 0 86554 800 6 wbs_dat_i[18]
port 423 nsew signal input
rlabel metal2 s 90454 0 90510 800 6 wbs_dat_i[19]
port 424 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 wbs_dat_i[1]
port 425 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 wbs_dat_i[20]
port 426 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 wbs_dat_i[21]
port 427 nsew signal input
rlabel metal2 s 102322 0 102378 800 6 wbs_dat_i[22]
port 428 nsew signal input
rlabel metal2 s 106278 0 106334 800 6 wbs_dat_i[23]
port 429 nsew signal input
rlabel metal2 s 110234 0 110290 800 6 wbs_dat_i[24]
port 430 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 wbs_dat_i[25]
port 431 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 wbs_dat_i[26]
port 432 nsew signal input
rlabel metal2 s 122102 0 122158 800 6 wbs_dat_i[27]
port 433 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 wbs_dat_i[28]
port 434 nsew signal input
rlabel metal2 s 130106 0 130162 800 6 wbs_dat_i[29]
port 435 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[2]
port 436 nsew signal input
rlabel metal2 s 134062 0 134118 800 6 wbs_dat_i[30]
port 437 nsew signal input
rlabel metal2 s 138018 0 138074 800 6 wbs_dat_i[31]
port 438 nsew signal input
rlabel metal2 s 25686 0 25742 800 6 wbs_dat_i[3]
port 439 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wbs_dat_i[4]
port 440 nsew signal input
rlabel metal2 s 34978 0 35034 800 6 wbs_dat_i[5]
port 441 nsew signal input
rlabel metal2 s 38934 0 38990 800 6 wbs_dat_i[6]
port 442 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_dat_i[7]
port 443 nsew signal input
rlabel metal2 s 46846 0 46902 800 6 wbs_dat_i[8]
port 444 nsew signal input
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_i[9]
port 445 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_dat_o[0]
port 446 nsew signal output
rlabel metal2 s 56138 0 56194 800 6 wbs_dat_o[10]
port 447 nsew signal output
rlabel metal2 s 60094 0 60150 800 6 wbs_dat_o[11]
port 448 nsew signal output
rlabel metal2 s 64050 0 64106 800 6 wbs_dat_o[12]
port 449 nsew signal output
rlabel metal2 s 68006 0 68062 800 6 wbs_dat_o[13]
port 450 nsew signal output
rlabel metal2 s 71962 0 72018 800 6 wbs_dat_o[14]
port 451 nsew signal output
rlabel metal2 s 75918 0 75974 800 6 wbs_dat_o[15]
port 452 nsew signal output
rlabel metal2 s 79874 0 79930 800 6 wbs_dat_o[16]
port 453 nsew signal output
rlabel metal2 s 83830 0 83886 800 6 wbs_dat_o[17]
port 454 nsew signal output
rlabel metal2 s 87786 0 87842 800 6 wbs_dat_o[18]
port 455 nsew signal output
rlabel metal2 s 91742 0 91798 800 6 wbs_dat_o[19]
port 456 nsew signal output
rlabel metal2 s 16486 0 16542 800 6 wbs_dat_o[1]
port 457 nsew signal output
rlabel metal2 s 95698 0 95754 800 6 wbs_dat_o[20]
port 458 nsew signal output
rlabel metal2 s 99654 0 99710 800 6 wbs_dat_o[21]
port 459 nsew signal output
rlabel metal2 s 103610 0 103666 800 6 wbs_dat_o[22]
port 460 nsew signal output
rlabel metal2 s 107658 0 107714 800 6 wbs_dat_o[23]
port 461 nsew signal output
rlabel metal2 s 111614 0 111670 800 6 wbs_dat_o[24]
port 462 nsew signal output
rlabel metal2 s 115570 0 115626 800 6 wbs_dat_o[25]
port 463 nsew signal output
rlabel metal2 s 119526 0 119582 800 6 wbs_dat_o[26]
port 464 nsew signal output
rlabel metal2 s 123482 0 123538 800 6 wbs_dat_o[27]
port 465 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 wbs_dat_o[28]
port 466 nsew signal output
rlabel metal2 s 131394 0 131450 800 6 wbs_dat_o[29]
port 467 nsew signal output
rlabel metal2 s 21730 0 21786 800 6 wbs_dat_o[2]
port 468 nsew signal output
rlabel metal2 s 135350 0 135406 800 6 wbs_dat_o[30]
port 469 nsew signal output
rlabel metal2 s 139306 0 139362 800 6 wbs_dat_o[31]
port 470 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[3]
port 471 nsew signal output
rlabel metal2 s 32310 0 32366 800 6 wbs_dat_o[4]
port 472 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 wbs_dat_o[5]
port 473 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 wbs_dat_o[6]
port 474 nsew signal output
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_o[7]
port 475 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 wbs_dat_o[8]
port 476 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 wbs_dat_o[9]
port 477 nsew signal output
rlabel metal2 s 12530 0 12586 800 6 wbs_sel_i[0]
port 478 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_sel_i[1]
port 479 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_sel_i[2]
port 480 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 wbs_sel_i[3]
port 481 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_stb_i
port 482 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_we_i
port 483 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 wmask_o[0]
port 484 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 wmask_o[1]
port 485 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 wmask_o[2]
port 486 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 wmask_o[3]
port 487 nsew signal output
rlabel metal4 s 127088 2128 127408 137680 6 vccd1
port 488 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 137680 6 vccd1
port 489 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 137680 6 vccd1
port 490 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 137680 6 vccd1
port 491 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 137680 6 vccd1
port 492 nsew power bidirectional
rlabel metal4 s 111728 2128 112048 137680 6 vssd1
port 493 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 137680 6 vssd1
port 494 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 137680 6 vssd1
port 495 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 137680 6 vssd1
port 496 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 140000 140000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 9370272
string GDS_START 638592
<< end >>

