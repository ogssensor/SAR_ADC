magic
tech sky130A
magscale 1 2
timestamp 1625379242
<< obsli1 >>
rect 1104 1445 179003 157777
<< obsm1 >>
rect 750 1436 179202 157808
<< metal2 >>
rect 1030 159200 1086 160000
rect 3146 159200 3202 160000
rect 5354 159200 5410 160000
rect 7562 159200 7618 160000
rect 9770 159200 9826 160000
rect 11978 159200 12034 160000
rect 14186 159200 14242 160000
rect 16394 159200 16450 160000
rect 18510 159200 18566 160000
rect 20718 159200 20774 160000
rect 22926 159200 22982 160000
rect 25134 159200 25190 160000
rect 27342 159200 27398 160000
rect 29550 159200 29606 160000
rect 31758 159200 31814 160000
rect 33874 159200 33930 160000
rect 36082 159200 36138 160000
rect 38290 159200 38346 160000
rect 40498 159200 40554 160000
rect 42706 159200 42762 160000
rect 44914 159200 44970 160000
rect 47122 159200 47178 160000
rect 49330 159200 49386 160000
rect 51446 159200 51502 160000
rect 53654 159200 53710 160000
rect 55862 159200 55918 160000
rect 58070 159200 58126 160000
rect 60278 159200 60334 160000
rect 62486 159200 62542 160000
rect 64694 159200 64750 160000
rect 66810 159200 66866 160000
rect 69018 159200 69074 160000
rect 71226 159200 71282 160000
rect 73434 159200 73490 160000
rect 75642 159200 75698 160000
rect 77850 159200 77906 160000
rect 80058 159200 80114 160000
rect 82266 159200 82322 160000
rect 84382 159200 84438 160000
rect 86590 159200 86646 160000
rect 88798 159200 88854 160000
rect 91006 159200 91062 160000
rect 93214 159200 93270 160000
rect 95422 159200 95478 160000
rect 97630 159200 97686 160000
rect 99746 159200 99802 160000
rect 101954 159200 102010 160000
rect 104162 159200 104218 160000
rect 106370 159200 106426 160000
rect 108578 159200 108634 160000
rect 110786 159200 110842 160000
rect 112994 159200 113050 160000
rect 115202 159200 115258 160000
rect 117318 159200 117374 160000
rect 119526 159200 119582 160000
rect 121734 159200 121790 160000
rect 123942 159200 123998 160000
rect 126150 159200 126206 160000
rect 128358 159200 128414 160000
rect 130566 159200 130622 160000
rect 132682 159200 132738 160000
rect 134890 159200 134946 160000
rect 137098 159200 137154 160000
rect 139306 159200 139362 160000
rect 141514 159200 141570 160000
rect 143722 159200 143778 160000
rect 145930 159200 145986 160000
rect 148138 159200 148194 160000
rect 150254 159200 150310 160000
rect 152462 159200 152518 160000
rect 154670 159200 154726 160000
rect 156878 159200 156934 160000
rect 159086 159200 159142 160000
rect 161294 159200 161350 160000
rect 163502 159200 163558 160000
rect 165618 159200 165674 160000
rect 167826 159200 167882 160000
rect 170034 159200 170090 160000
rect 172242 159200 172298 160000
rect 174450 159200 174506 160000
rect 176658 159200 176714 160000
rect 178866 159200 178922 160000
rect 754 0 810 800
rect 2318 0 2374 800
rect 3974 0 4030 800
rect 5630 0 5686 800
rect 7286 0 7342 800
rect 8942 0 8998 800
rect 10598 0 10654 800
rect 12254 0 12310 800
rect 13910 0 13966 800
rect 15566 0 15622 800
rect 17222 0 17278 800
rect 18878 0 18934 800
rect 20534 0 20590 800
rect 22190 0 22246 800
rect 23846 0 23902 800
rect 25502 0 25558 800
rect 27158 0 27214 800
rect 28814 0 28870 800
rect 30470 0 30526 800
rect 32126 0 32182 800
rect 33782 0 33838 800
rect 35438 0 35494 800
rect 37002 0 37058 800
rect 38658 0 38714 800
rect 40314 0 40370 800
rect 41970 0 42026 800
rect 43626 0 43682 800
rect 45282 0 45338 800
rect 46938 0 46994 800
rect 48594 0 48650 800
rect 50250 0 50306 800
rect 51906 0 51962 800
rect 53562 0 53618 800
rect 55218 0 55274 800
rect 56874 0 56930 800
rect 58530 0 58586 800
rect 60186 0 60242 800
rect 61842 0 61898 800
rect 63498 0 63554 800
rect 65154 0 65210 800
rect 66810 0 66866 800
rect 68466 0 68522 800
rect 70122 0 70178 800
rect 71778 0 71834 800
rect 73342 0 73398 800
rect 74998 0 75054 800
rect 76654 0 76710 800
rect 78310 0 78366 800
rect 79966 0 80022 800
rect 81622 0 81678 800
rect 83278 0 83334 800
rect 84934 0 84990 800
rect 86590 0 86646 800
rect 88246 0 88302 800
rect 89902 0 89958 800
rect 91558 0 91614 800
rect 93214 0 93270 800
rect 94870 0 94926 800
rect 96526 0 96582 800
rect 98182 0 98238 800
rect 99838 0 99894 800
rect 101494 0 101550 800
rect 103150 0 103206 800
rect 104806 0 104862 800
rect 106462 0 106518 800
rect 108118 0 108174 800
rect 109682 0 109738 800
rect 111338 0 111394 800
rect 112994 0 113050 800
rect 114650 0 114706 800
rect 116306 0 116362 800
rect 117962 0 118018 800
rect 119618 0 119674 800
rect 121274 0 121330 800
rect 122930 0 122986 800
rect 124586 0 124642 800
rect 126242 0 126298 800
rect 127898 0 127954 800
rect 129554 0 129610 800
rect 131210 0 131266 800
rect 132866 0 132922 800
rect 134522 0 134578 800
rect 136178 0 136234 800
rect 137834 0 137890 800
rect 139490 0 139546 800
rect 141146 0 141202 800
rect 142802 0 142858 800
rect 144458 0 144514 800
rect 146022 0 146078 800
rect 147678 0 147734 800
rect 149334 0 149390 800
rect 150990 0 151046 800
rect 152646 0 152702 800
rect 154302 0 154358 800
rect 155958 0 156014 800
rect 157614 0 157670 800
rect 159270 0 159326 800
rect 160926 0 160982 800
rect 162582 0 162638 800
rect 164238 0 164294 800
rect 165894 0 165950 800
rect 167550 0 167606 800
rect 169206 0 169262 800
rect 170862 0 170918 800
rect 172518 0 172574 800
rect 174174 0 174230 800
rect 175830 0 175886 800
rect 177486 0 177542 800
rect 179142 0 179198 800
<< obsm2 >>
rect 756 159144 974 159225
rect 1142 159144 3090 159225
rect 3258 159144 5298 159225
rect 5466 159144 7506 159225
rect 7674 159144 9714 159225
rect 9882 159144 11922 159225
rect 12090 159144 14130 159225
rect 14298 159144 16338 159225
rect 16506 159144 18454 159225
rect 18622 159144 20662 159225
rect 20830 159144 22870 159225
rect 23038 159144 25078 159225
rect 25246 159144 27286 159225
rect 27454 159144 29494 159225
rect 29662 159144 31702 159225
rect 31870 159144 33818 159225
rect 33986 159144 36026 159225
rect 36194 159144 38234 159225
rect 38402 159144 40442 159225
rect 40610 159144 42650 159225
rect 42818 159144 44858 159225
rect 45026 159144 47066 159225
rect 47234 159144 49274 159225
rect 49442 159144 51390 159225
rect 51558 159144 53598 159225
rect 53766 159144 55806 159225
rect 55974 159144 58014 159225
rect 58182 159144 60222 159225
rect 60390 159144 62430 159225
rect 62598 159144 64638 159225
rect 64806 159144 66754 159225
rect 66922 159144 68962 159225
rect 69130 159144 71170 159225
rect 71338 159144 73378 159225
rect 73546 159144 75586 159225
rect 75754 159144 77794 159225
rect 77962 159144 80002 159225
rect 80170 159144 82210 159225
rect 82378 159144 84326 159225
rect 84494 159144 86534 159225
rect 86702 159144 88742 159225
rect 88910 159144 90950 159225
rect 91118 159144 93158 159225
rect 93326 159144 95366 159225
rect 95534 159144 97574 159225
rect 97742 159144 99690 159225
rect 99858 159144 101898 159225
rect 102066 159144 104106 159225
rect 104274 159144 106314 159225
rect 106482 159144 108522 159225
rect 108690 159144 110730 159225
rect 110898 159144 112938 159225
rect 113106 159144 115146 159225
rect 115314 159144 117262 159225
rect 117430 159144 119470 159225
rect 119638 159144 121678 159225
rect 121846 159144 123886 159225
rect 124054 159144 126094 159225
rect 126262 159144 128302 159225
rect 128470 159144 130510 159225
rect 130678 159144 132626 159225
rect 132794 159144 134834 159225
rect 135002 159144 137042 159225
rect 137210 159144 139250 159225
rect 139418 159144 141458 159225
rect 141626 159144 143666 159225
rect 143834 159144 145874 159225
rect 146042 159144 148082 159225
rect 148250 159144 150198 159225
rect 150366 159144 152406 159225
rect 152574 159144 154614 159225
rect 154782 159144 156822 159225
rect 156990 159144 159030 159225
rect 159198 159144 161238 159225
rect 161406 159144 163446 159225
rect 163614 159144 165562 159225
rect 165730 159144 167770 159225
rect 167938 159144 169978 159225
rect 170146 159144 172186 159225
rect 172354 159144 174394 159225
rect 174562 159144 176602 159225
rect 176770 159144 178810 159225
rect 178978 159144 179196 159225
rect 756 856 179196 159144
rect 866 575 2262 856
rect 2430 575 3918 856
rect 4086 575 5574 856
rect 5742 575 7230 856
rect 7398 575 8886 856
rect 9054 575 10542 856
rect 10710 575 12198 856
rect 12366 575 13854 856
rect 14022 575 15510 856
rect 15678 575 17166 856
rect 17334 575 18822 856
rect 18990 575 20478 856
rect 20646 575 22134 856
rect 22302 575 23790 856
rect 23958 575 25446 856
rect 25614 575 27102 856
rect 27270 575 28758 856
rect 28926 575 30414 856
rect 30582 575 32070 856
rect 32238 575 33726 856
rect 33894 575 35382 856
rect 35550 575 36946 856
rect 37114 575 38602 856
rect 38770 575 40258 856
rect 40426 575 41914 856
rect 42082 575 43570 856
rect 43738 575 45226 856
rect 45394 575 46882 856
rect 47050 575 48538 856
rect 48706 575 50194 856
rect 50362 575 51850 856
rect 52018 575 53506 856
rect 53674 575 55162 856
rect 55330 575 56818 856
rect 56986 575 58474 856
rect 58642 575 60130 856
rect 60298 575 61786 856
rect 61954 575 63442 856
rect 63610 575 65098 856
rect 65266 575 66754 856
rect 66922 575 68410 856
rect 68578 575 70066 856
rect 70234 575 71722 856
rect 71890 575 73286 856
rect 73454 575 74942 856
rect 75110 575 76598 856
rect 76766 575 78254 856
rect 78422 575 79910 856
rect 80078 575 81566 856
rect 81734 575 83222 856
rect 83390 575 84878 856
rect 85046 575 86534 856
rect 86702 575 88190 856
rect 88358 575 89846 856
rect 90014 575 91502 856
rect 91670 575 93158 856
rect 93326 575 94814 856
rect 94982 575 96470 856
rect 96638 575 98126 856
rect 98294 575 99782 856
rect 99950 575 101438 856
rect 101606 575 103094 856
rect 103262 575 104750 856
rect 104918 575 106406 856
rect 106574 575 108062 856
rect 108230 575 109626 856
rect 109794 575 111282 856
rect 111450 575 112938 856
rect 113106 575 114594 856
rect 114762 575 116250 856
rect 116418 575 117906 856
rect 118074 575 119562 856
rect 119730 575 121218 856
rect 121386 575 122874 856
rect 123042 575 124530 856
rect 124698 575 126186 856
rect 126354 575 127842 856
rect 128010 575 129498 856
rect 129666 575 131154 856
rect 131322 575 132810 856
rect 132978 575 134466 856
rect 134634 575 136122 856
rect 136290 575 137778 856
rect 137946 575 139434 856
rect 139602 575 141090 856
rect 141258 575 142746 856
rect 142914 575 144402 856
rect 144570 575 145966 856
rect 146134 575 147622 856
rect 147790 575 149278 856
rect 149446 575 150934 856
rect 151102 575 152590 856
rect 152758 575 154246 856
rect 154414 575 155902 856
rect 156070 575 157558 856
rect 157726 575 159214 856
rect 159382 575 160870 856
rect 161038 575 162526 856
rect 162694 575 164182 856
rect 164350 575 165838 856
rect 166006 575 167494 856
rect 167662 575 169150 856
rect 169318 575 170806 856
rect 170974 575 172462 856
rect 172630 575 174118 856
rect 174286 575 175774 856
rect 175942 575 177430 856
rect 177598 575 179086 856
<< metal3 >>
rect 0 159128 800 159248
rect 179200 159128 180000 159248
rect 0 157768 800 157888
rect 179200 157632 180000 157752
rect 0 156544 800 156664
rect 179200 156136 180000 156256
rect 0 155184 800 155304
rect 179200 154640 180000 154760
rect 0 153824 800 153944
rect 179200 153280 180000 153400
rect 0 152600 800 152720
rect 179200 151784 180000 151904
rect 0 151240 800 151360
rect 179200 150288 180000 150408
rect 0 149880 800 150000
rect 0 148656 800 148776
rect 179200 148792 180000 148912
rect 0 147296 800 147416
rect 179200 147296 180000 147416
rect 0 145936 800 146056
rect 179200 145936 180000 146056
rect 0 144712 800 144832
rect 179200 144440 180000 144560
rect 0 143352 800 143472
rect 179200 142944 180000 143064
rect 0 142128 800 142248
rect 179200 141448 180000 141568
rect 0 140768 800 140888
rect 179200 139952 180000 140072
rect 0 139408 800 139528
rect 179200 138592 180000 138712
rect 0 138184 800 138304
rect 179200 137096 180000 137216
rect 0 136824 800 136944
rect 0 135464 800 135584
rect 179200 135600 180000 135720
rect 0 134240 800 134360
rect 179200 134104 180000 134224
rect 0 132880 800 133000
rect 179200 132744 180000 132864
rect 0 131520 800 131640
rect 179200 131248 180000 131368
rect 0 130296 800 130416
rect 179200 129752 180000 129872
rect 0 128936 800 129056
rect 179200 128256 180000 128376
rect 0 127712 800 127832
rect 179200 126760 180000 126880
rect 0 126352 800 126472
rect 179200 125400 180000 125520
rect 0 124992 800 125112
rect 0 123768 800 123888
rect 179200 123904 180000 124024
rect 0 122408 800 122528
rect 179200 122408 180000 122528
rect 0 121048 800 121168
rect 179200 120912 180000 121032
rect 0 119824 800 119944
rect 179200 119416 180000 119536
rect 0 118464 800 118584
rect 179200 118056 180000 118176
rect 0 117104 800 117224
rect 179200 116560 180000 116680
rect 0 115880 800 116000
rect 179200 115064 180000 115184
rect 0 114520 800 114640
rect 179200 113568 180000 113688
rect 0 113160 800 113280
rect 0 111936 800 112056
rect 179200 112072 180000 112192
rect 0 110576 800 110696
rect 179200 110712 180000 110832
rect 0 109352 800 109472
rect 179200 109216 180000 109336
rect 0 107992 800 108112
rect 179200 107720 180000 107840
rect 0 106632 800 106752
rect 179200 106224 180000 106344
rect 0 105408 800 105528
rect 179200 104864 180000 104984
rect 0 104048 800 104168
rect 179200 103368 180000 103488
rect 0 102688 800 102808
rect 179200 101872 180000 101992
rect 0 101464 800 101584
rect 179200 100376 180000 100496
rect 0 100104 800 100224
rect 0 98744 800 98864
rect 179200 98880 180000 99000
rect 0 97520 800 97640
rect 179200 97520 180000 97640
rect 0 96160 800 96280
rect 179200 96024 180000 96144
rect 0 94936 800 95056
rect 179200 94528 180000 94648
rect 0 93576 800 93696
rect 179200 93032 180000 93152
rect 0 92216 800 92336
rect 179200 91536 180000 91656
rect 0 90992 800 91112
rect 179200 90176 180000 90296
rect 0 89632 800 89752
rect 179200 88680 180000 88800
rect 0 88272 800 88392
rect 0 87048 800 87168
rect 179200 87184 180000 87304
rect 0 85688 800 85808
rect 179200 85688 180000 85808
rect 0 84328 800 84448
rect 179200 84192 180000 84312
rect 0 83104 800 83224
rect 179200 82832 180000 82952
rect 0 81744 800 81864
rect 179200 81336 180000 81456
rect 0 80520 800 80640
rect 179200 79840 180000 79960
rect 0 79160 800 79280
rect 179200 78344 180000 78464
rect 0 77800 800 77920
rect 179200 76984 180000 77104
rect 0 76576 800 76696
rect 179200 75488 180000 75608
rect 0 75216 800 75336
rect 0 73856 800 73976
rect 179200 73992 180000 74112
rect 0 72632 800 72752
rect 179200 72496 180000 72616
rect 0 71272 800 71392
rect 179200 71000 180000 71120
rect 0 69912 800 70032
rect 179200 69640 180000 69760
rect 0 68688 800 68808
rect 179200 68144 180000 68264
rect 0 67328 800 67448
rect 179200 66648 180000 66768
rect 0 65968 800 66088
rect 179200 65152 180000 65272
rect 0 64744 800 64864
rect 179200 63656 180000 63776
rect 0 63384 800 63504
rect 0 62160 800 62280
rect 179200 62296 180000 62416
rect 0 60800 800 60920
rect 179200 60800 180000 60920
rect 0 59440 800 59560
rect 179200 59304 180000 59424
rect 0 58216 800 58336
rect 179200 57808 180000 57928
rect 0 56856 800 56976
rect 179200 56312 180000 56432
rect 0 55496 800 55616
rect 179200 54952 180000 55072
rect 0 54272 800 54392
rect 179200 53456 180000 53576
rect 0 52912 800 53032
rect 179200 51960 180000 52080
rect 0 51552 800 51672
rect 0 50328 800 50448
rect 179200 50464 180000 50584
rect 0 48968 800 49088
rect 179200 49104 180000 49224
rect 0 47744 800 47864
rect 179200 47608 180000 47728
rect 0 46384 800 46504
rect 179200 46112 180000 46232
rect 0 45024 800 45144
rect 179200 44616 180000 44736
rect 0 43800 800 43920
rect 179200 43120 180000 43240
rect 0 42440 800 42560
rect 179200 41760 180000 41880
rect 0 41080 800 41200
rect 179200 40264 180000 40384
rect 0 39856 800 39976
rect 179200 38768 180000 38888
rect 0 38496 800 38616
rect 0 37136 800 37256
rect 179200 37272 180000 37392
rect 0 35912 800 36032
rect 179200 35776 180000 35896
rect 0 34552 800 34672
rect 179200 34416 180000 34536
rect 0 33192 800 33312
rect 179200 32920 180000 33040
rect 0 31968 800 32088
rect 179200 31424 180000 31544
rect 0 30608 800 30728
rect 179200 29928 180000 30048
rect 0 29384 800 29504
rect 179200 28432 180000 28552
rect 0 28024 800 28144
rect 179200 27072 180000 27192
rect 0 26664 800 26784
rect 0 25440 800 25560
rect 179200 25576 180000 25696
rect 0 24080 800 24200
rect 179200 24080 180000 24200
rect 0 22720 800 22840
rect 179200 22584 180000 22704
rect 0 21496 800 21616
rect 179200 21224 180000 21344
rect 0 20136 800 20256
rect 179200 19728 180000 19848
rect 0 18776 800 18896
rect 179200 18232 180000 18352
rect 0 17552 800 17672
rect 179200 16736 180000 16856
rect 0 16192 800 16312
rect 179200 15240 180000 15360
rect 0 14968 800 15088
rect 179200 13880 180000 14000
rect 0 13608 800 13728
rect 0 12248 800 12368
rect 179200 12384 180000 12504
rect 0 11024 800 11144
rect 179200 10888 180000 11008
rect 0 9664 800 9784
rect 179200 9392 180000 9512
rect 0 8304 800 8424
rect 179200 7896 180000 8016
rect 0 7080 800 7200
rect 179200 6536 180000 6656
rect 0 5720 800 5840
rect 179200 5040 180000 5160
rect 0 4360 800 4480
rect 179200 3544 180000 3664
rect 0 3136 800 3256
rect 179200 2048 180000 2168
rect 0 1776 800 1896
rect 0 552 800 672
rect 179200 688 180000 808
<< obsm3 >>
rect 880 159048 179120 159221
rect 800 157968 179200 159048
rect 880 157832 179200 157968
rect 880 157688 179120 157832
rect 800 157552 179120 157688
rect 800 156744 179200 157552
rect 880 156464 179200 156744
rect 800 156336 179200 156464
rect 800 156056 179120 156336
rect 800 155384 179200 156056
rect 880 155104 179200 155384
rect 800 154840 179200 155104
rect 800 154560 179120 154840
rect 800 154024 179200 154560
rect 880 153744 179200 154024
rect 800 153480 179200 153744
rect 800 153200 179120 153480
rect 800 152800 179200 153200
rect 880 152520 179200 152800
rect 800 151984 179200 152520
rect 800 151704 179120 151984
rect 800 151440 179200 151704
rect 880 151160 179200 151440
rect 800 150488 179200 151160
rect 800 150208 179120 150488
rect 800 150080 179200 150208
rect 880 149800 179200 150080
rect 800 148992 179200 149800
rect 800 148856 179120 148992
rect 880 148712 179120 148856
rect 880 148576 179200 148712
rect 800 147496 179200 148576
rect 880 147216 179120 147496
rect 800 146136 179200 147216
rect 880 145856 179120 146136
rect 800 144912 179200 145856
rect 880 144640 179200 144912
rect 880 144632 179120 144640
rect 800 144360 179120 144632
rect 800 143552 179200 144360
rect 880 143272 179200 143552
rect 800 143144 179200 143272
rect 800 142864 179120 143144
rect 800 142328 179200 142864
rect 880 142048 179200 142328
rect 800 141648 179200 142048
rect 800 141368 179120 141648
rect 800 140968 179200 141368
rect 880 140688 179200 140968
rect 800 140152 179200 140688
rect 800 139872 179120 140152
rect 800 139608 179200 139872
rect 880 139328 179200 139608
rect 800 138792 179200 139328
rect 800 138512 179120 138792
rect 800 138384 179200 138512
rect 880 138104 179200 138384
rect 800 137296 179200 138104
rect 800 137024 179120 137296
rect 880 137016 179120 137024
rect 880 136744 179200 137016
rect 800 135800 179200 136744
rect 800 135664 179120 135800
rect 880 135520 179120 135664
rect 880 135384 179200 135520
rect 800 134440 179200 135384
rect 880 134304 179200 134440
rect 880 134160 179120 134304
rect 800 134024 179120 134160
rect 800 133080 179200 134024
rect 880 132944 179200 133080
rect 880 132800 179120 132944
rect 800 132664 179120 132800
rect 800 131720 179200 132664
rect 880 131448 179200 131720
rect 880 131440 179120 131448
rect 800 131168 179120 131440
rect 800 130496 179200 131168
rect 880 130216 179200 130496
rect 800 129952 179200 130216
rect 800 129672 179120 129952
rect 800 129136 179200 129672
rect 880 128856 179200 129136
rect 800 128456 179200 128856
rect 800 128176 179120 128456
rect 800 127912 179200 128176
rect 880 127632 179200 127912
rect 800 126960 179200 127632
rect 800 126680 179120 126960
rect 800 126552 179200 126680
rect 880 126272 179200 126552
rect 800 125600 179200 126272
rect 800 125320 179120 125600
rect 800 125192 179200 125320
rect 880 124912 179200 125192
rect 800 124104 179200 124912
rect 800 123968 179120 124104
rect 880 123824 179120 123968
rect 880 123688 179200 123824
rect 800 122608 179200 123688
rect 880 122328 179120 122608
rect 800 121248 179200 122328
rect 880 121112 179200 121248
rect 880 120968 179120 121112
rect 800 120832 179120 120968
rect 800 120024 179200 120832
rect 880 119744 179200 120024
rect 800 119616 179200 119744
rect 800 119336 179120 119616
rect 800 118664 179200 119336
rect 880 118384 179200 118664
rect 800 118256 179200 118384
rect 800 117976 179120 118256
rect 800 117304 179200 117976
rect 880 117024 179200 117304
rect 800 116760 179200 117024
rect 800 116480 179120 116760
rect 800 116080 179200 116480
rect 880 115800 179200 116080
rect 800 115264 179200 115800
rect 800 114984 179120 115264
rect 800 114720 179200 114984
rect 880 114440 179200 114720
rect 800 113768 179200 114440
rect 800 113488 179120 113768
rect 800 113360 179200 113488
rect 880 113080 179200 113360
rect 800 112272 179200 113080
rect 800 112136 179120 112272
rect 880 111992 179120 112136
rect 880 111856 179200 111992
rect 800 110912 179200 111856
rect 800 110776 179120 110912
rect 880 110632 179120 110776
rect 880 110496 179200 110632
rect 800 109552 179200 110496
rect 880 109416 179200 109552
rect 880 109272 179120 109416
rect 800 109136 179120 109272
rect 800 108192 179200 109136
rect 880 107920 179200 108192
rect 880 107912 179120 107920
rect 800 107640 179120 107912
rect 800 106832 179200 107640
rect 880 106552 179200 106832
rect 800 106424 179200 106552
rect 800 106144 179120 106424
rect 800 105608 179200 106144
rect 880 105328 179200 105608
rect 800 105064 179200 105328
rect 800 104784 179120 105064
rect 800 104248 179200 104784
rect 880 103968 179200 104248
rect 800 103568 179200 103968
rect 800 103288 179120 103568
rect 800 102888 179200 103288
rect 880 102608 179200 102888
rect 800 102072 179200 102608
rect 800 101792 179120 102072
rect 800 101664 179200 101792
rect 880 101384 179200 101664
rect 800 100576 179200 101384
rect 800 100304 179120 100576
rect 880 100296 179120 100304
rect 880 100024 179200 100296
rect 800 99080 179200 100024
rect 800 98944 179120 99080
rect 880 98800 179120 98944
rect 880 98664 179200 98800
rect 800 97720 179200 98664
rect 880 97440 179120 97720
rect 800 96360 179200 97440
rect 880 96224 179200 96360
rect 880 96080 179120 96224
rect 800 95944 179120 96080
rect 800 95136 179200 95944
rect 880 94856 179200 95136
rect 800 94728 179200 94856
rect 800 94448 179120 94728
rect 800 93776 179200 94448
rect 880 93496 179200 93776
rect 800 93232 179200 93496
rect 800 92952 179120 93232
rect 800 92416 179200 92952
rect 880 92136 179200 92416
rect 800 91736 179200 92136
rect 800 91456 179120 91736
rect 800 91192 179200 91456
rect 880 90912 179200 91192
rect 800 90376 179200 90912
rect 800 90096 179120 90376
rect 800 89832 179200 90096
rect 880 89552 179200 89832
rect 800 88880 179200 89552
rect 800 88600 179120 88880
rect 800 88472 179200 88600
rect 880 88192 179200 88472
rect 800 87384 179200 88192
rect 800 87248 179120 87384
rect 880 87104 179120 87248
rect 880 86968 179200 87104
rect 800 85888 179200 86968
rect 880 85608 179120 85888
rect 800 84528 179200 85608
rect 880 84392 179200 84528
rect 880 84248 179120 84392
rect 800 84112 179120 84248
rect 800 83304 179200 84112
rect 880 83032 179200 83304
rect 880 83024 179120 83032
rect 800 82752 179120 83024
rect 800 81944 179200 82752
rect 880 81664 179200 81944
rect 800 81536 179200 81664
rect 800 81256 179120 81536
rect 800 80720 179200 81256
rect 880 80440 179200 80720
rect 800 80040 179200 80440
rect 800 79760 179120 80040
rect 800 79360 179200 79760
rect 880 79080 179200 79360
rect 800 78544 179200 79080
rect 800 78264 179120 78544
rect 800 78000 179200 78264
rect 880 77720 179200 78000
rect 800 77184 179200 77720
rect 800 76904 179120 77184
rect 800 76776 179200 76904
rect 880 76496 179200 76776
rect 800 75688 179200 76496
rect 800 75416 179120 75688
rect 880 75408 179120 75416
rect 880 75136 179200 75408
rect 800 74192 179200 75136
rect 800 74056 179120 74192
rect 880 73912 179120 74056
rect 880 73776 179200 73912
rect 800 72832 179200 73776
rect 880 72696 179200 72832
rect 880 72552 179120 72696
rect 800 72416 179120 72552
rect 800 71472 179200 72416
rect 880 71200 179200 71472
rect 880 71192 179120 71200
rect 800 70920 179120 71192
rect 800 70112 179200 70920
rect 880 69840 179200 70112
rect 880 69832 179120 69840
rect 800 69560 179120 69832
rect 800 68888 179200 69560
rect 880 68608 179200 68888
rect 800 68344 179200 68608
rect 800 68064 179120 68344
rect 800 67528 179200 68064
rect 880 67248 179200 67528
rect 800 66848 179200 67248
rect 800 66568 179120 66848
rect 800 66168 179200 66568
rect 880 65888 179200 66168
rect 800 65352 179200 65888
rect 800 65072 179120 65352
rect 800 64944 179200 65072
rect 880 64664 179200 64944
rect 800 63856 179200 64664
rect 800 63584 179120 63856
rect 880 63576 179120 63584
rect 880 63304 179200 63576
rect 800 62496 179200 63304
rect 800 62360 179120 62496
rect 880 62216 179120 62360
rect 880 62080 179200 62216
rect 800 61000 179200 62080
rect 880 60720 179120 61000
rect 800 59640 179200 60720
rect 880 59504 179200 59640
rect 880 59360 179120 59504
rect 800 59224 179120 59360
rect 800 58416 179200 59224
rect 880 58136 179200 58416
rect 800 58008 179200 58136
rect 800 57728 179120 58008
rect 800 57056 179200 57728
rect 880 56776 179200 57056
rect 800 56512 179200 56776
rect 800 56232 179120 56512
rect 800 55696 179200 56232
rect 880 55416 179200 55696
rect 800 55152 179200 55416
rect 800 54872 179120 55152
rect 800 54472 179200 54872
rect 880 54192 179200 54472
rect 800 53656 179200 54192
rect 800 53376 179120 53656
rect 800 53112 179200 53376
rect 880 52832 179200 53112
rect 800 52160 179200 52832
rect 800 51880 179120 52160
rect 800 51752 179200 51880
rect 880 51472 179200 51752
rect 800 50664 179200 51472
rect 800 50528 179120 50664
rect 880 50384 179120 50528
rect 880 50248 179200 50384
rect 800 49304 179200 50248
rect 800 49168 179120 49304
rect 880 49024 179120 49168
rect 880 48888 179200 49024
rect 800 47944 179200 48888
rect 880 47808 179200 47944
rect 880 47664 179120 47808
rect 800 47528 179120 47664
rect 800 46584 179200 47528
rect 880 46312 179200 46584
rect 880 46304 179120 46312
rect 800 46032 179120 46304
rect 800 45224 179200 46032
rect 880 44944 179200 45224
rect 800 44816 179200 44944
rect 800 44536 179120 44816
rect 800 44000 179200 44536
rect 880 43720 179200 44000
rect 800 43320 179200 43720
rect 800 43040 179120 43320
rect 800 42640 179200 43040
rect 880 42360 179200 42640
rect 800 41960 179200 42360
rect 800 41680 179120 41960
rect 800 41280 179200 41680
rect 880 41000 179200 41280
rect 800 40464 179200 41000
rect 800 40184 179120 40464
rect 800 40056 179200 40184
rect 880 39776 179200 40056
rect 800 38968 179200 39776
rect 800 38696 179120 38968
rect 880 38688 179120 38696
rect 880 38416 179200 38688
rect 800 37472 179200 38416
rect 800 37336 179120 37472
rect 880 37192 179120 37336
rect 880 37056 179200 37192
rect 800 36112 179200 37056
rect 880 35976 179200 36112
rect 880 35832 179120 35976
rect 800 35696 179120 35832
rect 800 34752 179200 35696
rect 880 34616 179200 34752
rect 880 34472 179120 34616
rect 800 34336 179120 34472
rect 800 33392 179200 34336
rect 880 33120 179200 33392
rect 880 33112 179120 33120
rect 800 32840 179120 33112
rect 800 32168 179200 32840
rect 880 31888 179200 32168
rect 800 31624 179200 31888
rect 800 31344 179120 31624
rect 800 30808 179200 31344
rect 880 30528 179200 30808
rect 800 30128 179200 30528
rect 800 29848 179120 30128
rect 800 29584 179200 29848
rect 880 29304 179200 29584
rect 800 28632 179200 29304
rect 800 28352 179120 28632
rect 800 28224 179200 28352
rect 880 27944 179200 28224
rect 800 27272 179200 27944
rect 800 26992 179120 27272
rect 800 26864 179200 26992
rect 880 26584 179200 26864
rect 800 25776 179200 26584
rect 800 25640 179120 25776
rect 880 25496 179120 25640
rect 880 25360 179200 25496
rect 800 24280 179200 25360
rect 880 24000 179120 24280
rect 800 22920 179200 24000
rect 880 22784 179200 22920
rect 880 22640 179120 22784
rect 800 22504 179120 22640
rect 800 21696 179200 22504
rect 880 21424 179200 21696
rect 880 21416 179120 21424
rect 800 21144 179120 21416
rect 800 20336 179200 21144
rect 880 20056 179200 20336
rect 800 19928 179200 20056
rect 800 19648 179120 19928
rect 800 18976 179200 19648
rect 880 18696 179200 18976
rect 800 18432 179200 18696
rect 800 18152 179120 18432
rect 800 17752 179200 18152
rect 880 17472 179200 17752
rect 800 16936 179200 17472
rect 800 16656 179120 16936
rect 800 16392 179200 16656
rect 880 16112 179200 16392
rect 800 15440 179200 16112
rect 800 15168 179120 15440
rect 880 15160 179120 15168
rect 880 14888 179200 15160
rect 800 14080 179200 14888
rect 800 13808 179120 14080
rect 880 13800 179120 13808
rect 880 13528 179200 13800
rect 800 12584 179200 13528
rect 800 12448 179120 12584
rect 880 12304 179120 12448
rect 880 12168 179200 12304
rect 800 11224 179200 12168
rect 880 11088 179200 11224
rect 880 10944 179120 11088
rect 800 10808 179120 10944
rect 800 9864 179200 10808
rect 880 9592 179200 9864
rect 880 9584 179120 9592
rect 800 9312 179120 9584
rect 800 8504 179200 9312
rect 880 8224 179200 8504
rect 800 8096 179200 8224
rect 800 7816 179120 8096
rect 800 7280 179200 7816
rect 880 7000 179200 7280
rect 800 6736 179200 7000
rect 800 6456 179120 6736
rect 800 5920 179200 6456
rect 880 5640 179200 5920
rect 800 5240 179200 5640
rect 800 4960 179120 5240
rect 800 4560 179200 4960
rect 880 4280 179200 4560
rect 800 3744 179200 4280
rect 800 3464 179120 3744
rect 800 3336 179200 3464
rect 880 3056 179200 3336
rect 800 2248 179200 3056
rect 800 1976 179120 2248
rect 880 1968 179120 1976
rect 880 1696 179200 1968
rect 800 888 179200 1696
rect 800 752 179120 888
rect 880 608 179120 752
rect 880 579 179200 608
<< metal4 >>
rect 4208 2128 4528 157808
rect 4868 2176 5188 157760
rect 5528 2176 5848 157760
rect 6188 2176 6508 157760
rect 19568 2128 19888 157808
rect 20228 2176 20548 157760
rect 20888 2176 21208 157760
rect 21548 2176 21868 157760
rect 34928 2128 35248 157808
rect 35588 2176 35908 157760
rect 36248 2176 36568 157760
rect 36908 2176 37228 157760
rect 50288 2128 50608 157808
rect 50948 2176 51268 157760
rect 51608 2176 51928 157760
rect 52268 2176 52588 157760
rect 65648 2128 65968 157808
rect 66308 2176 66628 157760
rect 66968 2176 67288 157760
rect 67628 2176 67948 157760
rect 81008 2128 81328 157808
rect 81668 2176 81988 157760
rect 82328 2176 82648 157760
rect 82988 2176 83308 157760
rect 96368 2128 96688 157808
rect 97028 2176 97348 157760
rect 97688 2176 98008 157760
rect 98348 2176 98668 157760
rect 111728 2128 112048 157808
rect 112388 2176 112708 157760
rect 113048 2176 113368 157760
rect 113708 2176 114028 157760
rect 127088 2128 127408 157808
rect 127748 2176 128068 157760
rect 128408 2176 128728 157760
rect 129068 2176 129388 157760
rect 142448 2128 142768 157808
rect 143108 2176 143428 157760
rect 143768 2176 144088 157760
rect 144428 2176 144748 157760
rect 157808 2128 158128 157808
rect 158468 2176 158788 157760
rect 159128 2176 159448 157760
rect 159788 2176 160108 157760
rect 173168 2128 173488 157808
rect 173828 2176 174148 157760
rect 174488 2176 174808 157760
rect 175148 2176 175468 157760
<< obsm4 >>
rect 177435 6155 177869 151877
<< labels >>
rlabel metal3 s 179200 688 180000 808 6 adc0_dat_i[0]
port 1 nsew signal input
rlabel metal3 s 179200 49104 180000 49224 6 adc0_dat_i[10]
port 2 nsew signal input
rlabel metal3 s 179200 53456 180000 53576 6 adc0_dat_i[11]
port 3 nsew signal input
rlabel metal3 s 179200 57808 180000 57928 6 adc0_dat_i[12]
port 4 nsew signal input
rlabel metal3 s 179200 62296 180000 62416 6 adc0_dat_i[13]
port 5 nsew signal input
rlabel metal3 s 179200 66648 180000 66768 6 adc0_dat_i[14]
port 6 nsew signal input
rlabel metal3 s 179200 71000 180000 71120 6 adc0_dat_i[15]
port 7 nsew signal input
rlabel metal3 s 179200 75488 180000 75608 6 adc0_dat_i[16]
port 8 nsew signal input
rlabel metal3 s 179200 79840 180000 79960 6 adc0_dat_i[17]
port 9 nsew signal input
rlabel metal3 s 179200 84192 180000 84312 6 adc0_dat_i[18]
port 10 nsew signal input
rlabel metal3 s 179200 88680 180000 88800 6 adc0_dat_i[19]
port 11 nsew signal input
rlabel metal3 s 179200 6536 180000 6656 6 adc0_dat_i[1]
port 12 nsew signal input
rlabel metal3 s 179200 93032 180000 93152 6 adc0_dat_i[20]
port 13 nsew signal input
rlabel metal3 s 179200 97520 180000 97640 6 adc0_dat_i[21]
port 14 nsew signal input
rlabel metal3 s 179200 101872 180000 101992 6 adc0_dat_i[22]
port 15 nsew signal input
rlabel metal3 s 179200 106224 180000 106344 6 adc0_dat_i[23]
port 16 nsew signal input
rlabel metal3 s 179200 110712 180000 110832 6 adc0_dat_i[24]
port 17 nsew signal input
rlabel metal3 s 179200 115064 180000 115184 6 adc0_dat_i[25]
port 18 nsew signal input
rlabel metal3 s 179200 119416 180000 119536 6 adc0_dat_i[26]
port 19 nsew signal input
rlabel metal3 s 179200 123904 180000 124024 6 adc0_dat_i[27]
port 20 nsew signal input
rlabel metal3 s 179200 128256 180000 128376 6 adc0_dat_i[28]
port 21 nsew signal input
rlabel metal3 s 179200 132744 180000 132864 6 adc0_dat_i[29]
port 22 nsew signal input
rlabel metal3 s 179200 12384 180000 12504 6 adc0_dat_i[2]
port 23 nsew signal input
rlabel metal3 s 179200 137096 180000 137216 6 adc0_dat_i[30]
port 24 nsew signal input
rlabel metal3 s 179200 141448 180000 141568 6 adc0_dat_i[31]
port 25 nsew signal input
rlabel metal3 s 179200 18232 180000 18352 6 adc0_dat_i[3]
port 26 nsew signal input
rlabel metal3 s 179200 22584 180000 22704 6 adc0_dat_i[4]
port 27 nsew signal input
rlabel metal3 s 179200 27072 180000 27192 6 adc0_dat_i[5]
port 28 nsew signal input
rlabel metal3 s 179200 31424 180000 31544 6 adc0_dat_i[6]
port 29 nsew signal input
rlabel metal3 s 179200 35776 180000 35896 6 adc0_dat_i[7]
port 30 nsew signal input
rlabel metal3 s 179200 40264 180000 40384 6 adc0_dat_i[8]
port 31 nsew signal input
rlabel metal3 s 179200 44616 180000 44736 6 adc0_dat_i[9]
port 32 nsew signal input
rlabel metal3 s 179200 2048 180000 2168 6 adc1_dat_i[0]
port 33 nsew signal input
rlabel metal3 s 179200 50464 180000 50584 6 adc1_dat_i[10]
port 34 nsew signal input
rlabel metal3 s 179200 54952 180000 55072 6 adc1_dat_i[11]
port 35 nsew signal input
rlabel metal3 s 179200 59304 180000 59424 6 adc1_dat_i[12]
port 36 nsew signal input
rlabel metal3 s 179200 63656 180000 63776 6 adc1_dat_i[13]
port 37 nsew signal input
rlabel metal3 s 179200 68144 180000 68264 6 adc1_dat_i[14]
port 38 nsew signal input
rlabel metal3 s 179200 72496 180000 72616 6 adc1_dat_i[15]
port 39 nsew signal input
rlabel metal3 s 179200 76984 180000 77104 6 adc1_dat_i[16]
port 40 nsew signal input
rlabel metal3 s 179200 81336 180000 81456 6 adc1_dat_i[17]
port 41 nsew signal input
rlabel metal3 s 179200 85688 180000 85808 6 adc1_dat_i[18]
port 42 nsew signal input
rlabel metal3 s 179200 90176 180000 90296 6 adc1_dat_i[19]
port 43 nsew signal input
rlabel metal3 s 179200 7896 180000 8016 6 adc1_dat_i[1]
port 44 nsew signal input
rlabel metal3 s 179200 94528 180000 94648 6 adc1_dat_i[20]
port 45 nsew signal input
rlabel metal3 s 179200 98880 180000 99000 6 adc1_dat_i[21]
port 46 nsew signal input
rlabel metal3 s 179200 103368 180000 103488 6 adc1_dat_i[22]
port 47 nsew signal input
rlabel metal3 s 179200 107720 180000 107840 6 adc1_dat_i[23]
port 48 nsew signal input
rlabel metal3 s 179200 112072 180000 112192 6 adc1_dat_i[24]
port 49 nsew signal input
rlabel metal3 s 179200 116560 180000 116680 6 adc1_dat_i[25]
port 50 nsew signal input
rlabel metal3 s 179200 120912 180000 121032 6 adc1_dat_i[26]
port 51 nsew signal input
rlabel metal3 s 179200 125400 180000 125520 6 adc1_dat_i[27]
port 52 nsew signal input
rlabel metal3 s 179200 129752 180000 129872 6 adc1_dat_i[28]
port 53 nsew signal input
rlabel metal3 s 179200 134104 180000 134224 6 adc1_dat_i[29]
port 54 nsew signal input
rlabel metal3 s 179200 13880 180000 14000 6 adc1_dat_i[2]
port 55 nsew signal input
rlabel metal3 s 179200 138592 180000 138712 6 adc1_dat_i[30]
port 56 nsew signal input
rlabel metal3 s 179200 142944 180000 143064 6 adc1_dat_i[31]
port 57 nsew signal input
rlabel metal3 s 179200 19728 180000 19848 6 adc1_dat_i[3]
port 58 nsew signal input
rlabel metal3 s 179200 24080 180000 24200 6 adc1_dat_i[4]
port 59 nsew signal input
rlabel metal3 s 179200 28432 180000 28552 6 adc1_dat_i[5]
port 60 nsew signal input
rlabel metal3 s 179200 32920 180000 33040 6 adc1_dat_i[6]
port 61 nsew signal input
rlabel metal3 s 179200 37272 180000 37392 6 adc1_dat_i[7]
port 62 nsew signal input
rlabel metal3 s 179200 41760 180000 41880 6 adc1_dat_i[8]
port 63 nsew signal input
rlabel metal3 s 179200 46112 180000 46232 6 adc1_dat_i[9]
port 64 nsew signal input
rlabel metal3 s 179200 3544 180000 3664 6 adc2_dat_i[0]
port 65 nsew signal input
rlabel metal3 s 179200 51960 180000 52080 6 adc2_dat_i[10]
port 66 nsew signal input
rlabel metal3 s 179200 56312 180000 56432 6 adc2_dat_i[11]
port 67 nsew signal input
rlabel metal3 s 179200 60800 180000 60920 6 adc2_dat_i[12]
port 68 nsew signal input
rlabel metal3 s 179200 65152 180000 65272 6 adc2_dat_i[13]
port 69 nsew signal input
rlabel metal3 s 179200 69640 180000 69760 6 adc2_dat_i[14]
port 70 nsew signal input
rlabel metal3 s 179200 73992 180000 74112 6 adc2_dat_i[15]
port 71 nsew signal input
rlabel metal3 s 179200 78344 180000 78464 6 adc2_dat_i[16]
port 72 nsew signal input
rlabel metal3 s 179200 82832 180000 82952 6 adc2_dat_i[17]
port 73 nsew signal input
rlabel metal3 s 179200 87184 180000 87304 6 adc2_dat_i[18]
port 74 nsew signal input
rlabel metal3 s 179200 91536 180000 91656 6 adc2_dat_i[19]
port 75 nsew signal input
rlabel metal3 s 179200 9392 180000 9512 6 adc2_dat_i[1]
port 76 nsew signal input
rlabel metal3 s 179200 96024 180000 96144 6 adc2_dat_i[20]
port 77 nsew signal input
rlabel metal3 s 179200 100376 180000 100496 6 adc2_dat_i[21]
port 78 nsew signal input
rlabel metal3 s 179200 104864 180000 104984 6 adc2_dat_i[22]
port 79 nsew signal input
rlabel metal3 s 179200 109216 180000 109336 6 adc2_dat_i[23]
port 80 nsew signal input
rlabel metal3 s 179200 113568 180000 113688 6 adc2_dat_i[24]
port 81 nsew signal input
rlabel metal3 s 179200 118056 180000 118176 6 adc2_dat_i[25]
port 82 nsew signal input
rlabel metal3 s 179200 122408 180000 122528 6 adc2_dat_i[26]
port 83 nsew signal input
rlabel metal3 s 179200 126760 180000 126880 6 adc2_dat_i[27]
port 84 nsew signal input
rlabel metal3 s 179200 131248 180000 131368 6 adc2_dat_i[28]
port 85 nsew signal input
rlabel metal3 s 179200 135600 180000 135720 6 adc2_dat_i[29]
port 86 nsew signal input
rlabel metal3 s 179200 15240 180000 15360 6 adc2_dat_i[2]
port 87 nsew signal input
rlabel metal3 s 179200 139952 180000 140072 6 adc2_dat_i[30]
port 88 nsew signal input
rlabel metal3 s 179200 144440 180000 144560 6 adc2_dat_i[31]
port 89 nsew signal input
rlabel metal3 s 179200 21224 180000 21344 6 adc2_dat_i[3]
port 90 nsew signal input
rlabel metal3 s 179200 25576 180000 25696 6 adc2_dat_i[4]
port 91 nsew signal input
rlabel metal3 s 179200 29928 180000 30048 6 adc2_dat_i[5]
port 92 nsew signal input
rlabel metal3 s 179200 34416 180000 34536 6 adc2_dat_i[6]
port 93 nsew signal input
rlabel metal3 s 179200 38768 180000 38888 6 adc2_dat_i[7]
port 94 nsew signal input
rlabel metal3 s 179200 43120 180000 43240 6 adc2_dat_i[8]
port 95 nsew signal input
rlabel metal3 s 179200 47608 180000 47728 6 adc2_dat_i[9]
port 96 nsew signal input
rlabel metal3 s 179200 5040 180000 5160 6 adc_dvalid_i[0]
port 97 nsew signal input
rlabel metal3 s 179200 10888 180000 11008 6 adc_dvalid_i[1]
port 98 nsew signal input
rlabel metal3 s 179200 16736 180000 16856 6 adc_dvalid_i[2]
port 99 nsew signal input
rlabel metal2 s 1030 159200 1086 160000 6 io_oeb[0]
port 100 nsew signal output
rlabel metal2 s 44914 159200 44970 160000 6 io_oeb[10]
port 101 nsew signal output
rlabel metal2 s 49330 159200 49386 160000 6 io_oeb[11]
port 102 nsew signal output
rlabel metal2 s 53654 159200 53710 160000 6 io_oeb[12]
port 103 nsew signal output
rlabel metal2 s 58070 159200 58126 160000 6 io_oeb[13]
port 104 nsew signal output
rlabel metal2 s 62486 159200 62542 160000 6 io_oeb[14]
port 105 nsew signal output
rlabel metal2 s 66810 159200 66866 160000 6 io_oeb[15]
port 106 nsew signal output
rlabel metal2 s 71226 159200 71282 160000 6 io_oeb[16]
port 107 nsew signal output
rlabel metal2 s 75642 159200 75698 160000 6 io_oeb[17]
port 108 nsew signal output
rlabel metal2 s 80058 159200 80114 160000 6 io_oeb[18]
port 109 nsew signal output
rlabel metal2 s 84382 159200 84438 160000 6 io_oeb[19]
port 110 nsew signal output
rlabel metal2 s 5354 159200 5410 160000 6 io_oeb[1]
port 111 nsew signal output
rlabel metal2 s 88798 159200 88854 160000 6 io_oeb[20]
port 112 nsew signal output
rlabel metal2 s 93214 159200 93270 160000 6 io_oeb[21]
port 113 nsew signal output
rlabel metal2 s 97630 159200 97686 160000 6 io_oeb[22]
port 114 nsew signal output
rlabel metal2 s 101954 159200 102010 160000 6 io_oeb[23]
port 115 nsew signal output
rlabel metal2 s 106370 159200 106426 160000 6 io_oeb[24]
port 116 nsew signal output
rlabel metal2 s 110786 159200 110842 160000 6 io_oeb[25]
port 117 nsew signal output
rlabel metal2 s 115202 159200 115258 160000 6 io_oeb[26]
port 118 nsew signal output
rlabel metal2 s 119526 159200 119582 160000 6 io_oeb[27]
port 119 nsew signal output
rlabel metal2 s 123942 159200 123998 160000 6 io_oeb[28]
port 120 nsew signal output
rlabel metal2 s 128358 159200 128414 160000 6 io_oeb[29]
port 121 nsew signal output
rlabel metal2 s 9770 159200 9826 160000 6 io_oeb[2]
port 122 nsew signal output
rlabel metal2 s 132682 159200 132738 160000 6 io_oeb[30]
port 123 nsew signal output
rlabel metal2 s 137098 159200 137154 160000 6 io_oeb[31]
port 124 nsew signal output
rlabel metal2 s 141514 159200 141570 160000 6 io_oeb[32]
port 125 nsew signal output
rlabel metal2 s 145930 159200 145986 160000 6 io_oeb[33]
port 126 nsew signal output
rlabel metal2 s 150254 159200 150310 160000 6 io_oeb[34]
port 127 nsew signal output
rlabel metal2 s 154670 159200 154726 160000 6 io_oeb[35]
port 128 nsew signal output
rlabel metal2 s 159086 159200 159142 160000 6 io_oeb[36]
port 129 nsew signal output
rlabel metal2 s 163502 159200 163558 160000 6 io_oeb[37]
port 130 nsew signal output
rlabel metal2 s 14186 159200 14242 160000 6 io_oeb[3]
port 131 nsew signal output
rlabel metal2 s 18510 159200 18566 160000 6 io_oeb[4]
port 132 nsew signal output
rlabel metal2 s 22926 159200 22982 160000 6 io_oeb[5]
port 133 nsew signal output
rlabel metal2 s 27342 159200 27398 160000 6 io_oeb[6]
port 134 nsew signal output
rlabel metal2 s 31758 159200 31814 160000 6 io_oeb[7]
port 135 nsew signal output
rlabel metal2 s 36082 159200 36138 160000 6 io_oeb[8]
port 136 nsew signal output
rlabel metal2 s 40498 159200 40554 160000 6 io_oeb[9]
port 137 nsew signal output
rlabel metal2 s 3146 159200 3202 160000 6 io_out[0]
port 138 nsew signal output
rlabel metal2 s 47122 159200 47178 160000 6 io_out[10]
port 139 nsew signal output
rlabel metal2 s 51446 159200 51502 160000 6 io_out[11]
port 140 nsew signal output
rlabel metal2 s 55862 159200 55918 160000 6 io_out[12]
port 141 nsew signal output
rlabel metal2 s 60278 159200 60334 160000 6 io_out[13]
port 142 nsew signal output
rlabel metal2 s 64694 159200 64750 160000 6 io_out[14]
port 143 nsew signal output
rlabel metal2 s 69018 159200 69074 160000 6 io_out[15]
port 144 nsew signal output
rlabel metal2 s 73434 159200 73490 160000 6 io_out[16]
port 145 nsew signal output
rlabel metal2 s 77850 159200 77906 160000 6 io_out[17]
port 146 nsew signal output
rlabel metal2 s 82266 159200 82322 160000 6 io_out[18]
port 147 nsew signal output
rlabel metal2 s 86590 159200 86646 160000 6 io_out[19]
port 148 nsew signal output
rlabel metal2 s 7562 159200 7618 160000 6 io_out[1]
port 149 nsew signal output
rlabel metal2 s 91006 159200 91062 160000 6 io_out[20]
port 150 nsew signal output
rlabel metal2 s 95422 159200 95478 160000 6 io_out[21]
port 151 nsew signal output
rlabel metal2 s 99746 159200 99802 160000 6 io_out[22]
port 152 nsew signal output
rlabel metal2 s 104162 159200 104218 160000 6 io_out[23]
port 153 nsew signal output
rlabel metal2 s 108578 159200 108634 160000 6 io_out[24]
port 154 nsew signal output
rlabel metal2 s 112994 159200 113050 160000 6 io_out[25]
port 155 nsew signal output
rlabel metal2 s 117318 159200 117374 160000 6 io_out[26]
port 156 nsew signal output
rlabel metal2 s 121734 159200 121790 160000 6 io_out[27]
port 157 nsew signal output
rlabel metal2 s 126150 159200 126206 160000 6 io_out[28]
port 158 nsew signal output
rlabel metal2 s 130566 159200 130622 160000 6 io_out[29]
port 159 nsew signal output
rlabel metal2 s 11978 159200 12034 160000 6 io_out[2]
port 160 nsew signal output
rlabel metal2 s 134890 159200 134946 160000 6 io_out[30]
port 161 nsew signal output
rlabel metal2 s 139306 159200 139362 160000 6 io_out[31]
port 162 nsew signal output
rlabel metal2 s 143722 159200 143778 160000 6 io_out[32]
port 163 nsew signal output
rlabel metal2 s 148138 159200 148194 160000 6 io_out[33]
port 164 nsew signal output
rlabel metal2 s 152462 159200 152518 160000 6 io_out[34]
port 165 nsew signal output
rlabel metal2 s 156878 159200 156934 160000 6 io_out[35]
port 166 nsew signal output
rlabel metal2 s 161294 159200 161350 160000 6 io_out[36]
port 167 nsew signal output
rlabel metal2 s 165618 159200 165674 160000 6 io_out[37]
port 168 nsew signal output
rlabel metal2 s 16394 159200 16450 160000 6 io_out[3]
port 169 nsew signal output
rlabel metal2 s 20718 159200 20774 160000 6 io_out[4]
port 170 nsew signal output
rlabel metal2 s 25134 159200 25190 160000 6 io_out[5]
port 171 nsew signal output
rlabel metal2 s 29550 159200 29606 160000 6 io_out[6]
port 172 nsew signal output
rlabel metal2 s 33874 159200 33930 160000 6 io_out[7]
port 173 nsew signal output
rlabel metal2 s 38290 159200 38346 160000 6 io_out[8]
port 174 nsew signal output
rlabel metal2 s 42706 159200 42762 160000 6 io_out[9]
port 175 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 irq[0]
port 176 nsew signal output
rlabel metal2 s 177486 0 177542 800 6 irq[1]
port 177 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 irq[2]
port 178 nsew signal output
rlabel metal3 s 0 5720 800 5840 6 mem1_data_i[0]
port 179 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 mem1_data_i[10]
port 180 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 mem1_data_i[11]
port 181 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 mem1_data_i[12]
port 182 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 mem1_data_i[13]
port 183 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 mem1_data_i[14]
port 184 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 mem1_data_i[15]
port 185 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 mem1_data_i[16]
port 186 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 mem1_data_i[17]
port 187 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 mem1_data_i[18]
port 188 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 mem1_data_i[19]
port 189 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 mem1_data_i[1]
port 190 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 mem1_data_i[20]
port 191 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 mem1_data_i[21]
port 192 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 mem1_data_i[22]
port 193 nsew signal input
rlabel metal3 s 0 124992 800 125112 6 mem1_data_i[23]
port 194 nsew signal input
rlabel metal3 s 0 128936 800 129056 6 mem1_data_i[24]
port 195 nsew signal input
rlabel metal3 s 0 132880 800 133000 6 mem1_data_i[25]
port 196 nsew signal input
rlabel metal3 s 0 136824 800 136944 6 mem1_data_i[26]
port 197 nsew signal input
rlabel metal3 s 0 140768 800 140888 6 mem1_data_i[27]
port 198 nsew signal input
rlabel metal3 s 0 144712 800 144832 6 mem1_data_i[28]
port 199 nsew signal input
rlabel metal3 s 0 148656 800 148776 6 mem1_data_i[29]
port 200 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 mem1_data_i[2]
port 201 nsew signal input
rlabel metal3 s 0 152600 800 152720 6 mem1_data_i[30]
port 202 nsew signal input
rlabel metal3 s 0 156544 800 156664 6 mem1_data_i[31]
port 203 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 mem1_data_i[3]
port 204 nsew signal input
rlabel metal3 s 0 37136 800 37256 6 mem1_data_i[4]
port 205 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 mem1_data_i[5]
port 206 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 mem1_data_i[6]
port 207 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 mem1_data_i[7]
port 208 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 mem1_data_i[8]
port 209 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 mem1_data_i[9]
port 210 nsew signal input
rlabel metal3 s 0 7080 800 7200 6 mem_data_i[0]
port 211 nsew signal input
rlabel metal3 s 0 75216 800 75336 6 mem_data_i[10]
port 212 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 mem_data_i[11]
port 213 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 mem_data_i[12]
port 214 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 mem_data_i[13]
port 215 nsew signal input
rlabel metal3 s 0 90992 800 91112 6 mem_data_i[14]
port 216 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 mem_data_i[15]
port 217 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 mem_data_i[16]
port 218 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 mem_data_i[17]
port 219 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 mem_data_i[18]
port 220 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 mem_data_i[19]
port 221 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 mem_data_i[1]
port 222 nsew signal input
rlabel metal3 s 0 114520 800 114640 6 mem_data_i[20]
port 223 nsew signal input
rlabel metal3 s 0 118464 800 118584 6 mem_data_i[21]
port 224 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 mem_data_i[22]
port 225 nsew signal input
rlabel metal3 s 0 126352 800 126472 6 mem_data_i[23]
port 226 nsew signal input
rlabel metal3 s 0 130296 800 130416 6 mem_data_i[24]
port 227 nsew signal input
rlabel metal3 s 0 134240 800 134360 6 mem_data_i[25]
port 228 nsew signal input
rlabel metal3 s 0 138184 800 138304 6 mem_data_i[26]
port 229 nsew signal input
rlabel metal3 s 0 142128 800 142248 6 mem_data_i[27]
port 230 nsew signal input
rlabel metal3 s 0 145936 800 146056 6 mem_data_i[28]
port 231 nsew signal input
rlabel metal3 s 0 149880 800 150000 6 mem_data_i[29]
port 232 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 mem_data_i[2]
port 233 nsew signal input
rlabel metal3 s 0 153824 800 153944 6 mem_data_i[30]
port 234 nsew signal input
rlabel metal3 s 0 157768 800 157888 6 mem_data_i[31]
port 235 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 mem_data_i[3]
port 236 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 mem_data_i[4]
port 237 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 mem_data_i[5]
port 238 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 mem_data_i[6]
port 239 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 mem_data_i[7]
port 240 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 mem_data_i[8]
port 241 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 mem_data_i[9]
port 242 nsew signal input
rlabel metal3 s 0 8304 800 8424 6 mem_data_o[0]
port 243 nsew signal output
rlabel metal3 s 0 76576 800 76696 6 mem_data_o[10]
port 244 nsew signal output
rlabel metal3 s 0 80520 800 80640 6 mem_data_o[11]
port 245 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 mem_data_o[12]
port 246 nsew signal output
rlabel metal3 s 0 88272 800 88392 6 mem_data_o[13]
port 247 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 mem_data_o[14]
port 248 nsew signal output
rlabel metal3 s 0 96160 800 96280 6 mem_data_o[15]
port 249 nsew signal output
rlabel metal3 s 0 100104 800 100224 6 mem_data_o[16]
port 250 nsew signal output
rlabel metal3 s 0 104048 800 104168 6 mem_data_o[17]
port 251 nsew signal output
rlabel metal3 s 0 107992 800 108112 6 mem_data_o[18]
port 252 nsew signal output
rlabel metal3 s 0 111936 800 112056 6 mem_data_o[19]
port 253 nsew signal output
rlabel metal3 s 0 17552 800 17672 6 mem_data_o[1]
port 254 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 mem_data_o[20]
port 255 nsew signal output
rlabel metal3 s 0 119824 800 119944 6 mem_data_o[21]
port 256 nsew signal output
rlabel metal3 s 0 123768 800 123888 6 mem_data_o[22]
port 257 nsew signal output
rlabel metal3 s 0 127712 800 127832 6 mem_data_o[23]
port 258 nsew signal output
rlabel metal3 s 0 131520 800 131640 6 mem_data_o[24]
port 259 nsew signal output
rlabel metal3 s 0 135464 800 135584 6 mem_data_o[25]
port 260 nsew signal output
rlabel metal3 s 0 139408 800 139528 6 mem_data_o[26]
port 261 nsew signal output
rlabel metal3 s 0 143352 800 143472 6 mem_data_o[27]
port 262 nsew signal output
rlabel metal3 s 0 147296 800 147416 6 mem_data_o[28]
port 263 nsew signal output
rlabel metal3 s 0 151240 800 151360 6 mem_data_o[29]
port 264 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 mem_data_o[2]
port 265 nsew signal output
rlabel metal3 s 0 155184 800 155304 6 mem_data_o[30]
port 266 nsew signal output
rlabel metal3 s 0 159128 800 159248 6 mem_data_o[31]
port 267 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 mem_data_o[3]
port 268 nsew signal output
rlabel metal3 s 0 39856 800 39976 6 mem_data_o[4]
port 269 nsew signal output
rlabel metal3 s 0 46384 800 46504 6 mem_data_o[5]
port 270 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 mem_data_o[6]
port 271 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 mem_data_o[7]
port 272 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 mem_data_o[8]
port 273 nsew signal output
rlabel metal3 s 0 72632 800 72752 6 mem_data_o[9]
port 274 nsew signal output
rlabel metal3 s 0 9664 800 9784 6 mem_raddr_o[0]
port 275 nsew signal output
rlabel metal3 s 0 18776 800 18896 6 mem_raddr_o[1]
port 276 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 mem_raddr_o[2]
port 277 nsew signal output
rlabel metal3 s 0 34552 800 34672 6 mem_raddr_o[3]
port 278 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 mem_raddr_o[4]
port 279 nsew signal output
rlabel metal3 s 0 47744 800 47864 6 mem_raddr_o[5]
port 280 nsew signal output
rlabel metal3 s 0 54272 800 54392 6 mem_raddr_o[6]
port 281 nsew signal output
rlabel metal3 s 0 60800 800 60920 6 mem_raddr_o[7]
port 282 nsew signal output
rlabel metal3 s 0 67328 800 67448 6 mem_raddr_o[8]
port 283 nsew signal output
rlabel metal3 s 0 11024 800 11144 6 mem_renb_o[0]
port 284 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 mem_renb_o[1]
port 285 nsew signal output
rlabel metal3 s 0 12248 800 12368 6 mem_waddr_o[0]
port 286 nsew signal output
rlabel metal3 s 0 21496 800 21616 6 mem_waddr_o[1]
port 287 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 mem_waddr_o[2]
port 288 nsew signal output
rlabel metal3 s 0 35912 800 36032 6 mem_waddr_o[3]
port 289 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 mem_waddr_o[4]
port 290 nsew signal output
rlabel metal3 s 0 48968 800 49088 6 mem_waddr_o[5]
port 291 nsew signal output
rlabel metal3 s 0 55496 800 55616 6 mem_waddr_o[6]
port 292 nsew signal output
rlabel metal3 s 0 62160 800 62280 6 mem_waddr_o[7]
port 293 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 mem_waddr_o[8]
port 294 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 mem_wenb_o[0]
port 295 nsew signal output
rlabel metal3 s 0 22720 800 22840 6 mem_wenb_o[1]
port 296 nsew signal output
rlabel metal3 s 179200 145936 180000 146056 6 oversample_o[0]
port 297 nsew signal output
rlabel metal3 s 179200 147296 180000 147416 6 oversample_o[1]
port 298 nsew signal output
rlabel metal3 s 179200 148792 180000 148912 6 oversample_o[2]
port 299 nsew signal output
rlabel metal3 s 179200 150288 180000 150408 6 oversample_o[3]
port 300 nsew signal output
rlabel metal3 s 179200 151784 180000 151904 6 oversample_o[4]
port 301 nsew signal output
rlabel metal3 s 179200 153280 180000 153400 6 oversample_o[5]
port 302 nsew signal output
rlabel metal3 s 179200 154640 180000 154760 6 oversample_o[6]
port 303 nsew signal output
rlabel metal3 s 179200 156136 180000 156256 6 oversample_o[7]
port 304 nsew signal output
rlabel metal3 s 179200 157632 180000 157752 6 oversample_o[8]
port 305 nsew signal output
rlabel metal3 s 179200 159128 180000 159248 6 oversample_o[9]
port 306 nsew signal output
rlabel metal2 s 174450 159200 174506 160000 6 sinc3_en_o[0]
port 307 nsew signal output
rlabel metal2 s 176658 159200 176714 160000 6 sinc3_en_o[1]
port 308 nsew signal output
rlabel metal2 s 178866 159200 178922 160000 6 sinc3_en_o[2]
port 309 nsew signal output
rlabel metal2 s 167826 159200 167882 160000 6 vco_enb_o[0]
port 310 nsew signal output
rlabel metal2 s 170034 159200 170090 160000 6 vco_enb_o[1]
port 311 nsew signal output
rlabel metal2 s 172242 159200 172298 160000 6 vco_enb_o[2]
port 312 nsew signal output
rlabel metal2 s 754 0 810 800 6 wb_clk_i
port 313 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wb_rst_i
port 314 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_ack_o
port 315 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_adr_i[0]
port 316 nsew signal input
rlabel metal2 s 66810 0 66866 800 6 wbs_adr_i[10]
port 317 nsew signal input
rlabel metal2 s 71778 0 71834 800 6 wbs_adr_i[11]
port 318 nsew signal input
rlabel metal2 s 76654 0 76710 800 6 wbs_adr_i[12]
port 319 nsew signal input
rlabel metal2 s 81622 0 81678 800 6 wbs_adr_i[13]
port 320 nsew signal input
rlabel metal2 s 86590 0 86646 800 6 wbs_adr_i[14]
port 321 nsew signal input
rlabel metal2 s 91558 0 91614 800 6 wbs_adr_i[15]
port 322 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 wbs_adr_i[16]
port 323 nsew signal input
rlabel metal2 s 101494 0 101550 800 6 wbs_adr_i[17]
port 324 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 wbs_adr_i[18]
port 325 nsew signal input
rlabel metal2 s 111338 0 111394 800 6 wbs_adr_i[19]
port 326 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wbs_adr_i[1]
port 327 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 wbs_adr_i[20]
port 328 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 wbs_adr_i[21]
port 329 nsew signal input
rlabel metal2 s 126242 0 126298 800 6 wbs_adr_i[22]
port 330 nsew signal input
rlabel metal2 s 131210 0 131266 800 6 wbs_adr_i[23]
port 331 nsew signal input
rlabel metal2 s 136178 0 136234 800 6 wbs_adr_i[24]
port 332 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 wbs_adr_i[25]
port 333 nsew signal input
rlabel metal2 s 146022 0 146078 800 6 wbs_adr_i[26]
port 334 nsew signal input
rlabel metal2 s 150990 0 151046 800 6 wbs_adr_i[27]
port 335 nsew signal input
rlabel metal2 s 155958 0 156014 800 6 wbs_adr_i[28]
port 336 nsew signal input
rlabel metal2 s 160926 0 160982 800 6 wbs_adr_i[29]
port 337 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_adr_i[2]
port 338 nsew signal input
rlabel metal2 s 165894 0 165950 800 6 wbs_adr_i[30]
port 339 nsew signal input
rlabel metal2 s 170862 0 170918 800 6 wbs_adr_i[31]
port 340 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wbs_adr_i[3]
port 341 nsew signal input
rlabel metal2 s 37002 0 37058 800 6 wbs_adr_i[4]
port 342 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 wbs_adr_i[5]
port 343 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 wbs_adr_i[6]
port 344 nsew signal input
rlabel metal2 s 51906 0 51962 800 6 wbs_adr_i[7]
port 345 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 wbs_adr_i[8]
port 346 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 wbs_adr_i[9]
port 347 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_cyc_i
port 348 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wbs_dat_i[0]
port 349 nsew signal input
rlabel metal2 s 68466 0 68522 800 6 wbs_dat_i[10]
port 350 nsew signal input
rlabel metal2 s 73342 0 73398 800 6 wbs_dat_i[11]
port 351 nsew signal input
rlabel metal2 s 78310 0 78366 800 6 wbs_dat_i[12]
port 352 nsew signal input
rlabel metal2 s 83278 0 83334 800 6 wbs_dat_i[13]
port 353 nsew signal input
rlabel metal2 s 88246 0 88302 800 6 wbs_dat_i[14]
port 354 nsew signal input
rlabel metal2 s 93214 0 93270 800 6 wbs_dat_i[15]
port 355 nsew signal input
rlabel metal2 s 98182 0 98238 800 6 wbs_dat_i[16]
port 356 nsew signal input
rlabel metal2 s 103150 0 103206 800 6 wbs_dat_i[17]
port 357 nsew signal input
rlabel metal2 s 108118 0 108174 800 6 wbs_dat_i[18]
port 358 nsew signal input
rlabel metal2 s 112994 0 113050 800 6 wbs_dat_i[19]
port 359 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 wbs_dat_i[1]
port 360 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 wbs_dat_i[20]
port 361 nsew signal input
rlabel metal2 s 122930 0 122986 800 6 wbs_dat_i[21]
port 362 nsew signal input
rlabel metal2 s 127898 0 127954 800 6 wbs_dat_i[22]
port 363 nsew signal input
rlabel metal2 s 132866 0 132922 800 6 wbs_dat_i[23]
port 364 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 wbs_dat_i[24]
port 365 nsew signal input
rlabel metal2 s 142802 0 142858 800 6 wbs_dat_i[25]
port 366 nsew signal input
rlabel metal2 s 147678 0 147734 800 6 wbs_dat_i[26]
port 367 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 wbs_dat_i[27]
port 368 nsew signal input
rlabel metal2 s 157614 0 157670 800 6 wbs_dat_i[28]
port 369 nsew signal input
rlabel metal2 s 162582 0 162638 800 6 wbs_dat_i[29]
port 370 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_dat_i[2]
port 371 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 wbs_dat_i[30]
port 372 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 wbs_dat_i[31]
port 373 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wbs_dat_i[3]
port 374 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[4]
port 375 nsew signal input
rlabel metal2 s 43626 0 43682 800 6 wbs_dat_i[5]
port 376 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 wbs_dat_i[6]
port 377 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 wbs_dat_i[7]
port 378 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_dat_i[8]
port 379 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 wbs_dat_i[9]
port 380 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wbs_dat_o[0]
port 381 nsew signal output
rlabel metal2 s 70122 0 70178 800 6 wbs_dat_o[10]
port 382 nsew signal output
rlabel metal2 s 74998 0 75054 800 6 wbs_dat_o[11]
port 383 nsew signal output
rlabel metal2 s 79966 0 80022 800 6 wbs_dat_o[12]
port 384 nsew signal output
rlabel metal2 s 84934 0 84990 800 6 wbs_dat_o[13]
port 385 nsew signal output
rlabel metal2 s 89902 0 89958 800 6 wbs_dat_o[14]
port 386 nsew signal output
rlabel metal2 s 94870 0 94926 800 6 wbs_dat_o[15]
port 387 nsew signal output
rlabel metal2 s 99838 0 99894 800 6 wbs_dat_o[16]
port 388 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 wbs_dat_o[17]
port 389 nsew signal output
rlabel metal2 s 109682 0 109738 800 6 wbs_dat_o[18]
port 390 nsew signal output
rlabel metal2 s 114650 0 114706 800 6 wbs_dat_o[19]
port 391 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wbs_dat_o[1]
port 392 nsew signal output
rlabel metal2 s 119618 0 119674 800 6 wbs_dat_o[20]
port 393 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 wbs_dat_o[21]
port 394 nsew signal output
rlabel metal2 s 129554 0 129610 800 6 wbs_dat_o[22]
port 395 nsew signal output
rlabel metal2 s 134522 0 134578 800 6 wbs_dat_o[23]
port 396 nsew signal output
rlabel metal2 s 139490 0 139546 800 6 wbs_dat_o[24]
port 397 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 wbs_dat_o[25]
port 398 nsew signal output
rlabel metal2 s 149334 0 149390 800 6 wbs_dat_o[26]
port 399 nsew signal output
rlabel metal2 s 154302 0 154358 800 6 wbs_dat_o[27]
port 400 nsew signal output
rlabel metal2 s 159270 0 159326 800 6 wbs_dat_o[28]
port 401 nsew signal output
rlabel metal2 s 164238 0 164294 800 6 wbs_dat_o[29]
port 402 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wbs_dat_o[2]
port 403 nsew signal output
rlabel metal2 s 169206 0 169262 800 6 wbs_dat_o[30]
port 404 nsew signal output
rlabel metal2 s 174174 0 174230 800 6 wbs_dat_o[31]
port 405 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 wbs_dat_o[3]
port 406 nsew signal output
rlabel metal2 s 40314 0 40370 800 6 wbs_dat_o[4]
port 407 nsew signal output
rlabel metal2 s 45282 0 45338 800 6 wbs_dat_o[5]
port 408 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_o[6]
port 409 nsew signal output
rlabel metal2 s 55218 0 55274 800 6 wbs_dat_o[7]
port 410 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 wbs_dat_o[8]
port 411 nsew signal output
rlabel metal2 s 65154 0 65210 800 6 wbs_dat_o[9]
port 412 nsew signal output
rlabel metal2 s 15566 0 15622 800 6 wbs_sel_i[0]
port 413 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_sel_i[1]
port 414 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wbs_sel_i[2]
port 415 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_sel_i[3]
port 416 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wbs_stb_i
port 417 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_we_i
port 418 nsew signal input
rlabel metal3 s 0 552 800 672 6 wmask_o[0]
port 419 nsew signal output
rlabel metal3 s 0 1776 800 1896 6 wmask_o[1]
port 420 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 wmask_o[2]
port 421 nsew signal output
rlabel metal3 s 0 4360 800 4480 6 wmask_o[3]
port 422 nsew signal output
rlabel metal4 s 157808 2128 158128 157808 6 vccd1
port 423 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 424 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 425 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 426 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 427 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 428 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 157808 6 vssd1
port 429 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 430 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 431 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 432 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 433 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 434 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 157760 6 vccd2
port 435 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 157760 6 vccd2
port 436 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 157760 6 vccd2
port 437 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 157760 6 vccd2
port 438 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 157760 6 vccd2
port 439 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 157760 6 vccd2
port 440 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 157760 6 vssd2
port 441 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 157760 6 vssd2
port 442 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 157760 6 vssd2
port 443 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 157760 6 vssd2
port 444 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 157760 6 vssd2
port 445 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 157760 6 vssd2
port 446 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 157760 6 vdda1
port 447 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 157760 6 vdda1
port 448 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 157760 6 vdda1
port 449 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 157760 6 vdda1
port 450 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 157760 6 vdda1
port 451 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 157760 6 vdda1
port 452 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 157760 6 vssa1
port 453 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 157760 6 vssa1
port 454 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 157760 6 vssa1
port 455 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 157760 6 vssa1
port 456 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 157760 6 vssa1
port 457 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 157760 6 vssa1
port 458 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 157760 6 vdda2
port 459 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 157760 6 vdda2
port 460 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 157760 6 vdda2
port 461 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 157760 6 vdda2
port 462 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 157760 6 vdda2
port 463 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 157760 6 vdda2
port 464 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 157760 6 vssa2
port 465 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 157760 6 vssa2
port 466 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 157760 6 vssa2
port 467 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 157760 6 vssa2
port 468 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 157760 6 vssa2
port 469 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 157760 6 vssa2
port 470 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 160000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 10758504
string GDS_START 647368
<< end >>

