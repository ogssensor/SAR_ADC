VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2889.020 -9.320 2892.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2709.020 -9.320 2712.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2529.020 2584.920 2532.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2349.020 -9.320 2352.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2169.020 -9.320 2172.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1989.020 2299.760 1992.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1809.020 2299.760 1812.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1629.020 2299.760 1632.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1449.020 2299.760 1452.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1269.020 2299.760 1272.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1089.020 -9.320 1092.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 909.020 -9.320 912.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 729.020 3279.860 732.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 549.020 3279.860 552.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 369.020 3279.860 372.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 189.020 3279.860 192.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.020 -9.320 12.020 3529.000 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 729.020 -9.320 732.020 2594.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 549.020 -9.320 552.020 2594.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 369.020 -9.320 372.020 2594.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 189.020 -9.320 192.020 2594.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2529.020 2046.160 2532.020 2446.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2529.020 1505.080 2532.020 1907.640 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1989.020 -9.320 1992.020 1680.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1809.020 -9.320 1812.020 1680.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1629.020 -9.320 1632.020 1680.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1449.020 -9.320 1452.020 1680.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1269.020 -9.320 1272.020 1680.240 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2529.020 -9.320 2532.020 1366.560 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 3434.140 2934.300 3437.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 3254.140 2934.300 3257.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 3074.140 2934.300 3077.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2894.140 2934.300 2897.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2714.140 2934.300 2717.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2534.140 2934.300 2537.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2354.140 2934.300 2357.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 2174.140 2934.300 2177.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1994.140 2934.300 1997.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1814.140 2934.300 1817.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1634.140 2934.300 1637.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1454.140 2934.300 1457.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1274.140 2934.300 1277.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 1094.140 2934.300 1097.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 914.140 2934.300 917.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 734.140 2934.300 737.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 554.140 2934.300 557.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 374.140 2934.300 377.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 194.140 2934.300 197.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -14.680 14.140 2934.300 17.140 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2931.300 -9.320 2934.300 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2799.020 -9.320 2802.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2619.020 2584.920 2622.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2439.020 -9.320 2442.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2259.020 -9.320 2262.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2079.020 2299.760 2082.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1899.020 2299.760 1902.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1719.020 2299.760 1722.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1539.020 2299.760 1542.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1359.020 2299.760 1362.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1179.020 2299.760 1182.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 999.020 -9.320 1002.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 819.020 3279.860 822.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 639.020 3279.860 642.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 459.020 3279.860 462.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 279.020 3279.860 282.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 99.020 -9.320 102.020 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.680 -9.320 -11.680 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 819.020 -9.320 822.020 2594.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 639.020 -9.320 642.020 2594.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 459.020 -9.320 462.020 2594.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 279.020 -9.320 282.020 2594.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2619.020 2046.160 2622.020 2446.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2619.020 1505.080 2622.020 1907.640 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2079.020 -9.320 2082.020 1680.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1899.020 -9.320 1902.020 1680.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1719.020 -9.320 1722.020 1680.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1539.020 -9.320 1542.020 1680.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1359.020 -9.320 1362.020 1680.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1179.020 -9.320 1182.020 1680.240 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2619.020 -9.320 2622.020 1366.560 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 3526.000 2934.300 3529.000 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 3344.140 2934.300 3347.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 3164.140 2934.300 3167.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2984.140 2934.300 2987.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2804.140 2934.300 2807.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2624.140 2934.300 2627.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2444.140 2934.300 2447.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2264.140 2934.300 2267.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 2084.140 2934.300 2087.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1904.140 2934.300 1907.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1724.140 2934.300 1727.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1544.140 2934.300 1547.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1364.140 2934.300 1367.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1184.140 2934.300 1187.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 1004.140 2934.300 1007.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 824.140 2934.300 827.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 644.140 2934.300 647.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 464.140 2934.300 467.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 284.140 2934.300 287.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 104.140 2934.300 107.140 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -14.680 -9.320 2934.300 -6.320 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2907.020 -18.720 2910.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2727.020 -18.720 2730.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2547.020 2585.160 2550.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2367.020 -18.720 2370.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2187.020 -18.720 2190.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2007.020 2300.000 2010.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1827.020 2300.000 1830.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1647.020 2300.000 1650.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1467.020 2300.000 1470.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1287.020 2300.000 1290.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1107.020 -18.720 1110.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 927.020 -18.720 930.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 747.020 3280.100 750.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 567.020 3280.100 570.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 387.020 3280.100 390.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 207.020 3280.100 210.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.020 -18.720 30.020 3538.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2936.000 -14.020 2939.000 3533.700 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.380 -14.020 -16.380 3533.700 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 747.020 -18.720 750.020 2594.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 567.020 -18.720 570.020 2594.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 387.020 -18.720 390.020 2594.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 207.020 -18.720 210.020 2594.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2547.020 2046.400 2550.020 2446.160 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2547.020 1505.320 2550.020 1907.400 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2007.020 -18.720 2010.020 1680.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1827.020 -18.720 1830.020 1680.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1647.020 -18.720 1650.020 1680.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1467.020 -18.720 1470.020 1680.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1287.020 -18.720 1290.020 1680.000 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2547.020 -18.720 2550.020 1366.320 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380 3530.700 2939.000 3533.700 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 3452.380 2943.700 3455.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 3272.380 2943.700 3275.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 3092.380 2943.700 3095.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 2912.380 2943.700 2915.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 2732.380 2943.700 2735.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 2552.380 2943.700 2555.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 2372.380 2943.700 2375.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 2192.380 2943.700 2195.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 2012.380 2943.700 2015.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 1832.380 2943.700 1835.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 1652.380 2943.700 1655.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 1472.380 2943.700 1475.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 1292.380 2943.700 1295.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 1112.380 2943.700 1115.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 932.380 2943.700 935.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 752.380 2943.700 755.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 572.380 2943.700 575.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 392.380 2943.700 395.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 212.380 2943.700 215.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -24.080 32.380 2943.700 35.380 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -19.380 -14.020 2939.000 -11.020 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2940.700 -18.720 2943.700 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2817.020 -18.720 2820.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2637.020 2585.160 2640.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2457.020 -18.720 2460.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2277.020 -18.720 2280.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2097.020 -18.720 2100.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1917.020 2300.000 1920.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1737.020 2300.000 1740.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1557.020 2300.000 1560.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1377.020 2300.000 1380.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1197.020 2300.000 1200.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1017.020 -18.720 1020.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 837.020 3280.100 840.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 657.020 3280.100 660.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 477.020 3280.100 480.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 297.020 3280.100 300.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 117.020 -18.720 120.020 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.080 -18.720 -21.080 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 837.020 -18.720 840.020 2594.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 657.020 -18.720 660.020 2594.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 477.020 -18.720 480.020 2594.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 297.020 -18.720 300.020 2594.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2637.020 2046.400 2640.020 2446.160 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2637.020 1505.320 2640.020 1907.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1917.020 -18.720 1920.020 1680.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1737.020 -18.720 1740.020 1680.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1557.020 -18.720 1560.020 1680.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1377.020 -18.720 1380.020 1680.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1197.020 -18.720 1200.020 1680.000 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2637.020 -18.720 2640.020 1366.320 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 3535.400 2943.700 3538.400 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 3362.380 2943.700 3365.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 3182.380 2943.700 3185.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 3002.380 2943.700 3005.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 2822.380 2943.700 2825.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 2642.380 2943.700 2645.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 2462.380 2943.700 2465.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 2282.380 2943.700 2285.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 2102.380 2943.700 2105.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 1922.380 2943.700 1925.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 1742.380 2943.700 1745.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 1562.380 2943.700 1565.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 1382.380 2943.700 1385.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 1202.380 2943.700 1205.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 1022.380 2943.700 1025.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 842.380 2943.700 845.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 662.380 2943.700 665.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 482.380 2943.700 485.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 302.380 2943.700 305.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 122.380 2943.700 125.380 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -24.080 -18.720 2943.700 -15.720 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2745.020 -28.120 2748.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2565.020 2585.160 2568.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2385.020 -28.120 2388.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2205.020 -28.120 2208.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2025.020 2300.000 2028.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1845.020 2300.000 1848.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1665.020 2300.000 1668.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1485.020 2300.000 1488.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1305.020 2300.000 1308.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1125.020 -28.120 1128.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 945.020 -28.120 948.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 765.020 3280.100 768.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 585.020 3280.100 588.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 405.020 3280.100 408.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 225.020 3280.100 228.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 45.020 -28.120 48.020 3547.800 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2945.400 -23.420 2948.400 3543.100 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -28.780 -23.420 -25.780 3543.100 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 765.020 -28.120 768.020 2594.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 585.020 -28.120 588.020 2594.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 405.020 -28.120 408.020 2594.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 225.020 -28.120 228.020 2594.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2565.020 2046.400 2568.020 2446.160 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2565.020 1505.320 2568.020 1907.400 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2025.020 -28.120 2028.020 1680.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1845.020 -28.120 1848.020 1680.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1665.020 -28.120 1668.020 1680.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1485.020 -28.120 1488.020 1680.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1305.020 -28.120 1308.020 1680.000 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2565.020 -28.120 2568.020 1366.320 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780 3540.100 2948.400 3543.100 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 3470.380 2953.100 3473.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 3290.380 2953.100 3293.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 3110.380 2953.100 3113.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 2930.380 2953.100 2933.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 2750.380 2953.100 2753.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 2570.380 2953.100 2573.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 2390.380 2953.100 2393.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 2210.380 2953.100 2213.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 2030.380 2953.100 2033.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 1850.380 2953.100 1853.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 1670.380 2953.100 1673.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 1490.380 2953.100 1493.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 1310.380 2953.100 1313.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 1130.380 2953.100 1133.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 950.380 2953.100 953.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 770.380 2953.100 773.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 590.380 2953.100 593.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 410.380 2953.100 413.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 230.380 2953.100 233.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -33.480 50.380 2953.100 53.380 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -28.780 -23.420 2948.400 -20.420 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2950.100 -28.120 2953.100 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2835.020 -28.120 2838.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2655.020 2585.160 2658.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2475.020 -28.120 2478.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2295.020 -28.120 2298.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2115.020 -28.120 2118.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1935.020 2300.000 1938.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1755.020 2300.000 1758.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1575.020 2300.000 1578.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1395.020 2300.000 1398.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1215.020 2300.000 1218.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1035.020 -28.120 1038.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 855.020 -28.120 858.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 675.020 3280.100 678.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 495.020 3280.100 498.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 315.020 3280.100 318.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 135.020 -28.120 138.020 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -33.480 -28.120 -30.480 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 675.020 -28.120 678.020 2594.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 495.020 -28.120 498.020 2594.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 315.020 -28.120 318.020 2594.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2655.020 2046.400 2658.020 2446.160 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2655.020 1505.320 2658.020 1907.400 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1935.020 -28.120 1938.020 1680.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1755.020 -28.120 1758.020 1680.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1575.020 -28.120 1578.020 1680.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1395.020 -28.120 1398.020 1680.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1215.020 -28.120 1218.020 1680.000 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2655.020 -28.120 2658.020 1366.320 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 3544.800 2953.100 3547.800 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 3380.380 2953.100 3383.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 3200.380 2953.100 3203.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 3020.380 2953.100 3023.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 2840.380 2953.100 2843.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 2660.380 2953.100 2663.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 2480.380 2953.100 2483.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 2300.380 2953.100 2303.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 2120.380 2953.100 2123.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 1940.380 2953.100 1943.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 1760.380 2953.100 1763.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 1580.380 2953.100 1583.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 1400.380 2953.100 1403.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 1220.380 2953.100 1223.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 1040.380 2953.100 1043.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 860.380 2953.100 863.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 680.380 2953.100 683.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 500.380 2953.100 503.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 320.380 2953.100 323.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 140.380 2953.100 143.380 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -33.480 -28.120 2953.100 -25.120 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2763.020 -37.520 2766.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2583.020 2585.160 2586.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2403.020 -37.520 2406.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2223.020 -37.520 2226.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2043.020 2300.000 2046.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1863.020 2300.000 1866.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1683.020 2300.000 1686.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1503.020 2300.000 1506.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1323.020 2300.000 1326.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1143.020 -37.520 1146.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 963.020 -37.520 966.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 783.020 3280.100 786.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 603.020 3280.100 606.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 423.020 3280.100 426.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 243.020 3280.100 246.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 63.020 -37.520 66.020 3557.200 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2954.800 -32.820 2957.800 3552.500 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.180 -32.820 -35.180 3552.500 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 783.020 -37.520 786.020 2594.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 603.020 -37.520 606.020 2594.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 423.020 -37.520 426.020 2594.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 243.020 -37.520 246.020 2594.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2583.020 2046.400 2586.020 2446.160 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2583.020 1505.320 2586.020 1907.400 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2043.020 -37.520 2046.020 1680.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1863.020 -37.520 1866.020 1680.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1683.020 -37.520 1686.020 1680.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1503.020 -37.520 1506.020 1680.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1323.020 -37.520 1326.020 1680.000 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 2583.020 -37.520 2586.020 1366.320 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180 3549.500 2957.800 3552.500 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 3488.380 2962.500 3491.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 3308.380 2962.500 3311.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 3128.380 2962.500 3131.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 2948.380 2962.500 2951.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 2768.380 2962.500 2771.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 2588.380 2962.500 2591.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 2408.380 2962.500 2411.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 2228.380 2962.500 2231.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 2048.380 2962.500 2051.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 1868.380 2962.500 1871.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 1688.380 2962.500 1691.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 1508.380 2962.500 1511.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 1328.380 2962.500 1331.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 1148.380 2962.500 1151.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 968.380 2962.500 971.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 788.380 2962.500 791.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 608.380 2962.500 611.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 428.380 2962.500 431.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 248.380 2962.500 251.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -42.880 68.380 2962.500 71.380 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT -38.180 -32.820 2957.800 -29.820 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2959.500 -37.520 2962.500 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2853.020 -37.520 2856.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2673.020 2585.160 2676.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2493.020 -37.520 2496.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2313.020 -37.520 2316.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2133.020 -37.520 2136.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1953.020 2300.000 1956.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1773.020 2300.000 1776.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1593.020 2300.000 1596.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1413.020 2300.000 1416.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1233.020 2300.000 1236.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1053.020 -37.520 1056.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 873.020 -37.520 876.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 693.020 3280.100 696.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 513.020 3280.100 516.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 333.020 3280.100 336.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 153.020 3280.100 156.020 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.880 -37.520 -39.880 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 693.020 -37.520 696.020 2594.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 513.020 -37.520 516.020 2594.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 333.020 -37.520 336.020 2594.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 153.020 -37.520 156.020 2594.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2673.020 2046.400 2676.020 2446.160 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2673.020 1505.320 2676.020 1907.400 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1953.020 -37.520 1956.020 1680.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1773.020 -37.520 1776.020 1680.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1593.020 -37.520 1596.020 1680.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1413.020 -37.520 1416.020 1680.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1233.020 -37.520 1236.020 1680.000 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 2673.020 -37.520 2676.020 1366.320 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 3554.200 2962.500 3557.200 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 3398.380 2962.500 3401.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 3218.380 2962.500 3221.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 3038.380 2962.500 3041.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 2858.380 2962.500 2861.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 2678.380 2962.500 2681.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 2498.380 2962.500 2501.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 2318.380 2962.500 2321.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 2138.380 2962.500 2141.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 1958.380 2962.500 1961.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 1778.380 2962.500 1781.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 1598.380 2962.500 1601.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 1418.380 2962.500 1421.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 1238.380 2962.500 1241.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 1058.380 2962.500 1061.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 878.380 2962.500 881.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 698.380 2962.500 701.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 518.380 2962.500 521.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 338.380 2962.500 341.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 158.380 2962.500 161.380 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT -42.880 -37.520 2962.500 -34.520 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 227.385 12.665 2690.580 3284.995 ;
      LAYER met1 ;
        RECT 2.830 10.640 2914.100 3509.040 ;
      LAYER met2 ;
        RECT 2.860 3517.320 40.150 3517.600 ;
        RECT 41.270 3517.320 121.110 3517.600 ;
        RECT 122.230 3517.320 202.070 3517.600 ;
        RECT 203.190 3517.320 283.490 3517.600 ;
        RECT 284.610 3517.320 364.450 3517.600 ;
        RECT 365.570 3517.320 445.410 3517.600 ;
        RECT 446.530 3517.320 526.830 3517.600 ;
        RECT 527.950 3517.320 607.790 3517.600 ;
        RECT 608.910 3517.320 688.750 3517.600 ;
        RECT 689.870 3517.320 770.170 3517.600 ;
        RECT 771.290 3517.320 851.130 3517.600 ;
        RECT 852.250 3517.320 932.090 3517.600 ;
        RECT 933.210 3517.320 1013.510 3517.600 ;
        RECT 1014.630 3517.320 1094.470 3517.600 ;
        RECT 1095.590 3517.320 1175.430 3517.600 ;
        RECT 1176.550 3517.320 1256.850 3517.600 ;
        RECT 1257.970 3517.320 1337.810 3517.600 ;
        RECT 1338.930 3517.320 1418.770 3517.600 ;
        RECT 1419.890 3517.320 1500.190 3517.600 ;
        RECT 1501.310 3517.320 1581.150 3517.600 ;
        RECT 1582.270 3517.320 1662.110 3517.600 ;
        RECT 1663.230 3517.320 1743.530 3517.600 ;
        RECT 1744.650 3517.320 1824.490 3517.600 ;
        RECT 1825.610 3517.320 1905.450 3517.600 ;
        RECT 1906.570 3517.320 1986.870 3517.600 ;
        RECT 1987.990 3517.320 2067.830 3517.600 ;
        RECT 2068.950 3517.320 2148.790 3517.600 ;
        RECT 2149.910 3517.320 2230.210 3517.600 ;
        RECT 2231.330 3517.320 2311.170 3517.600 ;
        RECT 2312.290 3517.320 2392.130 3517.600 ;
        RECT 2393.250 3517.320 2473.550 3517.600 ;
        RECT 2474.670 3517.320 2554.510 3517.600 ;
        RECT 2555.630 3517.320 2635.470 3517.600 ;
        RECT 2636.590 3517.320 2716.890 3517.600 ;
        RECT 2718.010 3517.320 2797.850 3517.600 ;
        RECT 2798.970 3517.320 2878.810 3517.600 ;
        RECT 2879.930 3517.320 2917.160 3517.600 ;
        RECT 2.860 2.680 2917.160 3517.320 ;
        RECT 3.550 2.400 7.950 2.680 ;
        RECT 9.070 2.400 13.930 2.680 ;
        RECT 15.050 2.400 19.910 2.680 ;
        RECT 21.030 2.400 25.890 2.680 ;
        RECT 27.010 2.400 31.870 2.680 ;
        RECT 32.990 2.400 37.850 2.680 ;
        RECT 38.970 2.400 43.370 2.680 ;
        RECT 44.490 2.400 49.350 2.680 ;
        RECT 50.470 2.400 55.330 2.680 ;
        RECT 56.450 2.400 61.310 2.680 ;
        RECT 62.430 2.400 67.290 2.680 ;
        RECT 68.410 2.400 73.270 2.680 ;
        RECT 74.390 2.400 79.250 2.680 ;
        RECT 80.370 2.400 84.770 2.680 ;
        RECT 85.890 2.400 90.750 2.680 ;
        RECT 91.870 2.400 96.730 2.680 ;
        RECT 97.850 2.400 102.710 2.680 ;
        RECT 103.830 2.400 108.690 2.680 ;
        RECT 109.810 2.400 114.670 2.680 ;
        RECT 115.790 2.400 120.650 2.680 ;
        RECT 121.770 2.400 126.170 2.680 ;
        RECT 127.290 2.400 132.150 2.680 ;
        RECT 133.270 2.400 138.130 2.680 ;
        RECT 139.250 2.400 144.110 2.680 ;
        RECT 145.230 2.400 150.090 2.680 ;
        RECT 151.210 2.400 156.070 2.680 ;
        RECT 157.190 2.400 161.590 2.680 ;
        RECT 162.710 2.400 167.570 2.680 ;
        RECT 168.690 2.400 173.550 2.680 ;
        RECT 174.670 2.400 179.530 2.680 ;
        RECT 180.650 2.400 185.510 2.680 ;
        RECT 186.630 2.400 191.490 2.680 ;
        RECT 192.610 2.400 197.470 2.680 ;
        RECT 198.590 2.400 202.990 2.680 ;
        RECT 204.110 2.400 208.970 2.680 ;
        RECT 210.090 2.400 214.950 2.680 ;
        RECT 216.070 2.400 220.930 2.680 ;
        RECT 222.050 2.400 226.910 2.680 ;
        RECT 228.030 2.400 232.890 2.680 ;
        RECT 234.010 2.400 238.870 2.680 ;
        RECT 239.990 2.400 244.390 2.680 ;
        RECT 245.510 2.400 250.370 2.680 ;
        RECT 251.490 2.400 256.350 2.680 ;
        RECT 257.470 2.400 262.330 2.680 ;
        RECT 263.450 2.400 268.310 2.680 ;
        RECT 269.430 2.400 274.290 2.680 ;
        RECT 275.410 2.400 279.810 2.680 ;
        RECT 280.930 2.400 285.790 2.680 ;
        RECT 286.910 2.400 291.770 2.680 ;
        RECT 292.890 2.400 297.750 2.680 ;
        RECT 298.870 2.400 303.730 2.680 ;
        RECT 304.850 2.400 309.710 2.680 ;
        RECT 310.830 2.400 315.690 2.680 ;
        RECT 316.810 2.400 321.210 2.680 ;
        RECT 322.330 2.400 327.190 2.680 ;
        RECT 328.310 2.400 333.170 2.680 ;
        RECT 334.290 2.400 339.150 2.680 ;
        RECT 340.270 2.400 345.130 2.680 ;
        RECT 346.250 2.400 351.110 2.680 ;
        RECT 352.230 2.400 357.090 2.680 ;
        RECT 358.210 2.400 362.610 2.680 ;
        RECT 363.730 2.400 368.590 2.680 ;
        RECT 369.710 2.400 374.570 2.680 ;
        RECT 375.690 2.400 380.550 2.680 ;
        RECT 381.670 2.400 386.530 2.680 ;
        RECT 387.650 2.400 392.510 2.680 ;
        RECT 393.630 2.400 398.030 2.680 ;
        RECT 399.150 2.400 404.010 2.680 ;
        RECT 405.130 2.400 409.990 2.680 ;
        RECT 411.110 2.400 415.970 2.680 ;
        RECT 417.090 2.400 421.950 2.680 ;
        RECT 423.070 2.400 427.930 2.680 ;
        RECT 429.050 2.400 433.910 2.680 ;
        RECT 435.030 2.400 439.430 2.680 ;
        RECT 440.550 2.400 445.410 2.680 ;
        RECT 446.530 2.400 451.390 2.680 ;
        RECT 452.510 2.400 457.370 2.680 ;
        RECT 458.490 2.400 463.350 2.680 ;
        RECT 464.470 2.400 469.330 2.680 ;
        RECT 470.450 2.400 475.310 2.680 ;
        RECT 476.430 2.400 480.830 2.680 ;
        RECT 481.950 2.400 486.810 2.680 ;
        RECT 487.930 2.400 492.790 2.680 ;
        RECT 493.910 2.400 498.770 2.680 ;
        RECT 499.890 2.400 504.750 2.680 ;
        RECT 505.870 2.400 510.730 2.680 ;
        RECT 511.850 2.400 516.250 2.680 ;
        RECT 517.370 2.400 522.230 2.680 ;
        RECT 523.350 2.400 528.210 2.680 ;
        RECT 529.330 2.400 534.190 2.680 ;
        RECT 535.310 2.400 540.170 2.680 ;
        RECT 541.290 2.400 546.150 2.680 ;
        RECT 547.270 2.400 552.130 2.680 ;
        RECT 553.250 2.400 557.650 2.680 ;
        RECT 558.770 2.400 563.630 2.680 ;
        RECT 564.750 2.400 569.610 2.680 ;
        RECT 570.730 2.400 575.590 2.680 ;
        RECT 576.710 2.400 581.570 2.680 ;
        RECT 582.690 2.400 587.550 2.680 ;
        RECT 588.670 2.400 593.530 2.680 ;
        RECT 594.650 2.400 599.050 2.680 ;
        RECT 600.170 2.400 605.030 2.680 ;
        RECT 606.150 2.400 611.010 2.680 ;
        RECT 612.130 2.400 616.990 2.680 ;
        RECT 618.110 2.400 622.970 2.680 ;
        RECT 624.090 2.400 628.950 2.680 ;
        RECT 630.070 2.400 634.470 2.680 ;
        RECT 635.590 2.400 640.450 2.680 ;
        RECT 641.570 2.400 646.430 2.680 ;
        RECT 647.550 2.400 652.410 2.680 ;
        RECT 653.530 2.400 658.390 2.680 ;
        RECT 659.510 2.400 664.370 2.680 ;
        RECT 665.490 2.400 670.350 2.680 ;
        RECT 671.470 2.400 675.870 2.680 ;
        RECT 676.990 2.400 681.850 2.680 ;
        RECT 682.970 2.400 687.830 2.680 ;
        RECT 688.950 2.400 693.810 2.680 ;
        RECT 694.930 2.400 699.790 2.680 ;
        RECT 700.910 2.400 705.770 2.680 ;
        RECT 706.890 2.400 711.750 2.680 ;
        RECT 712.870 2.400 717.270 2.680 ;
        RECT 718.390 2.400 723.250 2.680 ;
        RECT 724.370 2.400 729.230 2.680 ;
        RECT 730.350 2.400 735.210 2.680 ;
        RECT 736.330 2.400 741.190 2.680 ;
        RECT 742.310 2.400 747.170 2.680 ;
        RECT 748.290 2.400 752.690 2.680 ;
        RECT 753.810 2.400 758.670 2.680 ;
        RECT 759.790 2.400 764.650 2.680 ;
        RECT 765.770 2.400 770.630 2.680 ;
        RECT 771.750 2.400 776.610 2.680 ;
        RECT 777.730 2.400 782.590 2.680 ;
        RECT 783.710 2.400 788.570 2.680 ;
        RECT 789.690 2.400 794.090 2.680 ;
        RECT 795.210 2.400 800.070 2.680 ;
        RECT 801.190 2.400 806.050 2.680 ;
        RECT 807.170 2.400 812.030 2.680 ;
        RECT 813.150 2.400 818.010 2.680 ;
        RECT 819.130 2.400 823.990 2.680 ;
        RECT 825.110 2.400 829.970 2.680 ;
        RECT 831.090 2.400 835.490 2.680 ;
        RECT 836.610 2.400 841.470 2.680 ;
        RECT 842.590 2.400 847.450 2.680 ;
        RECT 848.570 2.400 853.430 2.680 ;
        RECT 854.550 2.400 859.410 2.680 ;
        RECT 860.530 2.400 865.390 2.680 ;
        RECT 866.510 2.400 870.910 2.680 ;
        RECT 872.030 2.400 876.890 2.680 ;
        RECT 878.010 2.400 882.870 2.680 ;
        RECT 883.990 2.400 888.850 2.680 ;
        RECT 889.970 2.400 894.830 2.680 ;
        RECT 895.950 2.400 900.810 2.680 ;
        RECT 901.930 2.400 906.790 2.680 ;
        RECT 907.910 2.400 912.310 2.680 ;
        RECT 913.430 2.400 918.290 2.680 ;
        RECT 919.410 2.400 924.270 2.680 ;
        RECT 925.390 2.400 930.250 2.680 ;
        RECT 931.370 2.400 936.230 2.680 ;
        RECT 937.350 2.400 942.210 2.680 ;
        RECT 943.330 2.400 948.190 2.680 ;
        RECT 949.310 2.400 953.710 2.680 ;
        RECT 954.830 2.400 959.690 2.680 ;
        RECT 960.810 2.400 965.670 2.680 ;
        RECT 966.790 2.400 971.650 2.680 ;
        RECT 972.770 2.400 977.630 2.680 ;
        RECT 978.750 2.400 983.610 2.680 ;
        RECT 984.730 2.400 989.130 2.680 ;
        RECT 990.250 2.400 995.110 2.680 ;
        RECT 996.230 2.400 1001.090 2.680 ;
        RECT 1002.210 2.400 1007.070 2.680 ;
        RECT 1008.190 2.400 1013.050 2.680 ;
        RECT 1014.170 2.400 1019.030 2.680 ;
        RECT 1020.150 2.400 1025.010 2.680 ;
        RECT 1026.130 2.400 1030.530 2.680 ;
        RECT 1031.650 2.400 1036.510 2.680 ;
        RECT 1037.630 2.400 1042.490 2.680 ;
        RECT 1043.610 2.400 1048.470 2.680 ;
        RECT 1049.590 2.400 1054.450 2.680 ;
        RECT 1055.570 2.400 1060.430 2.680 ;
        RECT 1061.550 2.400 1066.410 2.680 ;
        RECT 1067.530 2.400 1071.930 2.680 ;
        RECT 1073.050 2.400 1077.910 2.680 ;
        RECT 1079.030 2.400 1083.890 2.680 ;
        RECT 1085.010 2.400 1089.870 2.680 ;
        RECT 1090.990 2.400 1095.850 2.680 ;
        RECT 1096.970 2.400 1101.830 2.680 ;
        RECT 1102.950 2.400 1107.350 2.680 ;
        RECT 1108.470 2.400 1113.330 2.680 ;
        RECT 1114.450 2.400 1119.310 2.680 ;
        RECT 1120.430 2.400 1125.290 2.680 ;
        RECT 1126.410 2.400 1131.270 2.680 ;
        RECT 1132.390 2.400 1137.250 2.680 ;
        RECT 1138.370 2.400 1143.230 2.680 ;
        RECT 1144.350 2.400 1148.750 2.680 ;
        RECT 1149.870 2.400 1154.730 2.680 ;
        RECT 1155.850 2.400 1160.710 2.680 ;
        RECT 1161.830 2.400 1166.690 2.680 ;
        RECT 1167.810 2.400 1172.670 2.680 ;
        RECT 1173.790 2.400 1178.650 2.680 ;
        RECT 1179.770 2.400 1184.630 2.680 ;
        RECT 1185.750 2.400 1190.150 2.680 ;
        RECT 1191.270 2.400 1196.130 2.680 ;
        RECT 1197.250 2.400 1202.110 2.680 ;
        RECT 1203.230 2.400 1208.090 2.680 ;
        RECT 1209.210 2.400 1214.070 2.680 ;
        RECT 1215.190 2.400 1220.050 2.680 ;
        RECT 1221.170 2.400 1225.570 2.680 ;
        RECT 1226.690 2.400 1231.550 2.680 ;
        RECT 1232.670 2.400 1237.530 2.680 ;
        RECT 1238.650 2.400 1243.510 2.680 ;
        RECT 1244.630 2.400 1249.490 2.680 ;
        RECT 1250.610 2.400 1255.470 2.680 ;
        RECT 1256.590 2.400 1261.450 2.680 ;
        RECT 1262.570 2.400 1266.970 2.680 ;
        RECT 1268.090 2.400 1272.950 2.680 ;
        RECT 1274.070 2.400 1278.930 2.680 ;
        RECT 1280.050 2.400 1284.910 2.680 ;
        RECT 1286.030 2.400 1290.890 2.680 ;
        RECT 1292.010 2.400 1296.870 2.680 ;
        RECT 1297.990 2.400 1302.850 2.680 ;
        RECT 1303.970 2.400 1308.370 2.680 ;
        RECT 1309.490 2.400 1314.350 2.680 ;
        RECT 1315.470 2.400 1320.330 2.680 ;
        RECT 1321.450 2.400 1326.310 2.680 ;
        RECT 1327.430 2.400 1332.290 2.680 ;
        RECT 1333.410 2.400 1338.270 2.680 ;
        RECT 1339.390 2.400 1343.790 2.680 ;
        RECT 1344.910 2.400 1349.770 2.680 ;
        RECT 1350.890 2.400 1355.750 2.680 ;
        RECT 1356.870 2.400 1361.730 2.680 ;
        RECT 1362.850 2.400 1367.710 2.680 ;
        RECT 1368.830 2.400 1373.690 2.680 ;
        RECT 1374.810 2.400 1379.670 2.680 ;
        RECT 1380.790 2.400 1385.190 2.680 ;
        RECT 1386.310 2.400 1391.170 2.680 ;
        RECT 1392.290 2.400 1397.150 2.680 ;
        RECT 1398.270 2.400 1403.130 2.680 ;
        RECT 1404.250 2.400 1409.110 2.680 ;
        RECT 1410.230 2.400 1415.090 2.680 ;
        RECT 1416.210 2.400 1421.070 2.680 ;
        RECT 1422.190 2.400 1426.590 2.680 ;
        RECT 1427.710 2.400 1432.570 2.680 ;
        RECT 1433.690 2.400 1438.550 2.680 ;
        RECT 1439.670 2.400 1444.530 2.680 ;
        RECT 1445.650 2.400 1450.510 2.680 ;
        RECT 1451.630 2.400 1456.490 2.680 ;
        RECT 1457.610 2.400 1462.470 2.680 ;
        RECT 1463.590 2.400 1467.990 2.680 ;
        RECT 1469.110 2.400 1473.970 2.680 ;
        RECT 1475.090 2.400 1479.950 2.680 ;
        RECT 1481.070 2.400 1485.930 2.680 ;
        RECT 1487.050 2.400 1491.910 2.680 ;
        RECT 1493.030 2.400 1497.890 2.680 ;
        RECT 1499.010 2.400 1503.410 2.680 ;
        RECT 1504.530 2.400 1509.390 2.680 ;
        RECT 1510.510 2.400 1515.370 2.680 ;
        RECT 1516.490 2.400 1521.350 2.680 ;
        RECT 1522.470 2.400 1527.330 2.680 ;
        RECT 1528.450 2.400 1533.310 2.680 ;
        RECT 1534.430 2.400 1539.290 2.680 ;
        RECT 1540.410 2.400 1544.810 2.680 ;
        RECT 1545.930 2.400 1550.790 2.680 ;
        RECT 1551.910 2.400 1556.770 2.680 ;
        RECT 1557.890 2.400 1562.750 2.680 ;
        RECT 1563.870 2.400 1568.730 2.680 ;
        RECT 1569.850 2.400 1574.710 2.680 ;
        RECT 1575.830 2.400 1580.690 2.680 ;
        RECT 1581.810 2.400 1586.210 2.680 ;
        RECT 1587.330 2.400 1592.190 2.680 ;
        RECT 1593.310 2.400 1598.170 2.680 ;
        RECT 1599.290 2.400 1604.150 2.680 ;
        RECT 1605.270 2.400 1610.130 2.680 ;
        RECT 1611.250 2.400 1616.110 2.680 ;
        RECT 1617.230 2.400 1621.630 2.680 ;
        RECT 1622.750 2.400 1627.610 2.680 ;
        RECT 1628.730 2.400 1633.590 2.680 ;
        RECT 1634.710 2.400 1639.570 2.680 ;
        RECT 1640.690 2.400 1645.550 2.680 ;
        RECT 1646.670 2.400 1651.530 2.680 ;
        RECT 1652.650 2.400 1657.510 2.680 ;
        RECT 1658.630 2.400 1663.030 2.680 ;
        RECT 1664.150 2.400 1669.010 2.680 ;
        RECT 1670.130 2.400 1674.990 2.680 ;
        RECT 1676.110 2.400 1680.970 2.680 ;
        RECT 1682.090 2.400 1686.950 2.680 ;
        RECT 1688.070 2.400 1692.930 2.680 ;
        RECT 1694.050 2.400 1698.910 2.680 ;
        RECT 1700.030 2.400 1704.430 2.680 ;
        RECT 1705.550 2.400 1710.410 2.680 ;
        RECT 1711.530 2.400 1716.390 2.680 ;
        RECT 1717.510 2.400 1722.370 2.680 ;
        RECT 1723.490 2.400 1728.350 2.680 ;
        RECT 1729.470 2.400 1734.330 2.680 ;
        RECT 1735.450 2.400 1739.850 2.680 ;
        RECT 1740.970 2.400 1745.830 2.680 ;
        RECT 1746.950 2.400 1751.810 2.680 ;
        RECT 1752.930 2.400 1757.790 2.680 ;
        RECT 1758.910 2.400 1763.770 2.680 ;
        RECT 1764.890 2.400 1769.750 2.680 ;
        RECT 1770.870 2.400 1775.730 2.680 ;
        RECT 1776.850 2.400 1781.250 2.680 ;
        RECT 1782.370 2.400 1787.230 2.680 ;
        RECT 1788.350 2.400 1793.210 2.680 ;
        RECT 1794.330 2.400 1799.190 2.680 ;
        RECT 1800.310 2.400 1805.170 2.680 ;
        RECT 1806.290 2.400 1811.150 2.680 ;
        RECT 1812.270 2.400 1817.130 2.680 ;
        RECT 1818.250 2.400 1822.650 2.680 ;
        RECT 1823.770 2.400 1828.630 2.680 ;
        RECT 1829.750 2.400 1834.610 2.680 ;
        RECT 1835.730 2.400 1840.590 2.680 ;
        RECT 1841.710 2.400 1846.570 2.680 ;
        RECT 1847.690 2.400 1852.550 2.680 ;
        RECT 1853.670 2.400 1858.070 2.680 ;
        RECT 1859.190 2.400 1864.050 2.680 ;
        RECT 1865.170 2.400 1870.030 2.680 ;
        RECT 1871.150 2.400 1876.010 2.680 ;
        RECT 1877.130 2.400 1881.990 2.680 ;
        RECT 1883.110 2.400 1887.970 2.680 ;
        RECT 1889.090 2.400 1893.950 2.680 ;
        RECT 1895.070 2.400 1899.470 2.680 ;
        RECT 1900.590 2.400 1905.450 2.680 ;
        RECT 1906.570 2.400 1911.430 2.680 ;
        RECT 1912.550 2.400 1917.410 2.680 ;
        RECT 1918.530 2.400 1923.390 2.680 ;
        RECT 1924.510 2.400 1929.370 2.680 ;
        RECT 1930.490 2.400 1935.350 2.680 ;
        RECT 1936.470 2.400 1940.870 2.680 ;
        RECT 1941.990 2.400 1946.850 2.680 ;
        RECT 1947.970 2.400 1952.830 2.680 ;
        RECT 1953.950 2.400 1958.810 2.680 ;
        RECT 1959.930 2.400 1964.790 2.680 ;
        RECT 1965.910 2.400 1970.770 2.680 ;
        RECT 1971.890 2.400 1976.290 2.680 ;
        RECT 1977.410 2.400 1982.270 2.680 ;
        RECT 1983.390 2.400 1988.250 2.680 ;
        RECT 1989.370 2.400 1994.230 2.680 ;
        RECT 1995.350 2.400 2000.210 2.680 ;
        RECT 2001.330 2.400 2006.190 2.680 ;
        RECT 2007.310 2.400 2012.170 2.680 ;
        RECT 2013.290 2.400 2017.690 2.680 ;
        RECT 2018.810 2.400 2023.670 2.680 ;
        RECT 2024.790 2.400 2029.650 2.680 ;
        RECT 2030.770 2.400 2035.630 2.680 ;
        RECT 2036.750 2.400 2041.610 2.680 ;
        RECT 2042.730 2.400 2047.590 2.680 ;
        RECT 2048.710 2.400 2053.570 2.680 ;
        RECT 2054.690 2.400 2059.090 2.680 ;
        RECT 2060.210 2.400 2065.070 2.680 ;
        RECT 2066.190 2.400 2071.050 2.680 ;
        RECT 2072.170 2.400 2077.030 2.680 ;
        RECT 2078.150 2.400 2083.010 2.680 ;
        RECT 2084.130 2.400 2088.990 2.680 ;
        RECT 2090.110 2.400 2094.510 2.680 ;
        RECT 2095.630 2.400 2100.490 2.680 ;
        RECT 2101.610 2.400 2106.470 2.680 ;
        RECT 2107.590 2.400 2112.450 2.680 ;
        RECT 2113.570 2.400 2118.430 2.680 ;
        RECT 2119.550 2.400 2124.410 2.680 ;
        RECT 2125.530 2.400 2130.390 2.680 ;
        RECT 2131.510 2.400 2135.910 2.680 ;
        RECT 2137.030 2.400 2141.890 2.680 ;
        RECT 2143.010 2.400 2147.870 2.680 ;
        RECT 2148.990 2.400 2153.850 2.680 ;
        RECT 2154.970 2.400 2159.830 2.680 ;
        RECT 2160.950 2.400 2165.810 2.680 ;
        RECT 2166.930 2.400 2171.790 2.680 ;
        RECT 2172.910 2.400 2177.310 2.680 ;
        RECT 2178.430 2.400 2183.290 2.680 ;
        RECT 2184.410 2.400 2189.270 2.680 ;
        RECT 2190.390 2.400 2195.250 2.680 ;
        RECT 2196.370 2.400 2201.230 2.680 ;
        RECT 2202.350 2.400 2207.210 2.680 ;
        RECT 2208.330 2.400 2212.730 2.680 ;
        RECT 2213.850 2.400 2218.710 2.680 ;
        RECT 2219.830 2.400 2224.690 2.680 ;
        RECT 2225.810 2.400 2230.670 2.680 ;
        RECT 2231.790 2.400 2236.650 2.680 ;
        RECT 2237.770 2.400 2242.630 2.680 ;
        RECT 2243.750 2.400 2248.610 2.680 ;
        RECT 2249.730 2.400 2254.130 2.680 ;
        RECT 2255.250 2.400 2260.110 2.680 ;
        RECT 2261.230 2.400 2266.090 2.680 ;
        RECT 2267.210 2.400 2272.070 2.680 ;
        RECT 2273.190 2.400 2278.050 2.680 ;
        RECT 2279.170 2.400 2284.030 2.680 ;
        RECT 2285.150 2.400 2290.010 2.680 ;
        RECT 2291.130 2.400 2295.530 2.680 ;
        RECT 2296.650 2.400 2301.510 2.680 ;
        RECT 2302.630 2.400 2307.490 2.680 ;
        RECT 2308.610 2.400 2313.470 2.680 ;
        RECT 2314.590 2.400 2319.450 2.680 ;
        RECT 2320.570 2.400 2325.430 2.680 ;
        RECT 2326.550 2.400 2330.950 2.680 ;
        RECT 2332.070 2.400 2336.930 2.680 ;
        RECT 2338.050 2.400 2342.910 2.680 ;
        RECT 2344.030 2.400 2348.890 2.680 ;
        RECT 2350.010 2.400 2354.870 2.680 ;
        RECT 2355.990 2.400 2360.850 2.680 ;
        RECT 2361.970 2.400 2366.830 2.680 ;
        RECT 2367.950 2.400 2372.350 2.680 ;
        RECT 2373.470 2.400 2378.330 2.680 ;
        RECT 2379.450 2.400 2384.310 2.680 ;
        RECT 2385.430 2.400 2390.290 2.680 ;
        RECT 2391.410 2.400 2396.270 2.680 ;
        RECT 2397.390 2.400 2402.250 2.680 ;
        RECT 2403.370 2.400 2408.230 2.680 ;
        RECT 2409.350 2.400 2413.750 2.680 ;
        RECT 2414.870 2.400 2419.730 2.680 ;
        RECT 2420.850 2.400 2425.710 2.680 ;
        RECT 2426.830 2.400 2431.690 2.680 ;
        RECT 2432.810 2.400 2437.670 2.680 ;
        RECT 2438.790 2.400 2443.650 2.680 ;
        RECT 2444.770 2.400 2449.170 2.680 ;
        RECT 2450.290 2.400 2455.150 2.680 ;
        RECT 2456.270 2.400 2461.130 2.680 ;
        RECT 2462.250 2.400 2467.110 2.680 ;
        RECT 2468.230 2.400 2473.090 2.680 ;
        RECT 2474.210 2.400 2479.070 2.680 ;
        RECT 2480.190 2.400 2485.050 2.680 ;
        RECT 2486.170 2.400 2490.570 2.680 ;
        RECT 2491.690 2.400 2496.550 2.680 ;
        RECT 2497.670 2.400 2502.530 2.680 ;
        RECT 2503.650 2.400 2508.510 2.680 ;
        RECT 2509.630 2.400 2514.490 2.680 ;
        RECT 2515.610 2.400 2520.470 2.680 ;
        RECT 2521.590 2.400 2526.450 2.680 ;
        RECT 2527.570 2.400 2531.970 2.680 ;
        RECT 2533.090 2.400 2537.950 2.680 ;
        RECT 2539.070 2.400 2543.930 2.680 ;
        RECT 2545.050 2.400 2549.910 2.680 ;
        RECT 2551.030 2.400 2555.890 2.680 ;
        RECT 2557.010 2.400 2561.870 2.680 ;
        RECT 2562.990 2.400 2567.390 2.680 ;
        RECT 2568.510 2.400 2573.370 2.680 ;
        RECT 2574.490 2.400 2579.350 2.680 ;
        RECT 2580.470 2.400 2585.330 2.680 ;
        RECT 2586.450 2.400 2591.310 2.680 ;
        RECT 2592.430 2.400 2597.290 2.680 ;
        RECT 2598.410 2.400 2603.270 2.680 ;
        RECT 2604.390 2.400 2608.790 2.680 ;
        RECT 2609.910 2.400 2614.770 2.680 ;
        RECT 2615.890 2.400 2620.750 2.680 ;
        RECT 2621.870 2.400 2626.730 2.680 ;
        RECT 2627.850 2.400 2632.710 2.680 ;
        RECT 2633.830 2.400 2638.690 2.680 ;
        RECT 2639.810 2.400 2644.670 2.680 ;
        RECT 2645.790 2.400 2650.190 2.680 ;
        RECT 2651.310 2.400 2656.170 2.680 ;
        RECT 2657.290 2.400 2662.150 2.680 ;
        RECT 2663.270 2.400 2668.130 2.680 ;
        RECT 2669.250 2.400 2674.110 2.680 ;
        RECT 2675.230 2.400 2680.090 2.680 ;
        RECT 2681.210 2.400 2685.610 2.680 ;
        RECT 2686.730 2.400 2691.590 2.680 ;
        RECT 2692.710 2.400 2697.570 2.680 ;
        RECT 2698.690 2.400 2703.550 2.680 ;
        RECT 2704.670 2.400 2709.530 2.680 ;
        RECT 2710.650 2.400 2715.510 2.680 ;
        RECT 2716.630 2.400 2721.490 2.680 ;
        RECT 2722.610 2.400 2727.010 2.680 ;
        RECT 2728.130 2.400 2732.990 2.680 ;
        RECT 2734.110 2.400 2738.970 2.680 ;
        RECT 2740.090 2.400 2744.950 2.680 ;
        RECT 2746.070 2.400 2750.930 2.680 ;
        RECT 2752.050 2.400 2756.910 2.680 ;
        RECT 2758.030 2.400 2762.890 2.680 ;
        RECT 2764.010 2.400 2768.410 2.680 ;
        RECT 2769.530 2.400 2774.390 2.680 ;
        RECT 2775.510 2.400 2780.370 2.680 ;
        RECT 2781.490 2.400 2786.350 2.680 ;
        RECT 2787.470 2.400 2792.330 2.680 ;
        RECT 2793.450 2.400 2798.310 2.680 ;
        RECT 2799.430 2.400 2803.830 2.680 ;
        RECT 2804.950 2.400 2809.810 2.680 ;
        RECT 2810.930 2.400 2815.790 2.680 ;
        RECT 2816.910 2.400 2821.770 2.680 ;
        RECT 2822.890 2.400 2827.750 2.680 ;
        RECT 2828.870 2.400 2833.730 2.680 ;
        RECT 2834.850 2.400 2839.710 2.680 ;
        RECT 2840.830 2.400 2845.230 2.680 ;
        RECT 2846.350 2.400 2851.210 2.680 ;
        RECT 2852.330 2.400 2857.190 2.680 ;
        RECT 2858.310 2.400 2863.170 2.680 ;
        RECT 2864.290 2.400 2869.150 2.680 ;
        RECT 2870.270 2.400 2875.130 2.680 ;
        RECT 2876.250 2.400 2881.110 2.680 ;
        RECT 2882.230 2.400 2886.630 2.680 ;
        RECT 2887.750 2.400 2892.610 2.680 ;
        RECT 2893.730 2.400 2898.590 2.680 ;
        RECT 2899.710 2.400 2904.570 2.680 ;
        RECT 2905.690 2.400 2910.550 2.680 ;
        RECT 2911.670 2.400 2916.530 2.680 ;
      LAYER met3 ;
        RECT 2.400 3487.700 2917.600 3508.965 ;
        RECT 2.800 3487.020 2917.600 3487.700 ;
        RECT 2.800 3485.700 2917.200 3487.020 ;
        RECT 2.400 3485.020 2917.200 3485.700 ;
        RECT 2.400 3422.420 2917.600 3485.020 ;
        RECT 2.800 3420.420 2917.600 3422.420 ;
        RECT 2.400 3420.380 2917.600 3420.420 ;
        RECT 2.400 3418.380 2917.200 3420.380 ;
        RECT 2.400 3357.140 2917.600 3418.380 ;
        RECT 2.800 3355.140 2917.600 3357.140 ;
        RECT 2.400 3354.420 2917.600 3355.140 ;
        RECT 2.400 3352.420 2917.200 3354.420 ;
        RECT 2.400 3291.860 2917.600 3352.420 ;
        RECT 2.800 3289.860 2917.600 3291.860 ;
        RECT 2.400 3287.780 2917.600 3289.860 ;
        RECT 2.400 3285.780 2917.200 3287.780 ;
        RECT 2.400 3226.580 2917.600 3285.780 ;
        RECT 2.800 3224.580 2917.600 3226.580 ;
        RECT 2.400 3221.140 2917.600 3224.580 ;
        RECT 2.400 3219.140 2917.200 3221.140 ;
        RECT 2.400 3161.300 2917.600 3219.140 ;
        RECT 2.800 3159.300 2917.600 3161.300 ;
        RECT 2.400 3155.180 2917.600 3159.300 ;
        RECT 2.400 3153.180 2917.200 3155.180 ;
        RECT 2.400 3096.700 2917.600 3153.180 ;
        RECT 2.800 3094.700 2917.600 3096.700 ;
        RECT 2.400 3088.540 2917.600 3094.700 ;
        RECT 2.400 3086.540 2917.200 3088.540 ;
        RECT 2.400 3031.420 2917.600 3086.540 ;
        RECT 2.800 3029.420 2917.600 3031.420 ;
        RECT 2.400 3021.900 2917.600 3029.420 ;
        RECT 2.400 3019.900 2917.200 3021.900 ;
        RECT 2.400 2966.140 2917.600 3019.900 ;
        RECT 2.800 2964.140 2917.600 2966.140 ;
        RECT 2.400 2955.940 2917.600 2964.140 ;
        RECT 2.400 2953.940 2917.200 2955.940 ;
        RECT 2.400 2900.860 2917.600 2953.940 ;
        RECT 2.800 2898.860 2917.600 2900.860 ;
        RECT 2.400 2889.300 2917.600 2898.860 ;
        RECT 2.400 2887.300 2917.200 2889.300 ;
        RECT 2.400 2835.580 2917.600 2887.300 ;
        RECT 2.800 2833.580 2917.600 2835.580 ;
        RECT 2.400 2822.660 2917.600 2833.580 ;
        RECT 2.400 2820.660 2917.200 2822.660 ;
        RECT 2.400 2770.300 2917.600 2820.660 ;
        RECT 2.800 2768.300 2917.600 2770.300 ;
        RECT 2.400 2756.700 2917.600 2768.300 ;
        RECT 2.400 2754.700 2917.200 2756.700 ;
        RECT 2.400 2705.020 2917.600 2754.700 ;
        RECT 2.800 2703.020 2917.600 2705.020 ;
        RECT 2.400 2690.060 2917.600 2703.020 ;
        RECT 2.400 2688.060 2917.200 2690.060 ;
        RECT 2.400 2640.420 2917.600 2688.060 ;
        RECT 2.800 2638.420 2917.600 2640.420 ;
        RECT 2.400 2623.420 2917.600 2638.420 ;
        RECT 2.400 2621.420 2917.200 2623.420 ;
        RECT 2.400 2575.140 2917.600 2621.420 ;
        RECT 2.800 2573.140 2917.600 2575.140 ;
        RECT 2.400 2557.460 2917.600 2573.140 ;
        RECT 2.400 2555.460 2917.200 2557.460 ;
        RECT 2.400 2509.860 2917.600 2555.460 ;
        RECT 2.800 2507.860 2917.600 2509.860 ;
        RECT 2.400 2490.820 2917.600 2507.860 ;
        RECT 2.400 2488.820 2917.200 2490.820 ;
        RECT 2.400 2444.580 2917.600 2488.820 ;
        RECT 2.800 2442.580 2917.600 2444.580 ;
        RECT 2.400 2424.180 2917.600 2442.580 ;
        RECT 2.400 2422.180 2917.200 2424.180 ;
        RECT 2.400 2379.300 2917.600 2422.180 ;
        RECT 2.800 2377.300 2917.600 2379.300 ;
        RECT 2.400 2358.220 2917.600 2377.300 ;
        RECT 2.400 2356.220 2917.200 2358.220 ;
        RECT 2.400 2314.020 2917.600 2356.220 ;
        RECT 2.800 2312.020 2917.600 2314.020 ;
        RECT 2.400 2291.580 2917.600 2312.020 ;
        RECT 2.400 2289.580 2917.200 2291.580 ;
        RECT 2.400 2248.740 2917.600 2289.580 ;
        RECT 2.800 2246.740 2917.600 2248.740 ;
        RECT 2.400 2224.940 2917.600 2246.740 ;
        RECT 2.400 2222.940 2917.200 2224.940 ;
        RECT 2.400 2184.140 2917.600 2222.940 ;
        RECT 2.800 2182.140 2917.600 2184.140 ;
        RECT 2.400 2158.980 2917.600 2182.140 ;
        RECT 2.400 2156.980 2917.200 2158.980 ;
        RECT 2.400 2118.860 2917.600 2156.980 ;
        RECT 2.800 2116.860 2917.600 2118.860 ;
        RECT 2.400 2092.340 2917.600 2116.860 ;
        RECT 2.400 2090.340 2917.200 2092.340 ;
        RECT 2.400 2053.580 2917.600 2090.340 ;
        RECT 2.800 2051.580 2917.600 2053.580 ;
        RECT 2.400 2025.700 2917.600 2051.580 ;
        RECT 2.400 2023.700 2917.200 2025.700 ;
        RECT 2.400 1988.300 2917.600 2023.700 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 2.400 1959.740 2917.600 1986.300 ;
        RECT 2.400 1957.740 2917.200 1959.740 ;
        RECT 2.400 1923.020 2917.600 1957.740 ;
        RECT 2.800 1921.020 2917.600 1923.020 ;
        RECT 2.400 1893.100 2917.600 1921.020 ;
        RECT 2.400 1891.100 2917.200 1893.100 ;
        RECT 2.400 1857.740 2917.600 1891.100 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 2.400 1826.460 2917.600 1855.740 ;
        RECT 2.400 1824.460 2917.200 1826.460 ;
        RECT 2.400 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 2.400 1760.500 2917.600 1791.140 ;
        RECT 2.400 1758.500 2917.200 1760.500 ;
        RECT 2.400 1727.860 2917.600 1758.500 ;
        RECT 2.800 1725.860 2917.600 1727.860 ;
        RECT 2.400 1693.860 2917.600 1725.860 ;
        RECT 2.400 1691.860 2917.200 1693.860 ;
        RECT 2.400 1662.580 2917.600 1691.860 ;
        RECT 2.800 1660.580 2917.600 1662.580 ;
        RECT 2.400 1627.220 2917.600 1660.580 ;
        RECT 2.400 1625.220 2917.200 1627.220 ;
        RECT 2.400 1597.300 2917.600 1625.220 ;
        RECT 2.800 1595.300 2917.600 1597.300 ;
        RECT 2.400 1561.260 2917.600 1595.300 ;
        RECT 2.400 1559.260 2917.200 1561.260 ;
        RECT 2.400 1532.020 2917.600 1559.260 ;
        RECT 2.800 1530.020 2917.600 1532.020 ;
        RECT 2.400 1494.620 2917.600 1530.020 ;
        RECT 2.400 1492.620 2917.200 1494.620 ;
        RECT 2.400 1466.740 2917.600 1492.620 ;
        RECT 2.800 1464.740 2917.600 1466.740 ;
        RECT 2.400 1427.980 2917.600 1464.740 ;
        RECT 2.400 1425.980 2917.200 1427.980 ;
        RECT 2.400 1401.460 2917.600 1425.980 ;
        RECT 2.800 1399.460 2917.600 1401.460 ;
        RECT 2.400 1362.020 2917.600 1399.460 ;
        RECT 2.400 1360.020 2917.200 1362.020 ;
        RECT 2.400 1336.860 2917.600 1360.020 ;
        RECT 2.800 1334.860 2917.600 1336.860 ;
        RECT 2.400 1295.380 2917.600 1334.860 ;
        RECT 2.400 1293.380 2917.200 1295.380 ;
        RECT 2.400 1271.580 2917.600 1293.380 ;
        RECT 2.800 1269.580 2917.600 1271.580 ;
        RECT 2.400 1228.740 2917.600 1269.580 ;
        RECT 2.400 1226.740 2917.200 1228.740 ;
        RECT 2.400 1206.300 2917.600 1226.740 ;
        RECT 2.800 1204.300 2917.600 1206.300 ;
        RECT 2.400 1162.780 2917.600 1204.300 ;
        RECT 2.400 1160.780 2917.200 1162.780 ;
        RECT 2.400 1141.020 2917.600 1160.780 ;
        RECT 2.800 1139.020 2917.600 1141.020 ;
        RECT 2.400 1096.140 2917.600 1139.020 ;
        RECT 2.400 1094.140 2917.200 1096.140 ;
        RECT 2.400 1075.740 2917.600 1094.140 ;
        RECT 2.800 1073.740 2917.600 1075.740 ;
        RECT 2.400 1029.500 2917.600 1073.740 ;
        RECT 2.400 1027.500 2917.200 1029.500 ;
        RECT 2.400 1010.460 2917.600 1027.500 ;
        RECT 2.800 1008.460 2917.600 1010.460 ;
        RECT 2.400 963.540 2917.600 1008.460 ;
        RECT 2.400 961.540 2917.200 963.540 ;
        RECT 2.400 945.180 2917.600 961.540 ;
        RECT 2.800 943.180 2917.600 945.180 ;
        RECT 2.400 896.900 2917.600 943.180 ;
        RECT 2.400 894.900 2917.200 896.900 ;
        RECT 2.400 880.580 2917.600 894.900 ;
        RECT 2.800 878.580 2917.600 880.580 ;
        RECT 2.400 830.260 2917.600 878.580 ;
        RECT 2.400 828.260 2917.200 830.260 ;
        RECT 2.400 815.300 2917.600 828.260 ;
        RECT 2.800 813.300 2917.600 815.300 ;
        RECT 2.400 764.300 2917.600 813.300 ;
        RECT 2.400 762.300 2917.200 764.300 ;
        RECT 2.400 750.020 2917.600 762.300 ;
        RECT 2.800 748.020 2917.600 750.020 ;
        RECT 2.400 697.660 2917.600 748.020 ;
        RECT 2.400 695.660 2917.200 697.660 ;
        RECT 2.400 684.740 2917.600 695.660 ;
        RECT 2.800 682.740 2917.600 684.740 ;
        RECT 2.400 631.020 2917.600 682.740 ;
        RECT 2.400 629.020 2917.200 631.020 ;
        RECT 2.400 619.460 2917.600 629.020 ;
        RECT 2.800 617.460 2917.600 619.460 ;
        RECT 2.400 565.060 2917.600 617.460 ;
        RECT 2.400 563.060 2917.200 565.060 ;
        RECT 2.400 554.180 2917.600 563.060 ;
        RECT 2.800 552.180 2917.600 554.180 ;
        RECT 2.400 498.420 2917.600 552.180 ;
        RECT 2.400 496.420 2917.200 498.420 ;
        RECT 2.400 488.900 2917.600 496.420 ;
        RECT 2.800 486.900 2917.600 488.900 ;
        RECT 2.400 431.780 2917.600 486.900 ;
        RECT 2.400 429.780 2917.200 431.780 ;
        RECT 2.400 424.300 2917.600 429.780 ;
        RECT 2.800 422.300 2917.600 424.300 ;
        RECT 2.400 365.820 2917.600 422.300 ;
        RECT 2.400 363.820 2917.200 365.820 ;
        RECT 2.400 359.020 2917.600 363.820 ;
        RECT 2.800 357.020 2917.600 359.020 ;
        RECT 2.400 299.180 2917.600 357.020 ;
        RECT 2.400 297.180 2917.200 299.180 ;
        RECT 2.400 293.740 2917.600 297.180 ;
        RECT 2.800 291.740 2917.600 293.740 ;
        RECT 2.400 232.540 2917.600 291.740 ;
        RECT 2.400 230.540 2917.200 232.540 ;
        RECT 2.400 228.460 2917.600 230.540 ;
        RECT 2.800 226.460 2917.600 228.460 ;
        RECT 2.400 166.580 2917.600 226.460 ;
        RECT 2.400 164.580 2917.200 166.580 ;
        RECT 2.400 163.180 2917.600 164.580 ;
        RECT 2.800 161.180 2917.600 163.180 ;
        RECT 2.400 99.940 2917.600 161.180 ;
        RECT 2.400 97.940 2917.200 99.940 ;
        RECT 2.400 97.900 2917.600 97.940 ;
        RECT 2.800 95.900 2917.600 97.900 ;
        RECT 2.400 33.980 2917.600 95.900 ;
        RECT 2.400 33.300 2917.200 33.980 ;
        RECT 2.800 31.980 2917.200 33.300 ;
        RECT 2.800 31.300 2917.600 31.980 ;
        RECT 2.400 10.715 2917.600 31.300 ;
      LAYER met4 ;
        RECT 150.620 2594.640 854.620 3278.105 ;
        RECT 150.620 2594.400 188.620 2594.640 ;
        RECT 150.620 13.095 152.620 2594.400 ;
        RECT 156.420 13.095 188.620 2594.400 ;
        RECT 192.420 2594.400 278.620 2594.640 ;
        RECT 192.420 13.095 206.620 2594.400 ;
        RECT 210.420 13.095 224.620 2594.400 ;
        RECT 228.420 13.095 242.620 2594.400 ;
        RECT 246.420 13.095 278.620 2594.400 ;
        RECT 282.420 2594.400 368.620 2594.640 ;
        RECT 282.420 13.095 296.620 2594.400 ;
        RECT 300.420 13.095 314.620 2594.400 ;
        RECT 318.420 13.095 332.620 2594.400 ;
        RECT 336.420 13.095 368.620 2594.400 ;
        RECT 372.420 2594.400 458.620 2594.640 ;
        RECT 372.420 13.095 386.620 2594.400 ;
        RECT 390.420 13.095 404.620 2594.400 ;
        RECT 408.420 13.095 422.620 2594.400 ;
        RECT 426.420 13.095 458.620 2594.400 ;
        RECT 462.420 2594.400 548.620 2594.640 ;
        RECT 462.420 13.095 476.620 2594.400 ;
        RECT 480.420 13.095 494.620 2594.400 ;
        RECT 498.420 13.095 512.620 2594.400 ;
        RECT 516.420 13.095 548.620 2594.400 ;
        RECT 552.420 2594.400 638.620 2594.640 ;
        RECT 552.420 13.095 566.620 2594.400 ;
        RECT 570.420 13.095 584.620 2594.400 ;
        RECT 588.420 13.095 602.620 2594.400 ;
        RECT 606.420 13.095 638.620 2594.400 ;
        RECT 642.420 2594.400 728.620 2594.640 ;
        RECT 642.420 13.095 656.620 2594.400 ;
        RECT 660.420 13.095 674.620 2594.400 ;
        RECT 678.420 13.095 692.620 2594.400 ;
        RECT 696.420 13.095 728.620 2594.400 ;
        RECT 732.420 2594.400 818.620 2594.640 ;
        RECT 732.420 13.095 746.620 2594.400 ;
        RECT 750.420 13.095 764.620 2594.400 ;
        RECT 768.420 13.095 782.620 2594.400 ;
        RECT 786.420 13.095 818.620 2594.400 ;
        RECT 822.420 2594.400 854.620 2594.640 ;
        RECT 822.420 13.095 836.620 2594.400 ;
        RECT 840.420 13.095 854.620 2594.400 ;
        RECT 858.420 13.095 872.620 3278.105 ;
        RECT 876.420 13.095 908.620 3278.105 ;
        RECT 912.420 13.095 926.620 3278.105 ;
        RECT 930.420 13.095 944.620 3278.105 ;
        RECT 948.420 13.095 962.620 3278.105 ;
        RECT 966.420 13.095 998.620 3278.105 ;
        RECT 1002.420 13.095 1016.620 3278.105 ;
        RECT 1020.420 13.095 1034.620 3278.105 ;
        RECT 1038.420 13.095 1052.620 3278.105 ;
        RECT 1056.420 13.095 1088.620 3278.105 ;
        RECT 1092.420 13.095 1106.620 3278.105 ;
        RECT 1110.420 13.095 1124.620 3278.105 ;
        RECT 1128.420 13.095 1142.620 3278.105 ;
        RECT 1146.420 2299.360 1178.620 3278.105 ;
        RECT 1182.420 2299.600 1196.620 3278.105 ;
        RECT 1200.420 2299.600 1214.620 3278.105 ;
        RECT 1218.420 2299.600 1232.620 3278.105 ;
        RECT 1236.420 2299.600 1268.620 3278.105 ;
        RECT 1182.420 2299.360 1268.620 2299.600 ;
        RECT 1272.420 2299.600 1286.620 3278.105 ;
        RECT 1290.420 2299.600 1304.620 3278.105 ;
        RECT 1308.420 2299.600 1322.620 3278.105 ;
        RECT 1326.420 2299.600 1358.620 3278.105 ;
        RECT 1272.420 2299.360 1358.620 2299.600 ;
        RECT 1362.420 2299.600 1376.620 3278.105 ;
        RECT 1380.420 2299.600 1394.620 3278.105 ;
        RECT 1398.420 2299.600 1412.620 3278.105 ;
        RECT 1416.420 2299.600 1448.620 3278.105 ;
        RECT 1362.420 2299.360 1448.620 2299.600 ;
        RECT 1452.420 2299.600 1466.620 3278.105 ;
        RECT 1470.420 2299.600 1484.620 3278.105 ;
        RECT 1488.420 2299.600 1502.620 3278.105 ;
        RECT 1506.420 2299.600 1538.620 3278.105 ;
        RECT 1452.420 2299.360 1538.620 2299.600 ;
        RECT 1542.420 2299.600 1556.620 3278.105 ;
        RECT 1560.420 2299.600 1574.620 3278.105 ;
        RECT 1578.420 2299.600 1592.620 3278.105 ;
        RECT 1596.420 2299.600 1628.620 3278.105 ;
        RECT 1542.420 2299.360 1628.620 2299.600 ;
        RECT 1632.420 2299.600 1646.620 3278.105 ;
        RECT 1650.420 2299.600 1664.620 3278.105 ;
        RECT 1668.420 2299.600 1682.620 3278.105 ;
        RECT 1686.420 2299.600 1718.620 3278.105 ;
        RECT 1632.420 2299.360 1718.620 2299.600 ;
        RECT 1722.420 2299.600 1736.620 3278.105 ;
        RECT 1740.420 2299.600 1754.620 3278.105 ;
        RECT 1758.420 2299.600 1772.620 3278.105 ;
        RECT 1776.420 2299.600 1808.620 3278.105 ;
        RECT 1722.420 2299.360 1808.620 2299.600 ;
        RECT 1812.420 2299.600 1826.620 3278.105 ;
        RECT 1830.420 2299.600 1844.620 3278.105 ;
        RECT 1848.420 2299.600 1862.620 3278.105 ;
        RECT 1866.420 2299.600 1898.620 3278.105 ;
        RECT 1812.420 2299.360 1898.620 2299.600 ;
        RECT 1902.420 2299.600 1916.620 3278.105 ;
        RECT 1920.420 2299.600 1934.620 3278.105 ;
        RECT 1938.420 2299.600 1952.620 3278.105 ;
        RECT 1956.420 2299.600 1988.620 3278.105 ;
        RECT 1902.420 2299.360 1988.620 2299.600 ;
        RECT 1992.420 2299.600 2006.620 3278.105 ;
        RECT 2010.420 2299.600 2024.620 3278.105 ;
        RECT 2028.420 2299.600 2042.620 3278.105 ;
        RECT 2046.420 2299.600 2078.620 3278.105 ;
        RECT 1992.420 2299.360 2078.620 2299.600 ;
        RECT 2082.420 2299.360 2096.620 3278.105 ;
        RECT 1146.420 1680.640 2096.620 2299.360 ;
        RECT 1146.420 13.095 1178.620 1680.640 ;
        RECT 1182.420 1680.400 1268.620 1680.640 ;
        RECT 1182.420 13.095 1196.620 1680.400 ;
        RECT 1200.420 13.095 1214.620 1680.400 ;
        RECT 1218.420 13.095 1232.620 1680.400 ;
        RECT 1236.420 13.095 1268.620 1680.400 ;
        RECT 1272.420 1680.400 1358.620 1680.640 ;
        RECT 1272.420 13.095 1286.620 1680.400 ;
        RECT 1290.420 13.095 1304.620 1680.400 ;
        RECT 1308.420 13.095 1322.620 1680.400 ;
        RECT 1326.420 13.095 1358.620 1680.400 ;
        RECT 1362.420 1680.400 1448.620 1680.640 ;
        RECT 1362.420 13.095 1376.620 1680.400 ;
        RECT 1380.420 13.095 1394.620 1680.400 ;
        RECT 1398.420 13.095 1412.620 1680.400 ;
        RECT 1416.420 13.095 1448.620 1680.400 ;
        RECT 1452.420 1680.400 1538.620 1680.640 ;
        RECT 1452.420 13.095 1466.620 1680.400 ;
        RECT 1470.420 13.095 1484.620 1680.400 ;
        RECT 1488.420 13.095 1502.620 1680.400 ;
        RECT 1506.420 13.095 1538.620 1680.400 ;
        RECT 1542.420 1680.400 1628.620 1680.640 ;
        RECT 1542.420 13.095 1556.620 1680.400 ;
        RECT 1560.420 13.095 1574.620 1680.400 ;
        RECT 1578.420 13.095 1592.620 1680.400 ;
        RECT 1596.420 13.095 1628.620 1680.400 ;
        RECT 1632.420 1680.400 1718.620 1680.640 ;
        RECT 1632.420 13.095 1646.620 1680.400 ;
        RECT 1650.420 13.095 1664.620 1680.400 ;
        RECT 1668.420 13.095 1682.620 1680.400 ;
        RECT 1686.420 13.095 1718.620 1680.400 ;
        RECT 1722.420 1680.400 1808.620 1680.640 ;
        RECT 1722.420 13.095 1736.620 1680.400 ;
        RECT 1740.420 13.095 1754.620 1680.400 ;
        RECT 1758.420 13.095 1772.620 1680.400 ;
        RECT 1776.420 13.095 1808.620 1680.400 ;
        RECT 1812.420 1680.400 1898.620 1680.640 ;
        RECT 1812.420 13.095 1826.620 1680.400 ;
        RECT 1830.420 13.095 1844.620 1680.400 ;
        RECT 1848.420 13.095 1862.620 1680.400 ;
        RECT 1866.420 13.095 1898.620 1680.400 ;
        RECT 1902.420 1680.400 1988.620 1680.640 ;
        RECT 1902.420 13.095 1916.620 1680.400 ;
        RECT 1920.420 13.095 1934.620 1680.400 ;
        RECT 1938.420 13.095 1952.620 1680.400 ;
        RECT 1956.420 13.095 1988.620 1680.400 ;
        RECT 1992.420 1680.400 2078.620 1680.640 ;
        RECT 1992.420 13.095 2006.620 1680.400 ;
        RECT 2010.420 13.095 2024.620 1680.400 ;
        RECT 2028.420 13.095 2042.620 1680.400 ;
        RECT 2046.420 13.095 2078.620 1680.400 ;
        RECT 2082.420 13.095 2096.620 1680.640 ;
        RECT 2100.420 13.095 2114.620 3278.105 ;
        RECT 2118.420 13.095 2132.620 3278.105 ;
        RECT 2136.420 13.095 2168.620 3278.105 ;
        RECT 2172.420 13.095 2186.620 3278.105 ;
        RECT 2190.420 13.095 2204.620 3278.105 ;
        RECT 2208.420 13.095 2222.620 3278.105 ;
        RECT 2226.420 13.095 2258.620 3278.105 ;
        RECT 2262.420 13.095 2276.620 3278.105 ;
        RECT 2280.420 13.095 2294.620 3278.105 ;
        RECT 2298.420 13.095 2312.620 3278.105 ;
        RECT 2316.420 13.095 2348.620 3278.105 ;
        RECT 2352.420 13.095 2366.620 3278.105 ;
        RECT 2370.420 13.095 2384.620 3278.105 ;
        RECT 2388.420 13.095 2402.620 3278.105 ;
        RECT 2406.420 13.095 2438.620 3278.105 ;
        RECT 2442.420 13.095 2456.620 3278.105 ;
        RECT 2460.420 13.095 2474.620 3278.105 ;
        RECT 2478.420 13.095 2492.620 3278.105 ;
        RECT 2496.420 2584.520 2528.620 3278.105 ;
        RECT 2532.420 2584.760 2546.620 3278.105 ;
        RECT 2550.420 2584.760 2564.620 3278.105 ;
        RECT 2568.420 2584.760 2582.620 3278.105 ;
        RECT 2586.420 2584.760 2618.620 3278.105 ;
        RECT 2532.420 2584.520 2618.620 2584.760 ;
        RECT 2622.420 2584.760 2636.620 3278.105 ;
        RECT 2640.420 2584.760 2654.620 3278.105 ;
        RECT 2658.420 2584.760 2672.620 3278.105 ;
        RECT 2676.420 2584.760 2692.490 3278.105 ;
        RECT 2622.420 2584.520 2692.490 2584.760 ;
        RECT 2496.420 2446.800 2692.490 2584.520 ;
        RECT 2496.420 2045.760 2528.620 2446.800 ;
        RECT 2532.420 2446.560 2618.620 2446.800 ;
        RECT 2532.420 2046.000 2546.620 2446.560 ;
        RECT 2550.420 2046.000 2564.620 2446.560 ;
        RECT 2568.420 2046.000 2582.620 2446.560 ;
        RECT 2586.420 2046.000 2618.620 2446.560 ;
        RECT 2532.420 2045.760 2618.620 2046.000 ;
        RECT 2622.420 2446.560 2692.490 2446.800 ;
        RECT 2622.420 2046.000 2636.620 2446.560 ;
        RECT 2640.420 2046.000 2654.620 2446.560 ;
        RECT 2658.420 2046.000 2672.620 2446.560 ;
        RECT 2676.420 2046.000 2692.490 2446.560 ;
        RECT 2622.420 2045.760 2692.490 2046.000 ;
        RECT 2496.420 1908.040 2692.490 2045.760 ;
        RECT 2496.420 1504.680 2528.620 1908.040 ;
        RECT 2532.420 1907.800 2618.620 1908.040 ;
        RECT 2532.420 1504.920 2546.620 1907.800 ;
        RECT 2550.420 1504.920 2564.620 1907.800 ;
        RECT 2568.420 1504.920 2582.620 1907.800 ;
        RECT 2586.420 1504.920 2618.620 1907.800 ;
        RECT 2532.420 1504.680 2618.620 1504.920 ;
        RECT 2622.420 1907.800 2692.490 1908.040 ;
        RECT 2622.420 1504.920 2636.620 1907.800 ;
        RECT 2640.420 1504.920 2654.620 1907.800 ;
        RECT 2658.420 1504.920 2672.620 1907.800 ;
        RECT 2676.420 1504.920 2692.490 1907.800 ;
        RECT 2622.420 1504.680 2692.490 1504.920 ;
        RECT 2496.420 1366.960 2692.490 1504.680 ;
        RECT 2496.420 13.095 2528.620 1366.960 ;
        RECT 2532.420 1366.720 2618.620 1366.960 ;
        RECT 2532.420 13.095 2546.620 1366.720 ;
        RECT 2550.420 13.095 2564.620 1366.720 ;
        RECT 2568.420 13.095 2582.620 1366.720 ;
        RECT 2586.420 13.095 2618.620 1366.720 ;
        RECT 2622.420 1366.720 2692.490 1366.960 ;
        RECT 2622.420 13.095 2636.620 1366.720 ;
        RECT 2640.420 13.095 2654.620 1366.720 ;
        RECT 2658.420 13.095 2672.620 1366.720 ;
        RECT 2676.420 13.095 2692.490 1366.720 ;
      LAYER met5 ;
        RECT -42.880 3557.200 -39.880 3557.210 ;
        RECT 153.020 3557.200 156.020 3557.210 ;
        RECT 333.020 3557.200 336.020 3557.210 ;
        RECT 513.020 3557.200 516.020 3557.210 ;
        RECT 693.020 3557.200 696.020 3557.210 ;
        RECT 873.020 3557.200 876.020 3557.210 ;
        RECT 1053.020 3557.200 1056.020 3557.210 ;
        RECT 1233.020 3557.200 1236.020 3557.210 ;
        RECT 1413.020 3557.200 1416.020 3557.210 ;
        RECT 1593.020 3557.200 1596.020 3557.210 ;
        RECT 1773.020 3557.200 1776.020 3557.210 ;
        RECT 1953.020 3557.200 1956.020 3557.210 ;
        RECT 2133.020 3557.200 2136.020 3557.210 ;
        RECT 2313.020 3557.200 2316.020 3557.210 ;
        RECT 2493.020 3557.200 2496.020 3557.210 ;
        RECT 2673.020 3557.200 2676.020 3557.210 ;
        RECT 2853.020 3557.200 2856.020 3557.210 ;
        RECT 2959.500 3557.200 2962.500 3557.210 ;
        RECT -42.880 3554.190 -39.880 3554.200 ;
        RECT 153.020 3554.190 156.020 3554.200 ;
        RECT 333.020 3554.190 336.020 3554.200 ;
        RECT 513.020 3554.190 516.020 3554.200 ;
        RECT 693.020 3554.190 696.020 3554.200 ;
        RECT 873.020 3554.190 876.020 3554.200 ;
        RECT 1053.020 3554.190 1056.020 3554.200 ;
        RECT 1233.020 3554.190 1236.020 3554.200 ;
        RECT 1413.020 3554.190 1416.020 3554.200 ;
        RECT 1593.020 3554.190 1596.020 3554.200 ;
        RECT 1773.020 3554.190 1776.020 3554.200 ;
        RECT 1953.020 3554.190 1956.020 3554.200 ;
        RECT 2133.020 3554.190 2136.020 3554.200 ;
        RECT 2313.020 3554.190 2316.020 3554.200 ;
        RECT 2493.020 3554.190 2496.020 3554.200 ;
        RECT 2673.020 3554.190 2676.020 3554.200 ;
        RECT 2853.020 3554.190 2856.020 3554.200 ;
        RECT 2959.500 3554.190 2962.500 3554.200 ;
        RECT -38.180 3552.500 -35.180 3552.510 ;
        RECT 63.020 3552.500 66.020 3552.510 ;
        RECT 243.020 3552.500 246.020 3552.510 ;
        RECT 423.020 3552.500 426.020 3552.510 ;
        RECT 603.020 3552.500 606.020 3552.510 ;
        RECT 783.020 3552.500 786.020 3552.510 ;
        RECT 963.020 3552.500 966.020 3552.510 ;
        RECT 1143.020 3552.500 1146.020 3552.510 ;
        RECT 1323.020 3552.500 1326.020 3552.510 ;
        RECT 1503.020 3552.500 1506.020 3552.510 ;
        RECT 1683.020 3552.500 1686.020 3552.510 ;
        RECT 1863.020 3552.500 1866.020 3552.510 ;
        RECT 2043.020 3552.500 2046.020 3552.510 ;
        RECT 2223.020 3552.500 2226.020 3552.510 ;
        RECT 2403.020 3552.500 2406.020 3552.510 ;
        RECT 2583.020 3552.500 2586.020 3552.510 ;
        RECT 2763.020 3552.500 2766.020 3552.510 ;
        RECT 2954.800 3552.500 2957.800 3552.510 ;
        RECT -38.180 3549.490 -35.180 3549.500 ;
        RECT 63.020 3549.490 66.020 3549.500 ;
        RECT 243.020 3549.490 246.020 3549.500 ;
        RECT 423.020 3549.490 426.020 3549.500 ;
        RECT 603.020 3549.490 606.020 3549.500 ;
        RECT 783.020 3549.490 786.020 3549.500 ;
        RECT 963.020 3549.490 966.020 3549.500 ;
        RECT 1143.020 3549.490 1146.020 3549.500 ;
        RECT 1323.020 3549.490 1326.020 3549.500 ;
        RECT 1503.020 3549.490 1506.020 3549.500 ;
        RECT 1683.020 3549.490 1686.020 3549.500 ;
        RECT 1863.020 3549.490 1866.020 3549.500 ;
        RECT 2043.020 3549.490 2046.020 3549.500 ;
        RECT 2223.020 3549.490 2226.020 3549.500 ;
        RECT 2403.020 3549.490 2406.020 3549.500 ;
        RECT 2583.020 3549.490 2586.020 3549.500 ;
        RECT 2763.020 3549.490 2766.020 3549.500 ;
        RECT 2954.800 3549.490 2957.800 3549.500 ;
        RECT -33.480 3547.800 -30.480 3547.810 ;
        RECT 135.020 3547.800 138.020 3547.810 ;
        RECT 315.020 3547.800 318.020 3547.810 ;
        RECT 495.020 3547.800 498.020 3547.810 ;
        RECT 675.020 3547.800 678.020 3547.810 ;
        RECT 855.020 3547.800 858.020 3547.810 ;
        RECT 1035.020 3547.800 1038.020 3547.810 ;
        RECT 1215.020 3547.800 1218.020 3547.810 ;
        RECT 1395.020 3547.800 1398.020 3547.810 ;
        RECT 1575.020 3547.800 1578.020 3547.810 ;
        RECT 1755.020 3547.800 1758.020 3547.810 ;
        RECT 1935.020 3547.800 1938.020 3547.810 ;
        RECT 2115.020 3547.800 2118.020 3547.810 ;
        RECT 2295.020 3547.800 2298.020 3547.810 ;
        RECT 2475.020 3547.800 2478.020 3547.810 ;
        RECT 2655.020 3547.800 2658.020 3547.810 ;
        RECT 2835.020 3547.800 2838.020 3547.810 ;
        RECT 2950.100 3547.800 2953.100 3547.810 ;
        RECT -33.480 3544.790 -30.480 3544.800 ;
        RECT 135.020 3544.790 138.020 3544.800 ;
        RECT 315.020 3544.790 318.020 3544.800 ;
        RECT 495.020 3544.790 498.020 3544.800 ;
        RECT 675.020 3544.790 678.020 3544.800 ;
        RECT 855.020 3544.790 858.020 3544.800 ;
        RECT 1035.020 3544.790 1038.020 3544.800 ;
        RECT 1215.020 3544.790 1218.020 3544.800 ;
        RECT 1395.020 3544.790 1398.020 3544.800 ;
        RECT 1575.020 3544.790 1578.020 3544.800 ;
        RECT 1755.020 3544.790 1758.020 3544.800 ;
        RECT 1935.020 3544.790 1938.020 3544.800 ;
        RECT 2115.020 3544.790 2118.020 3544.800 ;
        RECT 2295.020 3544.790 2298.020 3544.800 ;
        RECT 2475.020 3544.790 2478.020 3544.800 ;
        RECT 2655.020 3544.790 2658.020 3544.800 ;
        RECT 2835.020 3544.790 2838.020 3544.800 ;
        RECT 2950.100 3544.790 2953.100 3544.800 ;
        RECT -28.780 3543.100 -25.780 3543.110 ;
        RECT 45.020 3543.100 48.020 3543.110 ;
        RECT 225.020 3543.100 228.020 3543.110 ;
        RECT 405.020 3543.100 408.020 3543.110 ;
        RECT 585.020 3543.100 588.020 3543.110 ;
        RECT 765.020 3543.100 768.020 3543.110 ;
        RECT 945.020 3543.100 948.020 3543.110 ;
        RECT 1125.020 3543.100 1128.020 3543.110 ;
        RECT 1305.020 3543.100 1308.020 3543.110 ;
        RECT 1485.020 3543.100 1488.020 3543.110 ;
        RECT 1665.020 3543.100 1668.020 3543.110 ;
        RECT 1845.020 3543.100 1848.020 3543.110 ;
        RECT 2025.020 3543.100 2028.020 3543.110 ;
        RECT 2205.020 3543.100 2208.020 3543.110 ;
        RECT 2385.020 3543.100 2388.020 3543.110 ;
        RECT 2565.020 3543.100 2568.020 3543.110 ;
        RECT 2745.020 3543.100 2748.020 3543.110 ;
        RECT 2945.400 3543.100 2948.400 3543.110 ;
        RECT -28.780 3540.090 -25.780 3540.100 ;
        RECT 45.020 3540.090 48.020 3540.100 ;
        RECT 225.020 3540.090 228.020 3540.100 ;
        RECT 405.020 3540.090 408.020 3540.100 ;
        RECT 585.020 3540.090 588.020 3540.100 ;
        RECT 765.020 3540.090 768.020 3540.100 ;
        RECT 945.020 3540.090 948.020 3540.100 ;
        RECT 1125.020 3540.090 1128.020 3540.100 ;
        RECT 1305.020 3540.090 1308.020 3540.100 ;
        RECT 1485.020 3540.090 1488.020 3540.100 ;
        RECT 1665.020 3540.090 1668.020 3540.100 ;
        RECT 1845.020 3540.090 1848.020 3540.100 ;
        RECT 2025.020 3540.090 2028.020 3540.100 ;
        RECT 2205.020 3540.090 2208.020 3540.100 ;
        RECT 2385.020 3540.090 2388.020 3540.100 ;
        RECT 2565.020 3540.090 2568.020 3540.100 ;
        RECT 2745.020 3540.090 2748.020 3540.100 ;
        RECT 2945.400 3540.090 2948.400 3540.100 ;
        RECT -24.080 3538.400 -21.080 3538.410 ;
        RECT 117.020 3538.400 120.020 3538.410 ;
        RECT 297.020 3538.400 300.020 3538.410 ;
        RECT 477.020 3538.400 480.020 3538.410 ;
        RECT 657.020 3538.400 660.020 3538.410 ;
        RECT 837.020 3538.400 840.020 3538.410 ;
        RECT 1017.020 3538.400 1020.020 3538.410 ;
        RECT 1197.020 3538.400 1200.020 3538.410 ;
        RECT 1377.020 3538.400 1380.020 3538.410 ;
        RECT 1557.020 3538.400 1560.020 3538.410 ;
        RECT 1737.020 3538.400 1740.020 3538.410 ;
        RECT 1917.020 3538.400 1920.020 3538.410 ;
        RECT 2097.020 3538.400 2100.020 3538.410 ;
        RECT 2277.020 3538.400 2280.020 3538.410 ;
        RECT 2457.020 3538.400 2460.020 3538.410 ;
        RECT 2637.020 3538.400 2640.020 3538.410 ;
        RECT 2817.020 3538.400 2820.020 3538.410 ;
        RECT 2940.700 3538.400 2943.700 3538.410 ;
        RECT -24.080 3535.390 -21.080 3535.400 ;
        RECT 117.020 3535.390 120.020 3535.400 ;
        RECT 297.020 3535.390 300.020 3535.400 ;
        RECT 477.020 3535.390 480.020 3535.400 ;
        RECT 657.020 3535.390 660.020 3535.400 ;
        RECT 837.020 3535.390 840.020 3535.400 ;
        RECT 1017.020 3535.390 1020.020 3535.400 ;
        RECT 1197.020 3535.390 1200.020 3535.400 ;
        RECT 1377.020 3535.390 1380.020 3535.400 ;
        RECT 1557.020 3535.390 1560.020 3535.400 ;
        RECT 1737.020 3535.390 1740.020 3535.400 ;
        RECT 1917.020 3535.390 1920.020 3535.400 ;
        RECT 2097.020 3535.390 2100.020 3535.400 ;
        RECT 2277.020 3535.390 2280.020 3535.400 ;
        RECT 2457.020 3535.390 2460.020 3535.400 ;
        RECT 2637.020 3535.390 2640.020 3535.400 ;
        RECT 2817.020 3535.390 2820.020 3535.400 ;
        RECT 2940.700 3535.390 2943.700 3535.400 ;
        RECT -19.380 3533.700 -16.380 3533.710 ;
        RECT 27.020 3533.700 30.020 3533.710 ;
        RECT 207.020 3533.700 210.020 3533.710 ;
        RECT 387.020 3533.700 390.020 3533.710 ;
        RECT 567.020 3533.700 570.020 3533.710 ;
        RECT 747.020 3533.700 750.020 3533.710 ;
        RECT 927.020 3533.700 930.020 3533.710 ;
        RECT 1107.020 3533.700 1110.020 3533.710 ;
        RECT 1287.020 3533.700 1290.020 3533.710 ;
        RECT 1467.020 3533.700 1470.020 3533.710 ;
        RECT 1647.020 3533.700 1650.020 3533.710 ;
        RECT 1827.020 3533.700 1830.020 3533.710 ;
        RECT 2007.020 3533.700 2010.020 3533.710 ;
        RECT 2187.020 3533.700 2190.020 3533.710 ;
        RECT 2367.020 3533.700 2370.020 3533.710 ;
        RECT 2547.020 3533.700 2550.020 3533.710 ;
        RECT 2727.020 3533.700 2730.020 3533.710 ;
        RECT 2907.020 3533.700 2910.020 3533.710 ;
        RECT 2936.000 3533.700 2939.000 3533.710 ;
        RECT -19.380 3530.690 -16.380 3530.700 ;
        RECT 27.020 3530.690 30.020 3530.700 ;
        RECT 207.020 3530.690 210.020 3530.700 ;
        RECT 387.020 3530.690 390.020 3530.700 ;
        RECT 567.020 3530.690 570.020 3530.700 ;
        RECT 747.020 3530.690 750.020 3530.700 ;
        RECT 927.020 3530.690 930.020 3530.700 ;
        RECT 1107.020 3530.690 1110.020 3530.700 ;
        RECT 1287.020 3530.690 1290.020 3530.700 ;
        RECT 1467.020 3530.690 1470.020 3530.700 ;
        RECT 1647.020 3530.690 1650.020 3530.700 ;
        RECT 1827.020 3530.690 1830.020 3530.700 ;
        RECT 2007.020 3530.690 2010.020 3530.700 ;
        RECT 2187.020 3530.690 2190.020 3530.700 ;
        RECT 2367.020 3530.690 2370.020 3530.700 ;
        RECT 2547.020 3530.690 2550.020 3530.700 ;
        RECT 2727.020 3530.690 2730.020 3530.700 ;
        RECT 2907.020 3530.690 2910.020 3530.700 ;
        RECT 2936.000 3530.690 2939.000 3530.700 ;
        RECT -14.680 3529.000 -11.680 3529.010 ;
        RECT 99.020 3529.000 102.020 3529.010 ;
        RECT 279.020 3529.000 282.020 3529.010 ;
        RECT 459.020 3529.000 462.020 3529.010 ;
        RECT 639.020 3529.000 642.020 3529.010 ;
        RECT 819.020 3529.000 822.020 3529.010 ;
        RECT 999.020 3529.000 1002.020 3529.010 ;
        RECT 1179.020 3529.000 1182.020 3529.010 ;
        RECT 1359.020 3529.000 1362.020 3529.010 ;
        RECT 1539.020 3529.000 1542.020 3529.010 ;
        RECT 1719.020 3529.000 1722.020 3529.010 ;
        RECT 1899.020 3529.000 1902.020 3529.010 ;
        RECT 2079.020 3529.000 2082.020 3529.010 ;
        RECT 2259.020 3529.000 2262.020 3529.010 ;
        RECT 2439.020 3529.000 2442.020 3529.010 ;
        RECT 2619.020 3529.000 2622.020 3529.010 ;
        RECT 2799.020 3529.000 2802.020 3529.010 ;
        RECT 2931.300 3529.000 2934.300 3529.010 ;
        RECT -14.680 3525.990 -11.680 3526.000 ;
        RECT 99.020 3525.990 102.020 3526.000 ;
        RECT 279.020 3525.990 282.020 3526.000 ;
        RECT 459.020 3525.990 462.020 3526.000 ;
        RECT 639.020 3525.990 642.020 3526.000 ;
        RECT 819.020 3525.990 822.020 3526.000 ;
        RECT 999.020 3525.990 1002.020 3526.000 ;
        RECT 1179.020 3525.990 1182.020 3526.000 ;
        RECT 1359.020 3525.990 1362.020 3526.000 ;
        RECT 1539.020 3525.990 1542.020 3526.000 ;
        RECT 1719.020 3525.990 1722.020 3526.000 ;
        RECT 1899.020 3525.990 1902.020 3526.000 ;
        RECT 2079.020 3525.990 2082.020 3526.000 ;
        RECT 2259.020 3525.990 2262.020 3526.000 ;
        RECT 2439.020 3525.990 2442.020 3526.000 ;
        RECT 2619.020 3525.990 2622.020 3526.000 ;
        RECT 2799.020 3525.990 2802.020 3526.000 ;
        RECT 2931.300 3525.990 2934.300 3526.000 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 9.020 3524.300 12.020 3524.310 ;
        RECT 189.020 3524.300 192.020 3524.310 ;
        RECT 369.020 3524.300 372.020 3524.310 ;
        RECT 549.020 3524.300 552.020 3524.310 ;
        RECT 729.020 3524.300 732.020 3524.310 ;
        RECT 909.020 3524.300 912.020 3524.310 ;
        RECT 1089.020 3524.300 1092.020 3524.310 ;
        RECT 1269.020 3524.300 1272.020 3524.310 ;
        RECT 1449.020 3524.300 1452.020 3524.310 ;
        RECT 1629.020 3524.300 1632.020 3524.310 ;
        RECT 1809.020 3524.300 1812.020 3524.310 ;
        RECT 1989.020 3524.300 1992.020 3524.310 ;
        RECT 2169.020 3524.300 2172.020 3524.310 ;
        RECT 2349.020 3524.300 2352.020 3524.310 ;
        RECT 2529.020 3524.300 2532.020 3524.310 ;
        RECT 2709.020 3524.300 2712.020 3524.310 ;
        RECT 2889.020 3524.300 2892.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 9.020 3521.290 12.020 3521.300 ;
        RECT 189.020 3521.290 192.020 3521.300 ;
        RECT 369.020 3521.290 372.020 3521.300 ;
        RECT 549.020 3521.290 552.020 3521.300 ;
        RECT 729.020 3521.290 732.020 3521.300 ;
        RECT 909.020 3521.290 912.020 3521.300 ;
        RECT 1089.020 3521.290 1092.020 3521.300 ;
        RECT 1269.020 3521.290 1272.020 3521.300 ;
        RECT 1449.020 3521.290 1452.020 3521.300 ;
        RECT 1629.020 3521.290 1632.020 3521.300 ;
        RECT 1809.020 3521.290 1812.020 3521.300 ;
        RECT 1989.020 3521.290 1992.020 3521.300 ;
        RECT 2169.020 3521.290 2172.020 3521.300 ;
        RECT 2349.020 3521.290 2352.020 3521.300 ;
        RECT 2529.020 3521.290 2532.020 3521.300 ;
        RECT 2709.020 3521.290 2712.020 3521.300 ;
        RECT 2889.020 3521.290 2892.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT 0.000 3492.980 2920.000 3519.700 ;
        RECT -38.180 3491.380 -35.180 3491.390 ;
        RECT 2954.800 3491.380 2957.800 3491.390 ;
        RECT -38.180 3488.370 -35.180 3488.380 ;
        RECT 2954.800 3488.370 2957.800 3488.380 ;
        RECT 0.000 3474.980 2920.000 3486.780 ;
        RECT -28.780 3473.380 -25.780 3473.390 ;
        RECT 2945.400 3473.380 2948.400 3473.390 ;
        RECT -28.780 3470.370 -25.780 3470.380 ;
        RECT 2945.400 3470.370 2948.400 3470.380 ;
        RECT 0.000 3456.980 2920.000 3468.780 ;
        RECT -19.380 3455.380 -16.380 3455.390 ;
        RECT 2936.000 3455.380 2939.000 3455.390 ;
        RECT -19.380 3452.370 -16.380 3452.380 ;
        RECT 2936.000 3452.370 2939.000 3452.380 ;
        RECT 0.000 3438.740 2920.000 3450.780 ;
        RECT -9.980 3437.140 -6.980 3437.150 ;
        RECT 2926.600 3437.140 2929.600 3437.150 ;
        RECT -9.980 3434.130 -6.980 3434.140 ;
        RECT 2926.600 3434.130 2929.600 3434.140 ;
        RECT 0.000 3402.980 2920.000 3432.540 ;
        RECT -42.880 3401.380 -39.880 3401.390 ;
        RECT 2959.500 3401.380 2962.500 3401.390 ;
        RECT -42.880 3398.370 -39.880 3398.380 ;
        RECT 2959.500 3398.370 2962.500 3398.380 ;
        RECT 0.000 3384.980 2920.000 3396.780 ;
        RECT -33.480 3383.380 -30.480 3383.390 ;
        RECT 2950.100 3383.380 2953.100 3383.390 ;
        RECT -33.480 3380.370 -30.480 3380.380 ;
        RECT 2950.100 3380.370 2953.100 3380.380 ;
        RECT 0.000 3366.980 2920.000 3378.780 ;
        RECT -24.080 3365.380 -21.080 3365.390 ;
        RECT 2940.700 3365.380 2943.700 3365.390 ;
        RECT -24.080 3362.370 -21.080 3362.380 ;
        RECT 2940.700 3362.370 2943.700 3362.380 ;
        RECT 0.000 3348.740 2920.000 3360.780 ;
        RECT -14.680 3347.140 -11.680 3347.150 ;
        RECT 2931.300 3347.140 2934.300 3347.150 ;
        RECT -14.680 3344.130 -11.680 3344.140 ;
        RECT 2931.300 3344.130 2934.300 3344.140 ;
        RECT 0.000 3312.980 2920.000 3342.540 ;
        RECT -38.180 3311.380 -35.180 3311.390 ;
        RECT 2954.800 3311.380 2957.800 3311.390 ;
        RECT -38.180 3308.370 -35.180 3308.380 ;
        RECT 2954.800 3308.370 2957.800 3308.380 ;
        RECT 0.000 3294.980 2920.000 3306.780 ;
        RECT -28.780 3293.380 -25.780 3293.390 ;
        RECT 2945.400 3293.380 2948.400 3293.390 ;
        RECT -28.780 3290.370 -25.780 3290.380 ;
        RECT 2945.400 3290.370 2948.400 3290.380 ;
        RECT 0.000 3276.980 2920.000 3288.780 ;
        RECT -19.380 3275.380 -16.380 3275.390 ;
        RECT 2936.000 3275.380 2939.000 3275.390 ;
        RECT -19.380 3272.370 -16.380 3272.380 ;
        RECT 2936.000 3272.370 2939.000 3272.380 ;
        RECT 0.000 3258.740 2920.000 3270.780 ;
        RECT -9.980 3257.140 -6.980 3257.150 ;
        RECT 2926.600 3257.140 2929.600 3257.150 ;
        RECT -9.980 3254.130 -6.980 3254.140 ;
        RECT 2926.600 3254.130 2929.600 3254.140 ;
        RECT 0.000 3222.980 2920.000 3252.540 ;
        RECT -42.880 3221.380 -39.880 3221.390 ;
        RECT 2959.500 3221.380 2962.500 3221.390 ;
        RECT -42.880 3218.370 -39.880 3218.380 ;
        RECT 2959.500 3218.370 2962.500 3218.380 ;
        RECT 0.000 3204.980 2920.000 3216.780 ;
        RECT -33.480 3203.380 -30.480 3203.390 ;
        RECT 2950.100 3203.380 2953.100 3203.390 ;
        RECT -33.480 3200.370 -30.480 3200.380 ;
        RECT 2950.100 3200.370 2953.100 3200.380 ;
        RECT 0.000 3186.980 2920.000 3198.780 ;
        RECT -24.080 3185.380 -21.080 3185.390 ;
        RECT 2940.700 3185.380 2943.700 3185.390 ;
        RECT -24.080 3182.370 -21.080 3182.380 ;
        RECT 2940.700 3182.370 2943.700 3182.380 ;
        RECT 0.000 3168.740 2920.000 3180.780 ;
        RECT -14.680 3167.140 -11.680 3167.150 ;
        RECT 2931.300 3167.140 2934.300 3167.150 ;
        RECT -14.680 3164.130 -11.680 3164.140 ;
        RECT 2931.300 3164.130 2934.300 3164.140 ;
        RECT 0.000 3132.980 2920.000 3162.540 ;
        RECT -38.180 3131.380 -35.180 3131.390 ;
        RECT 2954.800 3131.380 2957.800 3131.390 ;
        RECT -38.180 3128.370 -35.180 3128.380 ;
        RECT 2954.800 3128.370 2957.800 3128.380 ;
        RECT 0.000 3114.980 2920.000 3126.780 ;
        RECT -28.780 3113.380 -25.780 3113.390 ;
        RECT 2945.400 3113.380 2948.400 3113.390 ;
        RECT -28.780 3110.370 -25.780 3110.380 ;
        RECT 2945.400 3110.370 2948.400 3110.380 ;
        RECT 0.000 3096.980 2920.000 3108.780 ;
        RECT -19.380 3095.380 -16.380 3095.390 ;
        RECT 2936.000 3095.380 2939.000 3095.390 ;
        RECT -19.380 3092.370 -16.380 3092.380 ;
        RECT 2936.000 3092.370 2939.000 3092.380 ;
        RECT 0.000 3078.740 2920.000 3090.780 ;
        RECT -9.980 3077.140 -6.980 3077.150 ;
        RECT 2926.600 3077.140 2929.600 3077.150 ;
        RECT -9.980 3074.130 -6.980 3074.140 ;
        RECT 2926.600 3074.130 2929.600 3074.140 ;
        RECT 0.000 3042.980 2920.000 3072.540 ;
        RECT -42.880 3041.380 -39.880 3041.390 ;
        RECT 2959.500 3041.380 2962.500 3041.390 ;
        RECT -42.880 3038.370 -39.880 3038.380 ;
        RECT 2959.500 3038.370 2962.500 3038.380 ;
        RECT 0.000 3024.980 2920.000 3036.780 ;
        RECT -33.480 3023.380 -30.480 3023.390 ;
        RECT 2950.100 3023.380 2953.100 3023.390 ;
        RECT -33.480 3020.370 -30.480 3020.380 ;
        RECT 2950.100 3020.370 2953.100 3020.380 ;
        RECT 0.000 3006.980 2920.000 3018.780 ;
        RECT -24.080 3005.380 -21.080 3005.390 ;
        RECT 2940.700 3005.380 2943.700 3005.390 ;
        RECT -24.080 3002.370 -21.080 3002.380 ;
        RECT 2940.700 3002.370 2943.700 3002.380 ;
        RECT 0.000 2988.740 2920.000 3000.780 ;
        RECT -14.680 2987.140 -11.680 2987.150 ;
        RECT 2931.300 2987.140 2934.300 2987.150 ;
        RECT -14.680 2984.130 -11.680 2984.140 ;
        RECT 2931.300 2984.130 2934.300 2984.140 ;
        RECT 0.000 2952.980 2920.000 2982.540 ;
        RECT -38.180 2951.380 -35.180 2951.390 ;
        RECT 2954.800 2951.380 2957.800 2951.390 ;
        RECT -38.180 2948.370 -35.180 2948.380 ;
        RECT 2954.800 2948.370 2957.800 2948.380 ;
        RECT 0.000 2934.980 2920.000 2946.780 ;
        RECT -28.780 2933.380 -25.780 2933.390 ;
        RECT 2945.400 2933.380 2948.400 2933.390 ;
        RECT -28.780 2930.370 -25.780 2930.380 ;
        RECT 2945.400 2930.370 2948.400 2930.380 ;
        RECT 0.000 2916.980 2920.000 2928.780 ;
        RECT -19.380 2915.380 -16.380 2915.390 ;
        RECT 2936.000 2915.380 2939.000 2915.390 ;
        RECT -19.380 2912.370 -16.380 2912.380 ;
        RECT 2936.000 2912.370 2939.000 2912.380 ;
        RECT 0.000 2898.740 2920.000 2910.780 ;
        RECT -9.980 2897.140 -6.980 2897.150 ;
        RECT 2926.600 2897.140 2929.600 2897.150 ;
        RECT -9.980 2894.130 -6.980 2894.140 ;
        RECT 2926.600 2894.130 2929.600 2894.140 ;
        RECT 0.000 2862.980 2920.000 2892.540 ;
        RECT -42.880 2861.380 -39.880 2861.390 ;
        RECT 2959.500 2861.380 2962.500 2861.390 ;
        RECT -42.880 2858.370 -39.880 2858.380 ;
        RECT 2959.500 2858.370 2962.500 2858.380 ;
        RECT 0.000 2844.980 2920.000 2856.780 ;
        RECT -33.480 2843.380 -30.480 2843.390 ;
        RECT 2950.100 2843.380 2953.100 2843.390 ;
        RECT -33.480 2840.370 -30.480 2840.380 ;
        RECT 2950.100 2840.370 2953.100 2840.380 ;
        RECT 0.000 2826.980 2920.000 2838.780 ;
        RECT -24.080 2825.380 -21.080 2825.390 ;
        RECT 2940.700 2825.380 2943.700 2825.390 ;
        RECT -24.080 2822.370 -21.080 2822.380 ;
        RECT 2940.700 2822.370 2943.700 2822.380 ;
        RECT 0.000 2808.740 2920.000 2820.780 ;
        RECT -14.680 2807.140 -11.680 2807.150 ;
        RECT 2931.300 2807.140 2934.300 2807.150 ;
        RECT -14.680 2804.130 -11.680 2804.140 ;
        RECT 2931.300 2804.130 2934.300 2804.140 ;
        RECT 0.000 2772.980 2920.000 2802.540 ;
        RECT -38.180 2771.380 -35.180 2771.390 ;
        RECT 2954.800 2771.380 2957.800 2771.390 ;
        RECT -38.180 2768.370 -35.180 2768.380 ;
        RECT 2954.800 2768.370 2957.800 2768.380 ;
        RECT 0.000 2754.980 2920.000 2766.780 ;
        RECT -28.780 2753.380 -25.780 2753.390 ;
        RECT 2945.400 2753.380 2948.400 2753.390 ;
        RECT -28.780 2750.370 -25.780 2750.380 ;
        RECT 2945.400 2750.370 2948.400 2750.380 ;
        RECT 0.000 2736.980 2920.000 2748.780 ;
        RECT -19.380 2735.380 -16.380 2735.390 ;
        RECT 2936.000 2735.380 2939.000 2735.390 ;
        RECT -19.380 2732.370 -16.380 2732.380 ;
        RECT 2936.000 2732.370 2939.000 2732.380 ;
        RECT 0.000 2718.740 2920.000 2730.780 ;
        RECT -9.980 2717.140 -6.980 2717.150 ;
        RECT 2926.600 2717.140 2929.600 2717.150 ;
        RECT -9.980 2714.130 -6.980 2714.140 ;
        RECT 2926.600 2714.130 2929.600 2714.140 ;
        RECT 0.000 2682.980 2920.000 2712.540 ;
        RECT -42.880 2681.380 -39.880 2681.390 ;
        RECT 2959.500 2681.380 2962.500 2681.390 ;
        RECT -42.880 2678.370 -39.880 2678.380 ;
        RECT 2959.500 2678.370 2962.500 2678.380 ;
        RECT 0.000 2664.980 2920.000 2676.780 ;
        RECT -33.480 2663.380 -30.480 2663.390 ;
        RECT 2950.100 2663.380 2953.100 2663.390 ;
        RECT -33.480 2660.370 -30.480 2660.380 ;
        RECT 2950.100 2660.370 2953.100 2660.380 ;
        RECT 0.000 2646.980 2920.000 2658.780 ;
        RECT -24.080 2645.380 -21.080 2645.390 ;
        RECT 2940.700 2645.380 2943.700 2645.390 ;
        RECT -24.080 2642.370 -21.080 2642.380 ;
        RECT 2940.700 2642.370 2943.700 2642.380 ;
        RECT 0.000 2628.740 2920.000 2640.780 ;
        RECT -14.680 2627.140 -11.680 2627.150 ;
        RECT 2931.300 2627.140 2934.300 2627.150 ;
        RECT -14.680 2624.130 -11.680 2624.140 ;
        RECT 2931.300 2624.130 2934.300 2624.140 ;
        RECT 0.000 2592.980 2920.000 2622.540 ;
        RECT -38.180 2591.380 -35.180 2591.390 ;
        RECT 2954.800 2591.380 2957.800 2591.390 ;
        RECT -38.180 2588.370 -35.180 2588.380 ;
        RECT 2954.800 2588.370 2957.800 2588.380 ;
        RECT 0.000 2574.980 2920.000 2586.780 ;
        RECT -28.780 2573.380 -25.780 2573.390 ;
        RECT 2945.400 2573.380 2948.400 2573.390 ;
        RECT -28.780 2570.370 -25.780 2570.380 ;
        RECT 2945.400 2570.370 2948.400 2570.380 ;
        RECT 0.000 2556.980 2920.000 2568.780 ;
        RECT -19.380 2555.380 -16.380 2555.390 ;
        RECT 2936.000 2555.380 2939.000 2555.390 ;
        RECT -19.380 2552.370 -16.380 2552.380 ;
        RECT 2936.000 2552.370 2939.000 2552.380 ;
        RECT 0.000 2538.740 2920.000 2550.780 ;
        RECT -9.980 2537.140 -6.980 2537.150 ;
        RECT 2926.600 2537.140 2929.600 2537.150 ;
        RECT -9.980 2534.130 -6.980 2534.140 ;
        RECT 2926.600 2534.130 2929.600 2534.140 ;
        RECT 0.000 2502.980 2920.000 2532.540 ;
        RECT -42.880 2501.380 -39.880 2501.390 ;
        RECT 2959.500 2501.380 2962.500 2501.390 ;
        RECT -42.880 2498.370 -39.880 2498.380 ;
        RECT 2959.500 2498.370 2962.500 2498.380 ;
        RECT 0.000 2484.980 2920.000 2496.780 ;
        RECT -33.480 2483.380 -30.480 2483.390 ;
        RECT 2950.100 2483.380 2953.100 2483.390 ;
        RECT -33.480 2480.370 -30.480 2480.380 ;
        RECT 2950.100 2480.370 2953.100 2480.380 ;
        RECT 0.000 2466.980 2920.000 2478.780 ;
        RECT -24.080 2465.380 -21.080 2465.390 ;
        RECT 2940.700 2465.380 2943.700 2465.390 ;
        RECT -24.080 2462.370 -21.080 2462.380 ;
        RECT 2940.700 2462.370 2943.700 2462.380 ;
        RECT 0.000 2448.740 2920.000 2460.780 ;
        RECT -14.680 2447.140 -11.680 2447.150 ;
        RECT 2931.300 2447.140 2934.300 2447.150 ;
        RECT -14.680 2444.130 -11.680 2444.140 ;
        RECT 2931.300 2444.130 2934.300 2444.140 ;
        RECT 0.000 2412.980 2920.000 2442.540 ;
        RECT -38.180 2411.380 -35.180 2411.390 ;
        RECT 2954.800 2411.380 2957.800 2411.390 ;
        RECT -38.180 2408.370 -35.180 2408.380 ;
        RECT 2954.800 2408.370 2957.800 2408.380 ;
        RECT 0.000 2394.980 2920.000 2406.780 ;
        RECT -28.780 2393.380 -25.780 2393.390 ;
        RECT 2945.400 2393.380 2948.400 2393.390 ;
        RECT -28.780 2390.370 -25.780 2390.380 ;
        RECT 2945.400 2390.370 2948.400 2390.380 ;
        RECT 0.000 2376.980 2920.000 2388.780 ;
        RECT -19.380 2375.380 -16.380 2375.390 ;
        RECT 2936.000 2375.380 2939.000 2375.390 ;
        RECT -19.380 2372.370 -16.380 2372.380 ;
        RECT 2936.000 2372.370 2939.000 2372.380 ;
        RECT 0.000 2358.740 2920.000 2370.780 ;
        RECT -9.980 2357.140 -6.980 2357.150 ;
        RECT 2926.600 2357.140 2929.600 2357.150 ;
        RECT -9.980 2354.130 -6.980 2354.140 ;
        RECT 2926.600 2354.130 2929.600 2354.140 ;
        RECT 0.000 2322.980 2920.000 2352.540 ;
        RECT -42.880 2321.380 -39.880 2321.390 ;
        RECT 2959.500 2321.380 2962.500 2321.390 ;
        RECT -42.880 2318.370 -39.880 2318.380 ;
        RECT 2959.500 2318.370 2962.500 2318.380 ;
        RECT 0.000 2304.980 2920.000 2316.780 ;
        RECT -33.480 2303.380 -30.480 2303.390 ;
        RECT 2950.100 2303.380 2953.100 2303.390 ;
        RECT -33.480 2300.370 -30.480 2300.380 ;
        RECT 2950.100 2300.370 2953.100 2300.380 ;
        RECT 0.000 2286.980 2920.000 2298.780 ;
        RECT -24.080 2285.380 -21.080 2285.390 ;
        RECT 2940.700 2285.380 2943.700 2285.390 ;
        RECT -24.080 2282.370 -21.080 2282.380 ;
        RECT 2940.700 2282.370 2943.700 2282.380 ;
        RECT 0.000 2268.740 2920.000 2280.780 ;
        RECT -14.680 2267.140 -11.680 2267.150 ;
        RECT 2931.300 2267.140 2934.300 2267.150 ;
        RECT -14.680 2264.130 -11.680 2264.140 ;
        RECT 2931.300 2264.130 2934.300 2264.140 ;
        RECT 0.000 2232.980 2920.000 2262.540 ;
        RECT -38.180 2231.380 -35.180 2231.390 ;
        RECT 2954.800 2231.380 2957.800 2231.390 ;
        RECT -38.180 2228.370 -35.180 2228.380 ;
        RECT 2954.800 2228.370 2957.800 2228.380 ;
        RECT 0.000 2214.980 2920.000 2226.780 ;
        RECT -28.780 2213.380 -25.780 2213.390 ;
        RECT 2945.400 2213.380 2948.400 2213.390 ;
        RECT -28.780 2210.370 -25.780 2210.380 ;
        RECT 2945.400 2210.370 2948.400 2210.380 ;
        RECT 0.000 2196.980 2920.000 2208.780 ;
        RECT -19.380 2195.380 -16.380 2195.390 ;
        RECT 2936.000 2195.380 2939.000 2195.390 ;
        RECT -19.380 2192.370 -16.380 2192.380 ;
        RECT 2936.000 2192.370 2939.000 2192.380 ;
        RECT 0.000 2178.740 2920.000 2190.780 ;
        RECT -9.980 2177.140 -6.980 2177.150 ;
        RECT 2926.600 2177.140 2929.600 2177.150 ;
        RECT -9.980 2174.130 -6.980 2174.140 ;
        RECT 2926.600 2174.130 2929.600 2174.140 ;
        RECT 0.000 2142.980 2920.000 2172.540 ;
        RECT -42.880 2141.380 -39.880 2141.390 ;
        RECT 2959.500 2141.380 2962.500 2141.390 ;
        RECT -42.880 2138.370 -39.880 2138.380 ;
        RECT 2959.500 2138.370 2962.500 2138.380 ;
        RECT 0.000 2124.980 2920.000 2136.780 ;
        RECT -33.480 2123.380 -30.480 2123.390 ;
        RECT 2950.100 2123.380 2953.100 2123.390 ;
        RECT -33.480 2120.370 -30.480 2120.380 ;
        RECT 2950.100 2120.370 2953.100 2120.380 ;
        RECT 0.000 2106.980 2920.000 2118.780 ;
        RECT -24.080 2105.380 -21.080 2105.390 ;
        RECT 2940.700 2105.380 2943.700 2105.390 ;
        RECT -24.080 2102.370 -21.080 2102.380 ;
        RECT 2940.700 2102.370 2943.700 2102.380 ;
        RECT 0.000 2088.740 2920.000 2100.780 ;
        RECT -14.680 2087.140 -11.680 2087.150 ;
        RECT 2931.300 2087.140 2934.300 2087.150 ;
        RECT -14.680 2084.130 -11.680 2084.140 ;
        RECT 2931.300 2084.130 2934.300 2084.140 ;
        RECT 0.000 2052.980 2920.000 2082.540 ;
        RECT -38.180 2051.380 -35.180 2051.390 ;
        RECT 2954.800 2051.380 2957.800 2051.390 ;
        RECT -38.180 2048.370 -35.180 2048.380 ;
        RECT 2954.800 2048.370 2957.800 2048.380 ;
        RECT 0.000 2034.980 2920.000 2046.780 ;
        RECT -28.780 2033.380 -25.780 2033.390 ;
        RECT 2945.400 2033.380 2948.400 2033.390 ;
        RECT -28.780 2030.370 -25.780 2030.380 ;
        RECT 2945.400 2030.370 2948.400 2030.380 ;
        RECT 0.000 2016.980 2920.000 2028.780 ;
        RECT -19.380 2015.380 -16.380 2015.390 ;
        RECT 2936.000 2015.380 2939.000 2015.390 ;
        RECT -19.380 2012.370 -16.380 2012.380 ;
        RECT 2936.000 2012.370 2939.000 2012.380 ;
        RECT 0.000 1998.740 2920.000 2010.780 ;
        RECT -9.980 1997.140 -6.980 1997.150 ;
        RECT 2926.600 1997.140 2929.600 1997.150 ;
        RECT -9.980 1994.130 -6.980 1994.140 ;
        RECT 2926.600 1994.130 2929.600 1994.140 ;
        RECT 0.000 1962.980 2920.000 1992.540 ;
        RECT -42.880 1961.380 -39.880 1961.390 ;
        RECT 2959.500 1961.380 2962.500 1961.390 ;
        RECT -42.880 1958.370 -39.880 1958.380 ;
        RECT 2959.500 1958.370 2962.500 1958.380 ;
        RECT 0.000 1944.980 2920.000 1956.780 ;
        RECT -33.480 1943.380 -30.480 1943.390 ;
        RECT 2950.100 1943.380 2953.100 1943.390 ;
        RECT -33.480 1940.370 -30.480 1940.380 ;
        RECT 2950.100 1940.370 2953.100 1940.380 ;
        RECT 0.000 1926.980 2920.000 1938.780 ;
        RECT -24.080 1925.380 -21.080 1925.390 ;
        RECT 2940.700 1925.380 2943.700 1925.390 ;
        RECT -24.080 1922.370 -21.080 1922.380 ;
        RECT 2940.700 1922.370 2943.700 1922.380 ;
        RECT 0.000 1908.740 2920.000 1920.780 ;
        RECT -14.680 1907.140 -11.680 1907.150 ;
        RECT 2931.300 1907.140 2934.300 1907.150 ;
        RECT -14.680 1904.130 -11.680 1904.140 ;
        RECT 2931.300 1904.130 2934.300 1904.140 ;
        RECT 0.000 1872.980 2920.000 1902.540 ;
        RECT -38.180 1871.380 -35.180 1871.390 ;
        RECT 2954.800 1871.380 2957.800 1871.390 ;
        RECT -38.180 1868.370 -35.180 1868.380 ;
        RECT 2954.800 1868.370 2957.800 1868.380 ;
        RECT 0.000 1854.980 2920.000 1866.780 ;
        RECT -28.780 1853.380 -25.780 1853.390 ;
        RECT 2945.400 1853.380 2948.400 1853.390 ;
        RECT -28.780 1850.370 -25.780 1850.380 ;
        RECT 2945.400 1850.370 2948.400 1850.380 ;
        RECT 0.000 1836.980 2920.000 1848.780 ;
        RECT -19.380 1835.380 -16.380 1835.390 ;
        RECT 2936.000 1835.380 2939.000 1835.390 ;
        RECT -19.380 1832.370 -16.380 1832.380 ;
        RECT 2936.000 1832.370 2939.000 1832.380 ;
        RECT 0.000 1818.740 2920.000 1830.780 ;
        RECT -9.980 1817.140 -6.980 1817.150 ;
        RECT 2926.600 1817.140 2929.600 1817.150 ;
        RECT -9.980 1814.130 -6.980 1814.140 ;
        RECT 2926.600 1814.130 2929.600 1814.140 ;
        RECT 0.000 1782.980 2920.000 1812.540 ;
        RECT -42.880 1781.380 -39.880 1781.390 ;
        RECT 2959.500 1781.380 2962.500 1781.390 ;
        RECT -42.880 1778.370 -39.880 1778.380 ;
        RECT 2959.500 1778.370 2962.500 1778.380 ;
        RECT 0.000 1764.980 2920.000 1776.780 ;
        RECT -33.480 1763.380 -30.480 1763.390 ;
        RECT 2950.100 1763.380 2953.100 1763.390 ;
        RECT -33.480 1760.370 -30.480 1760.380 ;
        RECT 2950.100 1760.370 2953.100 1760.380 ;
        RECT 0.000 1746.980 2920.000 1758.780 ;
        RECT -24.080 1745.380 -21.080 1745.390 ;
        RECT 2940.700 1745.380 2943.700 1745.390 ;
        RECT -24.080 1742.370 -21.080 1742.380 ;
        RECT 2940.700 1742.370 2943.700 1742.380 ;
        RECT 0.000 1728.740 2920.000 1740.780 ;
        RECT -14.680 1727.140 -11.680 1727.150 ;
        RECT 2931.300 1727.140 2934.300 1727.150 ;
        RECT -14.680 1724.130 -11.680 1724.140 ;
        RECT 2931.300 1724.130 2934.300 1724.140 ;
        RECT 0.000 1692.980 2920.000 1722.540 ;
        RECT -38.180 1691.380 -35.180 1691.390 ;
        RECT 2954.800 1691.380 2957.800 1691.390 ;
        RECT -38.180 1688.370 -35.180 1688.380 ;
        RECT 2954.800 1688.370 2957.800 1688.380 ;
        RECT 0.000 1674.980 2920.000 1686.780 ;
        RECT -28.780 1673.380 -25.780 1673.390 ;
        RECT 2945.400 1673.380 2948.400 1673.390 ;
        RECT -28.780 1670.370 -25.780 1670.380 ;
        RECT 2945.400 1670.370 2948.400 1670.380 ;
        RECT 0.000 1656.980 2920.000 1668.780 ;
        RECT -19.380 1655.380 -16.380 1655.390 ;
        RECT 2936.000 1655.380 2939.000 1655.390 ;
        RECT -19.380 1652.370 -16.380 1652.380 ;
        RECT 2936.000 1652.370 2939.000 1652.380 ;
        RECT 0.000 1638.740 2920.000 1650.780 ;
        RECT -9.980 1637.140 -6.980 1637.150 ;
        RECT 2926.600 1637.140 2929.600 1637.150 ;
        RECT -9.980 1634.130 -6.980 1634.140 ;
        RECT 2926.600 1634.130 2929.600 1634.140 ;
        RECT 0.000 1602.980 2920.000 1632.540 ;
        RECT -42.880 1601.380 -39.880 1601.390 ;
        RECT 2959.500 1601.380 2962.500 1601.390 ;
        RECT -42.880 1598.370 -39.880 1598.380 ;
        RECT 2959.500 1598.370 2962.500 1598.380 ;
        RECT 0.000 1584.980 2920.000 1596.780 ;
        RECT -33.480 1583.380 -30.480 1583.390 ;
        RECT 2950.100 1583.380 2953.100 1583.390 ;
        RECT -33.480 1580.370 -30.480 1580.380 ;
        RECT 2950.100 1580.370 2953.100 1580.380 ;
        RECT 0.000 1566.980 2920.000 1578.780 ;
        RECT -24.080 1565.380 -21.080 1565.390 ;
        RECT 2940.700 1565.380 2943.700 1565.390 ;
        RECT -24.080 1562.370 -21.080 1562.380 ;
        RECT 2940.700 1562.370 2943.700 1562.380 ;
        RECT 0.000 1548.740 2920.000 1560.780 ;
        RECT -14.680 1547.140 -11.680 1547.150 ;
        RECT 2931.300 1547.140 2934.300 1547.150 ;
        RECT -14.680 1544.130 -11.680 1544.140 ;
        RECT 2931.300 1544.130 2934.300 1544.140 ;
        RECT 0.000 1512.980 2920.000 1542.540 ;
        RECT -38.180 1511.380 -35.180 1511.390 ;
        RECT 2954.800 1511.380 2957.800 1511.390 ;
        RECT -38.180 1508.370 -35.180 1508.380 ;
        RECT 2954.800 1508.370 2957.800 1508.380 ;
        RECT 0.000 1494.980 2920.000 1506.780 ;
        RECT -28.780 1493.380 -25.780 1493.390 ;
        RECT 2945.400 1493.380 2948.400 1493.390 ;
        RECT -28.780 1490.370 -25.780 1490.380 ;
        RECT 2945.400 1490.370 2948.400 1490.380 ;
        RECT 0.000 1476.980 2920.000 1488.780 ;
        RECT -19.380 1475.380 -16.380 1475.390 ;
        RECT 2936.000 1475.380 2939.000 1475.390 ;
        RECT -19.380 1472.370 -16.380 1472.380 ;
        RECT 2936.000 1472.370 2939.000 1472.380 ;
        RECT 0.000 1458.740 2920.000 1470.780 ;
        RECT -9.980 1457.140 -6.980 1457.150 ;
        RECT 2926.600 1457.140 2929.600 1457.150 ;
        RECT -9.980 1454.130 -6.980 1454.140 ;
        RECT 2926.600 1454.130 2929.600 1454.140 ;
        RECT 0.000 1422.980 2920.000 1452.540 ;
        RECT -42.880 1421.380 -39.880 1421.390 ;
        RECT 2959.500 1421.380 2962.500 1421.390 ;
        RECT -42.880 1418.370 -39.880 1418.380 ;
        RECT 2959.500 1418.370 2962.500 1418.380 ;
        RECT 0.000 1404.980 2920.000 1416.780 ;
        RECT -33.480 1403.380 -30.480 1403.390 ;
        RECT 2950.100 1403.380 2953.100 1403.390 ;
        RECT -33.480 1400.370 -30.480 1400.380 ;
        RECT 2950.100 1400.370 2953.100 1400.380 ;
        RECT 0.000 1386.980 2920.000 1398.780 ;
        RECT -24.080 1385.380 -21.080 1385.390 ;
        RECT 2940.700 1385.380 2943.700 1385.390 ;
        RECT -24.080 1382.370 -21.080 1382.380 ;
        RECT 2940.700 1382.370 2943.700 1382.380 ;
        RECT 0.000 1368.740 2920.000 1380.780 ;
        RECT -14.680 1367.140 -11.680 1367.150 ;
        RECT 2931.300 1367.140 2934.300 1367.150 ;
        RECT -14.680 1364.130 -11.680 1364.140 ;
        RECT 2931.300 1364.130 2934.300 1364.140 ;
        RECT 0.000 1332.980 2920.000 1362.540 ;
        RECT -38.180 1331.380 -35.180 1331.390 ;
        RECT 2954.800 1331.380 2957.800 1331.390 ;
        RECT -38.180 1328.370 -35.180 1328.380 ;
        RECT 2954.800 1328.370 2957.800 1328.380 ;
        RECT 0.000 1314.980 2920.000 1326.780 ;
        RECT -28.780 1313.380 -25.780 1313.390 ;
        RECT 2945.400 1313.380 2948.400 1313.390 ;
        RECT -28.780 1310.370 -25.780 1310.380 ;
        RECT 2945.400 1310.370 2948.400 1310.380 ;
        RECT 0.000 1296.980 2920.000 1308.780 ;
        RECT -19.380 1295.380 -16.380 1295.390 ;
        RECT 2936.000 1295.380 2939.000 1295.390 ;
        RECT -19.380 1292.370 -16.380 1292.380 ;
        RECT 2936.000 1292.370 2939.000 1292.380 ;
        RECT 0.000 1278.740 2920.000 1290.780 ;
        RECT -9.980 1277.140 -6.980 1277.150 ;
        RECT 2926.600 1277.140 2929.600 1277.150 ;
        RECT -9.980 1274.130 -6.980 1274.140 ;
        RECT 2926.600 1274.130 2929.600 1274.140 ;
        RECT 0.000 1242.980 2920.000 1272.540 ;
        RECT -42.880 1241.380 -39.880 1241.390 ;
        RECT 2959.500 1241.380 2962.500 1241.390 ;
        RECT -42.880 1238.370 -39.880 1238.380 ;
        RECT 2959.500 1238.370 2962.500 1238.380 ;
        RECT 0.000 1224.980 2920.000 1236.780 ;
        RECT -33.480 1223.380 -30.480 1223.390 ;
        RECT 2950.100 1223.380 2953.100 1223.390 ;
        RECT -33.480 1220.370 -30.480 1220.380 ;
        RECT 2950.100 1220.370 2953.100 1220.380 ;
        RECT 0.000 1206.980 2920.000 1218.780 ;
        RECT -24.080 1205.380 -21.080 1205.390 ;
        RECT 2940.700 1205.380 2943.700 1205.390 ;
        RECT -24.080 1202.370 -21.080 1202.380 ;
        RECT 2940.700 1202.370 2943.700 1202.380 ;
        RECT 0.000 1188.740 2920.000 1200.780 ;
        RECT -14.680 1187.140 -11.680 1187.150 ;
        RECT 2931.300 1187.140 2934.300 1187.150 ;
        RECT -14.680 1184.130 -11.680 1184.140 ;
        RECT 2931.300 1184.130 2934.300 1184.140 ;
        RECT 0.000 1152.980 2920.000 1182.540 ;
        RECT -38.180 1151.380 -35.180 1151.390 ;
        RECT 2954.800 1151.380 2957.800 1151.390 ;
        RECT -38.180 1148.370 -35.180 1148.380 ;
        RECT 2954.800 1148.370 2957.800 1148.380 ;
        RECT 0.000 1134.980 2920.000 1146.780 ;
        RECT -28.780 1133.380 -25.780 1133.390 ;
        RECT 2945.400 1133.380 2948.400 1133.390 ;
        RECT -28.780 1130.370 -25.780 1130.380 ;
        RECT 2945.400 1130.370 2948.400 1130.380 ;
        RECT 0.000 1116.980 2920.000 1128.780 ;
        RECT -19.380 1115.380 -16.380 1115.390 ;
        RECT 2936.000 1115.380 2939.000 1115.390 ;
        RECT -19.380 1112.370 -16.380 1112.380 ;
        RECT 2936.000 1112.370 2939.000 1112.380 ;
        RECT 0.000 1098.740 2920.000 1110.780 ;
        RECT -9.980 1097.140 -6.980 1097.150 ;
        RECT 2926.600 1097.140 2929.600 1097.150 ;
        RECT -9.980 1094.130 -6.980 1094.140 ;
        RECT 2926.600 1094.130 2929.600 1094.140 ;
        RECT 0.000 1062.980 2920.000 1092.540 ;
        RECT -42.880 1061.380 -39.880 1061.390 ;
        RECT 2959.500 1061.380 2962.500 1061.390 ;
        RECT -42.880 1058.370 -39.880 1058.380 ;
        RECT 2959.500 1058.370 2962.500 1058.380 ;
        RECT 0.000 1044.980 2920.000 1056.780 ;
        RECT -33.480 1043.380 -30.480 1043.390 ;
        RECT 2950.100 1043.380 2953.100 1043.390 ;
        RECT -33.480 1040.370 -30.480 1040.380 ;
        RECT 2950.100 1040.370 2953.100 1040.380 ;
        RECT 0.000 1026.980 2920.000 1038.780 ;
        RECT -24.080 1025.380 -21.080 1025.390 ;
        RECT 2940.700 1025.380 2943.700 1025.390 ;
        RECT -24.080 1022.370 -21.080 1022.380 ;
        RECT 2940.700 1022.370 2943.700 1022.380 ;
        RECT 0.000 1008.740 2920.000 1020.780 ;
        RECT -14.680 1007.140 -11.680 1007.150 ;
        RECT 2931.300 1007.140 2934.300 1007.150 ;
        RECT -14.680 1004.130 -11.680 1004.140 ;
        RECT 2931.300 1004.130 2934.300 1004.140 ;
        RECT 0.000 972.980 2920.000 1002.540 ;
        RECT -38.180 971.380 -35.180 971.390 ;
        RECT 2954.800 971.380 2957.800 971.390 ;
        RECT -38.180 968.370 -35.180 968.380 ;
        RECT 2954.800 968.370 2957.800 968.380 ;
        RECT 0.000 954.980 2920.000 966.780 ;
        RECT -28.780 953.380 -25.780 953.390 ;
        RECT 2945.400 953.380 2948.400 953.390 ;
        RECT -28.780 950.370 -25.780 950.380 ;
        RECT 2945.400 950.370 2948.400 950.380 ;
        RECT 0.000 936.980 2920.000 948.780 ;
        RECT -19.380 935.380 -16.380 935.390 ;
        RECT 2936.000 935.380 2939.000 935.390 ;
        RECT -19.380 932.370 -16.380 932.380 ;
        RECT 2936.000 932.370 2939.000 932.380 ;
        RECT 0.000 918.740 2920.000 930.780 ;
        RECT -9.980 917.140 -6.980 917.150 ;
        RECT 2926.600 917.140 2929.600 917.150 ;
        RECT -9.980 914.130 -6.980 914.140 ;
        RECT 2926.600 914.130 2929.600 914.140 ;
        RECT 0.000 882.980 2920.000 912.540 ;
        RECT -42.880 881.380 -39.880 881.390 ;
        RECT 2959.500 881.380 2962.500 881.390 ;
        RECT -42.880 878.370 -39.880 878.380 ;
        RECT 2959.500 878.370 2962.500 878.380 ;
        RECT 0.000 864.980 2920.000 876.780 ;
        RECT -33.480 863.380 -30.480 863.390 ;
        RECT 2950.100 863.380 2953.100 863.390 ;
        RECT -33.480 860.370 -30.480 860.380 ;
        RECT 2950.100 860.370 2953.100 860.380 ;
        RECT 0.000 846.980 2920.000 858.780 ;
        RECT -24.080 845.380 -21.080 845.390 ;
        RECT 2940.700 845.380 2943.700 845.390 ;
        RECT -24.080 842.370 -21.080 842.380 ;
        RECT 2940.700 842.370 2943.700 842.380 ;
        RECT 0.000 828.740 2920.000 840.780 ;
        RECT -14.680 827.140 -11.680 827.150 ;
        RECT 2931.300 827.140 2934.300 827.150 ;
        RECT -14.680 824.130 -11.680 824.140 ;
        RECT 2931.300 824.130 2934.300 824.140 ;
        RECT 0.000 792.980 2920.000 822.540 ;
        RECT -38.180 791.380 -35.180 791.390 ;
        RECT 2954.800 791.380 2957.800 791.390 ;
        RECT -38.180 788.370 -35.180 788.380 ;
        RECT 2954.800 788.370 2957.800 788.380 ;
        RECT 0.000 774.980 2920.000 786.780 ;
        RECT -28.780 773.380 -25.780 773.390 ;
        RECT 2945.400 773.380 2948.400 773.390 ;
        RECT -28.780 770.370 -25.780 770.380 ;
        RECT 2945.400 770.370 2948.400 770.380 ;
        RECT 0.000 756.980 2920.000 768.780 ;
        RECT -19.380 755.380 -16.380 755.390 ;
        RECT 2936.000 755.380 2939.000 755.390 ;
        RECT -19.380 752.370 -16.380 752.380 ;
        RECT 2936.000 752.370 2939.000 752.380 ;
        RECT 0.000 738.740 2920.000 750.780 ;
        RECT -9.980 737.140 -6.980 737.150 ;
        RECT 2926.600 737.140 2929.600 737.150 ;
        RECT -9.980 734.130 -6.980 734.140 ;
        RECT 2926.600 734.130 2929.600 734.140 ;
        RECT 0.000 702.980 2920.000 732.540 ;
        RECT -42.880 701.380 -39.880 701.390 ;
        RECT 2959.500 701.380 2962.500 701.390 ;
        RECT -42.880 698.370 -39.880 698.380 ;
        RECT 2959.500 698.370 2962.500 698.380 ;
        RECT 0.000 684.980 2920.000 696.780 ;
        RECT -33.480 683.380 -30.480 683.390 ;
        RECT 2950.100 683.380 2953.100 683.390 ;
        RECT -33.480 680.370 -30.480 680.380 ;
        RECT 2950.100 680.370 2953.100 680.380 ;
        RECT 0.000 666.980 2920.000 678.780 ;
        RECT -24.080 665.380 -21.080 665.390 ;
        RECT 2940.700 665.380 2943.700 665.390 ;
        RECT -24.080 662.370 -21.080 662.380 ;
        RECT 2940.700 662.370 2943.700 662.380 ;
        RECT 0.000 648.740 2920.000 660.780 ;
        RECT -14.680 647.140 -11.680 647.150 ;
        RECT 2931.300 647.140 2934.300 647.150 ;
        RECT -14.680 644.130 -11.680 644.140 ;
        RECT 2931.300 644.130 2934.300 644.140 ;
        RECT 0.000 612.980 2920.000 642.540 ;
        RECT -38.180 611.380 -35.180 611.390 ;
        RECT 2954.800 611.380 2957.800 611.390 ;
        RECT -38.180 608.370 -35.180 608.380 ;
        RECT 2954.800 608.370 2957.800 608.380 ;
        RECT 0.000 594.980 2920.000 606.780 ;
        RECT -28.780 593.380 -25.780 593.390 ;
        RECT 2945.400 593.380 2948.400 593.390 ;
        RECT -28.780 590.370 -25.780 590.380 ;
        RECT 2945.400 590.370 2948.400 590.380 ;
        RECT 0.000 576.980 2920.000 588.780 ;
        RECT -19.380 575.380 -16.380 575.390 ;
        RECT 2936.000 575.380 2939.000 575.390 ;
        RECT -19.380 572.370 -16.380 572.380 ;
        RECT 2936.000 572.370 2939.000 572.380 ;
        RECT 0.000 558.740 2920.000 570.780 ;
        RECT -9.980 557.140 -6.980 557.150 ;
        RECT 2926.600 557.140 2929.600 557.150 ;
        RECT -9.980 554.130 -6.980 554.140 ;
        RECT 2926.600 554.130 2929.600 554.140 ;
        RECT 0.000 522.980 2920.000 552.540 ;
        RECT -42.880 521.380 -39.880 521.390 ;
        RECT 2959.500 521.380 2962.500 521.390 ;
        RECT -42.880 518.370 -39.880 518.380 ;
        RECT 2959.500 518.370 2962.500 518.380 ;
        RECT 0.000 504.980 2920.000 516.780 ;
        RECT -33.480 503.380 -30.480 503.390 ;
        RECT 2950.100 503.380 2953.100 503.390 ;
        RECT -33.480 500.370 -30.480 500.380 ;
        RECT 2950.100 500.370 2953.100 500.380 ;
        RECT 0.000 486.980 2920.000 498.780 ;
        RECT -24.080 485.380 -21.080 485.390 ;
        RECT 2940.700 485.380 2943.700 485.390 ;
        RECT -24.080 482.370 -21.080 482.380 ;
        RECT 2940.700 482.370 2943.700 482.380 ;
        RECT 0.000 468.740 2920.000 480.780 ;
        RECT -14.680 467.140 -11.680 467.150 ;
        RECT 2931.300 467.140 2934.300 467.150 ;
        RECT -14.680 464.130 -11.680 464.140 ;
        RECT 2931.300 464.130 2934.300 464.140 ;
        RECT 0.000 432.980 2920.000 462.540 ;
        RECT -38.180 431.380 -35.180 431.390 ;
        RECT 2954.800 431.380 2957.800 431.390 ;
        RECT -38.180 428.370 -35.180 428.380 ;
        RECT 2954.800 428.370 2957.800 428.380 ;
        RECT 0.000 414.980 2920.000 426.780 ;
        RECT -28.780 413.380 -25.780 413.390 ;
        RECT 2945.400 413.380 2948.400 413.390 ;
        RECT -28.780 410.370 -25.780 410.380 ;
        RECT 2945.400 410.370 2948.400 410.380 ;
        RECT 0.000 396.980 2920.000 408.780 ;
        RECT -19.380 395.380 -16.380 395.390 ;
        RECT 2936.000 395.380 2939.000 395.390 ;
        RECT -19.380 392.370 -16.380 392.380 ;
        RECT 2936.000 392.370 2939.000 392.380 ;
        RECT 0.000 378.740 2920.000 390.780 ;
        RECT -9.980 377.140 -6.980 377.150 ;
        RECT 2926.600 377.140 2929.600 377.150 ;
        RECT -9.980 374.130 -6.980 374.140 ;
        RECT 2926.600 374.130 2929.600 374.140 ;
        RECT 0.000 342.980 2920.000 372.540 ;
        RECT -42.880 341.380 -39.880 341.390 ;
        RECT 2959.500 341.380 2962.500 341.390 ;
        RECT -42.880 338.370 -39.880 338.380 ;
        RECT 2959.500 338.370 2962.500 338.380 ;
        RECT 0.000 324.980 2920.000 336.780 ;
        RECT -33.480 323.380 -30.480 323.390 ;
        RECT 2950.100 323.380 2953.100 323.390 ;
        RECT -33.480 320.370 -30.480 320.380 ;
        RECT 2950.100 320.370 2953.100 320.380 ;
        RECT 0.000 306.980 2920.000 318.780 ;
        RECT -24.080 305.380 -21.080 305.390 ;
        RECT 2940.700 305.380 2943.700 305.390 ;
        RECT -24.080 302.370 -21.080 302.380 ;
        RECT 2940.700 302.370 2943.700 302.380 ;
        RECT 0.000 288.740 2920.000 300.780 ;
        RECT -14.680 287.140 -11.680 287.150 ;
        RECT 2931.300 287.140 2934.300 287.150 ;
        RECT -14.680 284.130 -11.680 284.140 ;
        RECT 2931.300 284.130 2934.300 284.140 ;
        RECT 0.000 252.980 2920.000 282.540 ;
        RECT -38.180 251.380 -35.180 251.390 ;
        RECT 2954.800 251.380 2957.800 251.390 ;
        RECT -38.180 248.370 -35.180 248.380 ;
        RECT 2954.800 248.370 2957.800 248.380 ;
        RECT 0.000 234.980 2920.000 246.780 ;
        RECT -28.780 233.380 -25.780 233.390 ;
        RECT 2945.400 233.380 2948.400 233.390 ;
        RECT -28.780 230.370 -25.780 230.380 ;
        RECT 2945.400 230.370 2948.400 230.380 ;
        RECT 0.000 216.980 2920.000 228.780 ;
        RECT -19.380 215.380 -16.380 215.390 ;
        RECT 2936.000 215.380 2939.000 215.390 ;
        RECT -19.380 212.370 -16.380 212.380 ;
        RECT 2936.000 212.370 2939.000 212.380 ;
        RECT 0.000 198.740 2920.000 210.780 ;
        RECT -9.980 197.140 -6.980 197.150 ;
        RECT 2926.600 197.140 2929.600 197.150 ;
        RECT -9.980 194.130 -6.980 194.140 ;
        RECT 2926.600 194.130 2929.600 194.140 ;
        RECT 0.000 162.980 2920.000 192.540 ;
        RECT -42.880 161.380 -39.880 161.390 ;
        RECT 2959.500 161.380 2962.500 161.390 ;
        RECT -42.880 158.370 -39.880 158.380 ;
        RECT 2959.500 158.370 2962.500 158.380 ;
        RECT 0.000 144.980 2920.000 156.780 ;
        RECT -33.480 143.380 -30.480 143.390 ;
        RECT 2950.100 143.380 2953.100 143.390 ;
        RECT -33.480 140.370 -30.480 140.380 ;
        RECT 2950.100 140.370 2953.100 140.380 ;
        RECT 0.000 126.980 2920.000 138.780 ;
        RECT -24.080 125.380 -21.080 125.390 ;
        RECT 2940.700 125.380 2943.700 125.390 ;
        RECT -24.080 122.370 -21.080 122.380 ;
        RECT 2940.700 122.370 2943.700 122.380 ;
        RECT 0.000 108.740 2920.000 120.780 ;
        RECT -14.680 107.140 -11.680 107.150 ;
        RECT 2931.300 107.140 2934.300 107.150 ;
        RECT -14.680 104.130 -11.680 104.140 ;
        RECT 2931.300 104.130 2934.300 104.140 ;
        RECT 0.000 72.980 2920.000 102.540 ;
        RECT -38.180 71.380 -35.180 71.390 ;
        RECT 2954.800 71.380 2957.800 71.390 ;
        RECT -38.180 68.370 -35.180 68.380 ;
        RECT 2954.800 68.370 2957.800 68.380 ;
        RECT 0.000 54.980 2920.000 66.780 ;
        RECT -28.780 53.380 -25.780 53.390 ;
        RECT 2945.400 53.380 2948.400 53.390 ;
        RECT -28.780 50.370 -25.780 50.380 ;
        RECT 2945.400 50.370 2948.400 50.380 ;
        RECT 0.000 36.980 2920.000 48.780 ;
        RECT -19.380 35.380 -16.380 35.390 ;
        RECT 2936.000 35.380 2939.000 35.390 ;
        RECT -19.380 32.370 -16.380 32.380 ;
        RECT 2936.000 32.370 2939.000 32.380 ;
        RECT 0.000 18.740 2920.000 30.780 ;
        RECT -9.980 17.140 -6.980 17.150 ;
        RECT 2926.600 17.140 2929.600 17.150 ;
        RECT -9.980 14.130 -6.980 14.140 ;
        RECT 2926.600 14.130 2929.600 14.140 ;
        RECT 0.000 0.000 2920.000 12.540 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 9.020 -1.620 12.020 -1.610 ;
        RECT 189.020 -1.620 192.020 -1.610 ;
        RECT 369.020 -1.620 372.020 -1.610 ;
        RECT 549.020 -1.620 552.020 -1.610 ;
        RECT 729.020 -1.620 732.020 -1.610 ;
        RECT 909.020 -1.620 912.020 -1.610 ;
        RECT 1089.020 -1.620 1092.020 -1.610 ;
        RECT 1269.020 -1.620 1272.020 -1.610 ;
        RECT 1449.020 -1.620 1452.020 -1.610 ;
        RECT 1629.020 -1.620 1632.020 -1.610 ;
        RECT 1809.020 -1.620 1812.020 -1.610 ;
        RECT 1989.020 -1.620 1992.020 -1.610 ;
        RECT 2169.020 -1.620 2172.020 -1.610 ;
        RECT 2349.020 -1.620 2352.020 -1.610 ;
        RECT 2529.020 -1.620 2532.020 -1.610 ;
        RECT 2709.020 -1.620 2712.020 -1.610 ;
        RECT 2889.020 -1.620 2892.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 9.020 -4.630 12.020 -4.620 ;
        RECT 189.020 -4.630 192.020 -4.620 ;
        RECT 369.020 -4.630 372.020 -4.620 ;
        RECT 549.020 -4.630 552.020 -4.620 ;
        RECT 729.020 -4.630 732.020 -4.620 ;
        RECT 909.020 -4.630 912.020 -4.620 ;
        RECT 1089.020 -4.630 1092.020 -4.620 ;
        RECT 1269.020 -4.630 1272.020 -4.620 ;
        RECT 1449.020 -4.630 1452.020 -4.620 ;
        RECT 1629.020 -4.630 1632.020 -4.620 ;
        RECT 1809.020 -4.630 1812.020 -4.620 ;
        RECT 1989.020 -4.630 1992.020 -4.620 ;
        RECT 2169.020 -4.630 2172.020 -4.620 ;
        RECT 2349.020 -4.630 2352.020 -4.620 ;
        RECT 2529.020 -4.630 2532.020 -4.620 ;
        RECT 2709.020 -4.630 2712.020 -4.620 ;
        RECT 2889.020 -4.630 2892.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
        RECT -14.680 -6.320 -11.680 -6.310 ;
        RECT 99.020 -6.320 102.020 -6.310 ;
        RECT 279.020 -6.320 282.020 -6.310 ;
        RECT 459.020 -6.320 462.020 -6.310 ;
        RECT 639.020 -6.320 642.020 -6.310 ;
        RECT 819.020 -6.320 822.020 -6.310 ;
        RECT 999.020 -6.320 1002.020 -6.310 ;
        RECT 1179.020 -6.320 1182.020 -6.310 ;
        RECT 1359.020 -6.320 1362.020 -6.310 ;
        RECT 1539.020 -6.320 1542.020 -6.310 ;
        RECT 1719.020 -6.320 1722.020 -6.310 ;
        RECT 1899.020 -6.320 1902.020 -6.310 ;
        RECT 2079.020 -6.320 2082.020 -6.310 ;
        RECT 2259.020 -6.320 2262.020 -6.310 ;
        RECT 2439.020 -6.320 2442.020 -6.310 ;
        RECT 2619.020 -6.320 2622.020 -6.310 ;
        RECT 2799.020 -6.320 2802.020 -6.310 ;
        RECT 2931.300 -6.320 2934.300 -6.310 ;
        RECT -14.680 -9.330 -11.680 -9.320 ;
        RECT 99.020 -9.330 102.020 -9.320 ;
        RECT 279.020 -9.330 282.020 -9.320 ;
        RECT 459.020 -9.330 462.020 -9.320 ;
        RECT 639.020 -9.330 642.020 -9.320 ;
        RECT 819.020 -9.330 822.020 -9.320 ;
        RECT 999.020 -9.330 1002.020 -9.320 ;
        RECT 1179.020 -9.330 1182.020 -9.320 ;
        RECT 1359.020 -9.330 1362.020 -9.320 ;
        RECT 1539.020 -9.330 1542.020 -9.320 ;
        RECT 1719.020 -9.330 1722.020 -9.320 ;
        RECT 1899.020 -9.330 1902.020 -9.320 ;
        RECT 2079.020 -9.330 2082.020 -9.320 ;
        RECT 2259.020 -9.330 2262.020 -9.320 ;
        RECT 2439.020 -9.330 2442.020 -9.320 ;
        RECT 2619.020 -9.330 2622.020 -9.320 ;
        RECT 2799.020 -9.330 2802.020 -9.320 ;
        RECT 2931.300 -9.330 2934.300 -9.320 ;
        RECT -19.380 -11.020 -16.380 -11.010 ;
        RECT 27.020 -11.020 30.020 -11.010 ;
        RECT 207.020 -11.020 210.020 -11.010 ;
        RECT 387.020 -11.020 390.020 -11.010 ;
        RECT 567.020 -11.020 570.020 -11.010 ;
        RECT 747.020 -11.020 750.020 -11.010 ;
        RECT 927.020 -11.020 930.020 -11.010 ;
        RECT 1107.020 -11.020 1110.020 -11.010 ;
        RECT 1287.020 -11.020 1290.020 -11.010 ;
        RECT 1467.020 -11.020 1470.020 -11.010 ;
        RECT 1647.020 -11.020 1650.020 -11.010 ;
        RECT 1827.020 -11.020 1830.020 -11.010 ;
        RECT 2007.020 -11.020 2010.020 -11.010 ;
        RECT 2187.020 -11.020 2190.020 -11.010 ;
        RECT 2367.020 -11.020 2370.020 -11.010 ;
        RECT 2547.020 -11.020 2550.020 -11.010 ;
        RECT 2727.020 -11.020 2730.020 -11.010 ;
        RECT 2907.020 -11.020 2910.020 -11.010 ;
        RECT 2936.000 -11.020 2939.000 -11.010 ;
        RECT -19.380 -14.030 -16.380 -14.020 ;
        RECT 27.020 -14.030 30.020 -14.020 ;
        RECT 207.020 -14.030 210.020 -14.020 ;
        RECT 387.020 -14.030 390.020 -14.020 ;
        RECT 567.020 -14.030 570.020 -14.020 ;
        RECT 747.020 -14.030 750.020 -14.020 ;
        RECT 927.020 -14.030 930.020 -14.020 ;
        RECT 1107.020 -14.030 1110.020 -14.020 ;
        RECT 1287.020 -14.030 1290.020 -14.020 ;
        RECT 1467.020 -14.030 1470.020 -14.020 ;
        RECT 1647.020 -14.030 1650.020 -14.020 ;
        RECT 1827.020 -14.030 1830.020 -14.020 ;
        RECT 2007.020 -14.030 2010.020 -14.020 ;
        RECT 2187.020 -14.030 2190.020 -14.020 ;
        RECT 2367.020 -14.030 2370.020 -14.020 ;
        RECT 2547.020 -14.030 2550.020 -14.020 ;
        RECT 2727.020 -14.030 2730.020 -14.020 ;
        RECT 2907.020 -14.030 2910.020 -14.020 ;
        RECT 2936.000 -14.030 2939.000 -14.020 ;
        RECT -24.080 -15.720 -21.080 -15.710 ;
        RECT 117.020 -15.720 120.020 -15.710 ;
        RECT 297.020 -15.720 300.020 -15.710 ;
        RECT 477.020 -15.720 480.020 -15.710 ;
        RECT 657.020 -15.720 660.020 -15.710 ;
        RECT 837.020 -15.720 840.020 -15.710 ;
        RECT 1017.020 -15.720 1020.020 -15.710 ;
        RECT 1197.020 -15.720 1200.020 -15.710 ;
        RECT 1377.020 -15.720 1380.020 -15.710 ;
        RECT 1557.020 -15.720 1560.020 -15.710 ;
        RECT 1737.020 -15.720 1740.020 -15.710 ;
        RECT 1917.020 -15.720 1920.020 -15.710 ;
        RECT 2097.020 -15.720 2100.020 -15.710 ;
        RECT 2277.020 -15.720 2280.020 -15.710 ;
        RECT 2457.020 -15.720 2460.020 -15.710 ;
        RECT 2637.020 -15.720 2640.020 -15.710 ;
        RECT 2817.020 -15.720 2820.020 -15.710 ;
        RECT 2940.700 -15.720 2943.700 -15.710 ;
        RECT -24.080 -18.730 -21.080 -18.720 ;
        RECT 117.020 -18.730 120.020 -18.720 ;
        RECT 297.020 -18.730 300.020 -18.720 ;
        RECT 477.020 -18.730 480.020 -18.720 ;
        RECT 657.020 -18.730 660.020 -18.720 ;
        RECT 837.020 -18.730 840.020 -18.720 ;
        RECT 1017.020 -18.730 1020.020 -18.720 ;
        RECT 1197.020 -18.730 1200.020 -18.720 ;
        RECT 1377.020 -18.730 1380.020 -18.720 ;
        RECT 1557.020 -18.730 1560.020 -18.720 ;
        RECT 1737.020 -18.730 1740.020 -18.720 ;
        RECT 1917.020 -18.730 1920.020 -18.720 ;
        RECT 2097.020 -18.730 2100.020 -18.720 ;
        RECT 2277.020 -18.730 2280.020 -18.720 ;
        RECT 2457.020 -18.730 2460.020 -18.720 ;
        RECT 2637.020 -18.730 2640.020 -18.720 ;
        RECT 2817.020 -18.730 2820.020 -18.720 ;
        RECT 2940.700 -18.730 2943.700 -18.720 ;
        RECT -28.780 -20.420 -25.780 -20.410 ;
        RECT 45.020 -20.420 48.020 -20.410 ;
        RECT 225.020 -20.420 228.020 -20.410 ;
        RECT 405.020 -20.420 408.020 -20.410 ;
        RECT 585.020 -20.420 588.020 -20.410 ;
        RECT 765.020 -20.420 768.020 -20.410 ;
        RECT 945.020 -20.420 948.020 -20.410 ;
        RECT 1125.020 -20.420 1128.020 -20.410 ;
        RECT 1305.020 -20.420 1308.020 -20.410 ;
        RECT 1485.020 -20.420 1488.020 -20.410 ;
        RECT 1665.020 -20.420 1668.020 -20.410 ;
        RECT 1845.020 -20.420 1848.020 -20.410 ;
        RECT 2025.020 -20.420 2028.020 -20.410 ;
        RECT 2205.020 -20.420 2208.020 -20.410 ;
        RECT 2385.020 -20.420 2388.020 -20.410 ;
        RECT 2565.020 -20.420 2568.020 -20.410 ;
        RECT 2745.020 -20.420 2748.020 -20.410 ;
        RECT 2945.400 -20.420 2948.400 -20.410 ;
        RECT -28.780 -23.430 -25.780 -23.420 ;
        RECT 45.020 -23.430 48.020 -23.420 ;
        RECT 225.020 -23.430 228.020 -23.420 ;
        RECT 405.020 -23.430 408.020 -23.420 ;
        RECT 585.020 -23.430 588.020 -23.420 ;
        RECT 765.020 -23.430 768.020 -23.420 ;
        RECT 945.020 -23.430 948.020 -23.420 ;
        RECT 1125.020 -23.430 1128.020 -23.420 ;
        RECT 1305.020 -23.430 1308.020 -23.420 ;
        RECT 1485.020 -23.430 1488.020 -23.420 ;
        RECT 1665.020 -23.430 1668.020 -23.420 ;
        RECT 1845.020 -23.430 1848.020 -23.420 ;
        RECT 2025.020 -23.430 2028.020 -23.420 ;
        RECT 2205.020 -23.430 2208.020 -23.420 ;
        RECT 2385.020 -23.430 2388.020 -23.420 ;
        RECT 2565.020 -23.430 2568.020 -23.420 ;
        RECT 2745.020 -23.430 2748.020 -23.420 ;
        RECT 2945.400 -23.430 2948.400 -23.420 ;
        RECT -33.480 -25.120 -30.480 -25.110 ;
        RECT 135.020 -25.120 138.020 -25.110 ;
        RECT 315.020 -25.120 318.020 -25.110 ;
        RECT 495.020 -25.120 498.020 -25.110 ;
        RECT 675.020 -25.120 678.020 -25.110 ;
        RECT 855.020 -25.120 858.020 -25.110 ;
        RECT 1035.020 -25.120 1038.020 -25.110 ;
        RECT 1215.020 -25.120 1218.020 -25.110 ;
        RECT 1395.020 -25.120 1398.020 -25.110 ;
        RECT 1575.020 -25.120 1578.020 -25.110 ;
        RECT 1755.020 -25.120 1758.020 -25.110 ;
        RECT 1935.020 -25.120 1938.020 -25.110 ;
        RECT 2115.020 -25.120 2118.020 -25.110 ;
        RECT 2295.020 -25.120 2298.020 -25.110 ;
        RECT 2475.020 -25.120 2478.020 -25.110 ;
        RECT 2655.020 -25.120 2658.020 -25.110 ;
        RECT 2835.020 -25.120 2838.020 -25.110 ;
        RECT 2950.100 -25.120 2953.100 -25.110 ;
        RECT -33.480 -28.130 -30.480 -28.120 ;
        RECT 135.020 -28.130 138.020 -28.120 ;
        RECT 315.020 -28.130 318.020 -28.120 ;
        RECT 495.020 -28.130 498.020 -28.120 ;
        RECT 675.020 -28.130 678.020 -28.120 ;
        RECT 855.020 -28.130 858.020 -28.120 ;
        RECT 1035.020 -28.130 1038.020 -28.120 ;
        RECT 1215.020 -28.130 1218.020 -28.120 ;
        RECT 1395.020 -28.130 1398.020 -28.120 ;
        RECT 1575.020 -28.130 1578.020 -28.120 ;
        RECT 1755.020 -28.130 1758.020 -28.120 ;
        RECT 1935.020 -28.130 1938.020 -28.120 ;
        RECT 2115.020 -28.130 2118.020 -28.120 ;
        RECT 2295.020 -28.130 2298.020 -28.120 ;
        RECT 2475.020 -28.130 2478.020 -28.120 ;
        RECT 2655.020 -28.130 2658.020 -28.120 ;
        RECT 2835.020 -28.130 2838.020 -28.120 ;
        RECT 2950.100 -28.130 2953.100 -28.120 ;
        RECT -38.180 -29.820 -35.180 -29.810 ;
        RECT 63.020 -29.820 66.020 -29.810 ;
        RECT 243.020 -29.820 246.020 -29.810 ;
        RECT 423.020 -29.820 426.020 -29.810 ;
        RECT 603.020 -29.820 606.020 -29.810 ;
        RECT 783.020 -29.820 786.020 -29.810 ;
        RECT 963.020 -29.820 966.020 -29.810 ;
        RECT 1143.020 -29.820 1146.020 -29.810 ;
        RECT 1323.020 -29.820 1326.020 -29.810 ;
        RECT 1503.020 -29.820 1506.020 -29.810 ;
        RECT 1683.020 -29.820 1686.020 -29.810 ;
        RECT 1863.020 -29.820 1866.020 -29.810 ;
        RECT 2043.020 -29.820 2046.020 -29.810 ;
        RECT 2223.020 -29.820 2226.020 -29.810 ;
        RECT 2403.020 -29.820 2406.020 -29.810 ;
        RECT 2583.020 -29.820 2586.020 -29.810 ;
        RECT 2763.020 -29.820 2766.020 -29.810 ;
        RECT 2954.800 -29.820 2957.800 -29.810 ;
        RECT -38.180 -32.830 -35.180 -32.820 ;
        RECT 63.020 -32.830 66.020 -32.820 ;
        RECT 243.020 -32.830 246.020 -32.820 ;
        RECT 423.020 -32.830 426.020 -32.820 ;
        RECT 603.020 -32.830 606.020 -32.820 ;
        RECT 783.020 -32.830 786.020 -32.820 ;
        RECT 963.020 -32.830 966.020 -32.820 ;
        RECT 1143.020 -32.830 1146.020 -32.820 ;
        RECT 1323.020 -32.830 1326.020 -32.820 ;
        RECT 1503.020 -32.830 1506.020 -32.820 ;
        RECT 1683.020 -32.830 1686.020 -32.820 ;
        RECT 1863.020 -32.830 1866.020 -32.820 ;
        RECT 2043.020 -32.830 2046.020 -32.820 ;
        RECT 2223.020 -32.830 2226.020 -32.820 ;
        RECT 2403.020 -32.830 2406.020 -32.820 ;
        RECT 2583.020 -32.830 2586.020 -32.820 ;
        RECT 2763.020 -32.830 2766.020 -32.820 ;
        RECT 2954.800 -32.830 2957.800 -32.820 ;
        RECT -42.880 -34.520 -39.880 -34.510 ;
        RECT 153.020 -34.520 156.020 -34.510 ;
        RECT 333.020 -34.520 336.020 -34.510 ;
        RECT 513.020 -34.520 516.020 -34.510 ;
        RECT 693.020 -34.520 696.020 -34.510 ;
        RECT 873.020 -34.520 876.020 -34.510 ;
        RECT 1053.020 -34.520 1056.020 -34.510 ;
        RECT 1233.020 -34.520 1236.020 -34.510 ;
        RECT 1413.020 -34.520 1416.020 -34.510 ;
        RECT 1593.020 -34.520 1596.020 -34.510 ;
        RECT 1773.020 -34.520 1776.020 -34.510 ;
        RECT 1953.020 -34.520 1956.020 -34.510 ;
        RECT 2133.020 -34.520 2136.020 -34.510 ;
        RECT 2313.020 -34.520 2316.020 -34.510 ;
        RECT 2493.020 -34.520 2496.020 -34.510 ;
        RECT 2673.020 -34.520 2676.020 -34.510 ;
        RECT 2853.020 -34.520 2856.020 -34.510 ;
        RECT 2959.500 -34.520 2962.500 -34.510 ;
        RECT -42.880 -37.530 -39.880 -37.520 ;
        RECT 153.020 -37.530 156.020 -37.520 ;
        RECT 333.020 -37.530 336.020 -37.520 ;
        RECT 513.020 -37.530 516.020 -37.520 ;
        RECT 693.020 -37.530 696.020 -37.520 ;
        RECT 873.020 -37.530 876.020 -37.520 ;
        RECT 1053.020 -37.530 1056.020 -37.520 ;
        RECT 1233.020 -37.530 1236.020 -37.520 ;
        RECT 1413.020 -37.530 1416.020 -37.520 ;
        RECT 1593.020 -37.530 1596.020 -37.520 ;
        RECT 1773.020 -37.530 1776.020 -37.520 ;
        RECT 1953.020 -37.530 1956.020 -37.520 ;
        RECT 2133.020 -37.530 2136.020 -37.520 ;
        RECT 2313.020 -37.530 2316.020 -37.520 ;
        RECT 2493.020 -37.530 2496.020 -37.520 ;
        RECT 2673.020 -37.530 2676.020 -37.520 ;
        RECT 2853.020 -37.530 2856.020 -37.520 ;
        RECT 2959.500 -37.530 2962.500 -37.520 ;
  END
END user_project_wrapper
END LIBRARY

