magic
tech sky130A
magscale 1 2
timestamp 1623702531
<< obsli1 >>
rect 1104 1377 178848 117521
<< obsm1 >>
rect 474 756 179570 118040
<< metal2 >>
rect 478 119200 534 120000
rect 1398 119200 1454 120000
rect 2410 119200 2466 120000
rect 3422 119200 3478 120000
rect 4342 119200 4398 120000
rect 5354 119200 5410 120000
rect 6366 119200 6422 120000
rect 7286 119200 7342 120000
rect 8298 119200 8354 120000
rect 9310 119200 9366 120000
rect 10230 119200 10286 120000
rect 11242 119200 11298 120000
rect 12254 119200 12310 120000
rect 13266 119200 13322 120000
rect 14186 119200 14242 120000
rect 15198 119200 15254 120000
rect 16210 119200 16266 120000
rect 17130 119200 17186 120000
rect 18142 119200 18198 120000
rect 19154 119200 19210 120000
rect 20074 119200 20130 120000
rect 21086 119200 21142 120000
rect 22098 119200 22154 120000
rect 23018 119200 23074 120000
rect 24030 119200 24086 120000
rect 25042 119200 25098 120000
rect 26054 119200 26110 120000
rect 26974 119200 27030 120000
rect 27986 119200 28042 120000
rect 28998 119200 29054 120000
rect 29918 119200 29974 120000
rect 30930 119200 30986 120000
rect 31942 119200 31998 120000
rect 32862 119200 32918 120000
rect 33874 119200 33930 120000
rect 34886 119200 34942 120000
rect 35806 119200 35862 120000
rect 36818 119200 36874 120000
rect 37830 119200 37886 120000
rect 38842 119200 38898 120000
rect 39762 119200 39818 120000
rect 40774 119200 40830 120000
rect 41786 119200 41842 120000
rect 42706 119200 42762 120000
rect 43718 119200 43774 120000
rect 44730 119200 44786 120000
rect 45650 119200 45706 120000
rect 46662 119200 46718 120000
rect 47674 119200 47730 120000
rect 48686 119200 48742 120000
rect 49606 119200 49662 120000
rect 50618 119200 50674 120000
rect 51630 119200 51686 120000
rect 52550 119200 52606 120000
rect 53562 119200 53618 120000
rect 54574 119200 54630 120000
rect 55494 119200 55550 120000
rect 56506 119200 56562 120000
rect 57518 119200 57574 120000
rect 58438 119200 58494 120000
rect 59450 119200 59506 120000
rect 60462 119200 60518 120000
rect 61474 119200 61530 120000
rect 62394 119200 62450 120000
rect 63406 119200 63462 120000
rect 64418 119200 64474 120000
rect 65338 119200 65394 120000
rect 66350 119200 66406 120000
rect 67362 119200 67418 120000
rect 68282 119200 68338 120000
rect 69294 119200 69350 120000
rect 70306 119200 70362 120000
rect 71226 119200 71282 120000
rect 72238 119200 72294 120000
rect 73250 119200 73306 120000
rect 74262 119200 74318 120000
rect 75182 119200 75238 120000
rect 76194 119200 76250 120000
rect 77206 119200 77262 120000
rect 78126 119200 78182 120000
rect 79138 119200 79194 120000
rect 80150 119200 80206 120000
rect 81070 119200 81126 120000
rect 82082 119200 82138 120000
rect 83094 119200 83150 120000
rect 84014 119200 84070 120000
rect 85026 119200 85082 120000
rect 86038 119200 86094 120000
rect 87050 119200 87106 120000
rect 87970 119200 88026 120000
rect 88982 119200 89038 120000
rect 89994 119200 90050 120000
rect 90914 119200 90970 120000
rect 91926 119200 91982 120000
rect 92938 119200 92994 120000
rect 93858 119200 93914 120000
rect 94870 119200 94926 120000
rect 95882 119200 95938 120000
rect 96894 119200 96950 120000
rect 97814 119200 97870 120000
rect 98826 119200 98882 120000
rect 99838 119200 99894 120000
rect 100758 119200 100814 120000
rect 101770 119200 101826 120000
rect 102782 119200 102838 120000
rect 103702 119200 103758 120000
rect 104714 119200 104770 120000
rect 105726 119200 105782 120000
rect 106646 119200 106702 120000
rect 107658 119200 107714 120000
rect 108670 119200 108726 120000
rect 109682 119200 109738 120000
rect 110602 119200 110658 120000
rect 111614 119200 111670 120000
rect 112626 119200 112682 120000
rect 113546 119200 113602 120000
rect 114558 119200 114614 120000
rect 115570 119200 115626 120000
rect 116490 119200 116546 120000
rect 117502 119200 117558 120000
rect 118514 119200 118570 120000
rect 119434 119200 119490 120000
rect 120446 119200 120502 120000
rect 121458 119200 121514 120000
rect 122470 119200 122526 120000
rect 123390 119200 123446 120000
rect 124402 119200 124458 120000
rect 125414 119200 125470 120000
rect 126334 119200 126390 120000
rect 127346 119200 127402 120000
rect 128358 119200 128414 120000
rect 129278 119200 129334 120000
rect 130290 119200 130346 120000
rect 131302 119200 131358 120000
rect 132222 119200 132278 120000
rect 133234 119200 133290 120000
rect 134246 119200 134302 120000
rect 135258 119200 135314 120000
rect 136178 119200 136234 120000
rect 137190 119200 137246 120000
rect 138202 119200 138258 120000
rect 139122 119200 139178 120000
rect 140134 119200 140190 120000
rect 141146 119200 141202 120000
rect 142066 119200 142122 120000
rect 143078 119200 143134 120000
rect 144090 119200 144146 120000
rect 145102 119200 145158 120000
rect 146022 119200 146078 120000
rect 147034 119200 147090 120000
rect 148046 119200 148102 120000
rect 148966 119200 149022 120000
rect 149978 119200 150034 120000
rect 150990 119200 151046 120000
rect 151910 119200 151966 120000
rect 152922 119200 152978 120000
rect 153934 119200 153990 120000
rect 154854 119200 154910 120000
rect 155866 119200 155922 120000
rect 156878 119200 156934 120000
rect 157890 119200 157946 120000
rect 158810 119200 158866 120000
rect 159822 119200 159878 120000
rect 160834 119200 160890 120000
rect 161754 119200 161810 120000
rect 162766 119200 162822 120000
rect 163778 119200 163834 120000
rect 164698 119200 164754 120000
rect 165710 119200 165766 120000
rect 166722 119200 166778 120000
rect 167642 119200 167698 120000
rect 168654 119200 168710 120000
rect 169666 119200 169722 120000
rect 170678 119200 170734 120000
rect 171598 119200 171654 120000
rect 172610 119200 172666 120000
rect 173622 119200 173678 120000
rect 174542 119200 174598 120000
rect 175554 119200 175610 120000
rect 176566 119200 176622 120000
rect 177486 119200 177542 120000
rect 178498 119200 178554 120000
rect 179510 119200 179566 120000
rect 662 0 718 800
rect 1950 0 2006 800
rect 3330 0 3386 800
rect 4710 0 4766 800
rect 6090 0 6146 800
rect 7470 0 7526 800
rect 8758 0 8814 800
rect 10138 0 10194 800
rect 11518 0 11574 800
rect 12898 0 12954 800
rect 14278 0 14334 800
rect 15658 0 15714 800
rect 16946 0 17002 800
rect 18326 0 18382 800
rect 19706 0 19762 800
rect 21086 0 21142 800
rect 22466 0 22522 800
rect 23846 0 23902 800
rect 25134 0 25190 800
rect 26514 0 26570 800
rect 27894 0 27950 800
rect 29274 0 29330 800
rect 30654 0 30710 800
rect 31942 0 31998 800
rect 33322 0 33378 800
rect 34702 0 34758 800
rect 36082 0 36138 800
rect 37462 0 37518 800
rect 38842 0 38898 800
rect 40130 0 40186 800
rect 41510 0 41566 800
rect 42890 0 42946 800
rect 44270 0 44326 800
rect 45650 0 45706 800
rect 47030 0 47086 800
rect 48318 0 48374 800
rect 49698 0 49754 800
rect 51078 0 51134 800
rect 52458 0 52514 800
rect 53838 0 53894 800
rect 55218 0 55274 800
rect 56506 0 56562 800
rect 57886 0 57942 800
rect 59266 0 59322 800
rect 60646 0 60702 800
rect 62026 0 62082 800
rect 63314 0 63370 800
rect 64694 0 64750 800
rect 66074 0 66130 800
rect 67454 0 67510 800
rect 68834 0 68890 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 72882 0 72938 800
rect 74262 0 74318 800
rect 75642 0 75698 800
rect 77022 0 77078 800
rect 78402 0 78458 800
rect 79690 0 79746 800
rect 81070 0 81126 800
rect 82450 0 82506 800
rect 83830 0 83886 800
rect 85210 0 85266 800
rect 86590 0 86646 800
rect 87878 0 87934 800
rect 89258 0 89314 800
rect 90638 0 90694 800
rect 92018 0 92074 800
rect 93398 0 93454 800
rect 94686 0 94742 800
rect 96066 0 96122 800
rect 97446 0 97502 800
rect 98826 0 98882 800
rect 100206 0 100262 800
rect 101586 0 101642 800
rect 102874 0 102930 800
rect 104254 0 104310 800
rect 105634 0 105690 800
rect 107014 0 107070 800
rect 108394 0 108450 800
rect 109774 0 109830 800
rect 111062 0 111118 800
rect 112442 0 112498 800
rect 113822 0 113878 800
rect 115202 0 115258 800
rect 116582 0 116638 800
rect 117962 0 118018 800
rect 119250 0 119306 800
rect 120630 0 120686 800
rect 122010 0 122066 800
rect 123390 0 123446 800
rect 124770 0 124826 800
rect 126058 0 126114 800
rect 127438 0 127494 800
rect 128818 0 128874 800
rect 130198 0 130254 800
rect 131578 0 131634 800
rect 132958 0 133014 800
rect 134246 0 134302 800
rect 135626 0 135682 800
rect 137006 0 137062 800
rect 138386 0 138442 800
rect 139766 0 139822 800
rect 141146 0 141202 800
rect 142434 0 142490 800
rect 143814 0 143870 800
rect 145194 0 145250 800
rect 146574 0 146630 800
rect 147954 0 148010 800
rect 149334 0 149390 800
rect 150622 0 150678 800
rect 152002 0 152058 800
rect 153382 0 153438 800
rect 154762 0 154818 800
rect 156142 0 156198 800
rect 157430 0 157486 800
rect 158810 0 158866 800
rect 160190 0 160246 800
rect 161570 0 161626 800
rect 162950 0 163006 800
rect 164330 0 164386 800
rect 165618 0 165674 800
rect 166998 0 167054 800
rect 168378 0 168434 800
rect 169758 0 169814 800
rect 171138 0 171194 800
rect 172518 0 172574 800
rect 173806 0 173862 800
rect 175186 0 175242 800
rect 176566 0 176622 800
rect 177946 0 178002 800
rect 179326 0 179382 800
<< obsm2 >>
rect 590 119144 1342 119785
rect 1510 119144 2354 119785
rect 2522 119144 3366 119785
rect 3534 119144 4286 119785
rect 4454 119144 5298 119785
rect 5466 119144 6310 119785
rect 6478 119144 7230 119785
rect 7398 119144 8242 119785
rect 8410 119144 9254 119785
rect 9422 119144 10174 119785
rect 10342 119144 11186 119785
rect 11354 119144 12198 119785
rect 12366 119144 13210 119785
rect 13378 119144 14130 119785
rect 14298 119144 15142 119785
rect 15310 119144 16154 119785
rect 16322 119144 17074 119785
rect 17242 119144 18086 119785
rect 18254 119144 19098 119785
rect 19266 119144 20018 119785
rect 20186 119144 21030 119785
rect 21198 119144 22042 119785
rect 22210 119144 22962 119785
rect 23130 119144 23974 119785
rect 24142 119144 24986 119785
rect 25154 119144 25998 119785
rect 26166 119144 26918 119785
rect 27086 119144 27930 119785
rect 28098 119144 28942 119785
rect 29110 119144 29862 119785
rect 30030 119144 30874 119785
rect 31042 119144 31886 119785
rect 32054 119144 32806 119785
rect 32974 119144 33818 119785
rect 33986 119144 34830 119785
rect 34998 119144 35750 119785
rect 35918 119144 36762 119785
rect 36930 119144 37774 119785
rect 37942 119144 38786 119785
rect 38954 119144 39706 119785
rect 39874 119144 40718 119785
rect 40886 119144 41730 119785
rect 41898 119144 42650 119785
rect 42818 119144 43662 119785
rect 43830 119144 44674 119785
rect 44842 119144 45594 119785
rect 45762 119144 46606 119785
rect 46774 119144 47618 119785
rect 47786 119144 48630 119785
rect 48798 119144 49550 119785
rect 49718 119144 50562 119785
rect 50730 119144 51574 119785
rect 51742 119144 52494 119785
rect 52662 119144 53506 119785
rect 53674 119144 54518 119785
rect 54686 119144 55438 119785
rect 55606 119144 56450 119785
rect 56618 119144 57462 119785
rect 57630 119144 58382 119785
rect 58550 119144 59394 119785
rect 59562 119144 60406 119785
rect 60574 119144 61418 119785
rect 61586 119144 62338 119785
rect 62506 119144 63350 119785
rect 63518 119144 64362 119785
rect 64530 119144 65282 119785
rect 65450 119144 66294 119785
rect 66462 119144 67306 119785
rect 67474 119144 68226 119785
rect 68394 119144 69238 119785
rect 69406 119144 70250 119785
rect 70418 119144 71170 119785
rect 71338 119144 72182 119785
rect 72350 119144 73194 119785
rect 73362 119144 74206 119785
rect 74374 119144 75126 119785
rect 75294 119144 76138 119785
rect 76306 119144 77150 119785
rect 77318 119144 78070 119785
rect 78238 119144 79082 119785
rect 79250 119144 80094 119785
rect 80262 119144 81014 119785
rect 81182 119144 82026 119785
rect 82194 119144 83038 119785
rect 83206 119144 83958 119785
rect 84126 119144 84970 119785
rect 85138 119144 85982 119785
rect 86150 119144 86994 119785
rect 87162 119144 87914 119785
rect 88082 119144 88926 119785
rect 89094 119144 89938 119785
rect 90106 119144 90858 119785
rect 91026 119144 91870 119785
rect 92038 119144 92882 119785
rect 93050 119144 93802 119785
rect 93970 119144 94814 119785
rect 94982 119144 95826 119785
rect 95994 119144 96838 119785
rect 97006 119144 97758 119785
rect 97926 119144 98770 119785
rect 98938 119144 99782 119785
rect 99950 119144 100702 119785
rect 100870 119144 101714 119785
rect 101882 119144 102726 119785
rect 102894 119144 103646 119785
rect 103814 119144 104658 119785
rect 104826 119144 105670 119785
rect 105838 119144 106590 119785
rect 106758 119144 107602 119785
rect 107770 119144 108614 119785
rect 108782 119144 109626 119785
rect 109794 119144 110546 119785
rect 110714 119144 111558 119785
rect 111726 119144 112570 119785
rect 112738 119144 113490 119785
rect 113658 119144 114502 119785
rect 114670 119144 115514 119785
rect 115682 119144 116434 119785
rect 116602 119144 117446 119785
rect 117614 119144 118458 119785
rect 118626 119144 119378 119785
rect 119546 119144 120390 119785
rect 120558 119144 121402 119785
rect 121570 119144 122414 119785
rect 122582 119144 123334 119785
rect 123502 119144 124346 119785
rect 124514 119144 125358 119785
rect 125526 119144 126278 119785
rect 126446 119144 127290 119785
rect 127458 119144 128302 119785
rect 128470 119144 129222 119785
rect 129390 119144 130234 119785
rect 130402 119144 131246 119785
rect 131414 119144 132166 119785
rect 132334 119144 133178 119785
rect 133346 119144 134190 119785
rect 134358 119144 135202 119785
rect 135370 119144 136122 119785
rect 136290 119144 137134 119785
rect 137302 119144 138146 119785
rect 138314 119144 139066 119785
rect 139234 119144 140078 119785
rect 140246 119144 141090 119785
rect 141258 119144 142010 119785
rect 142178 119144 143022 119785
rect 143190 119144 144034 119785
rect 144202 119144 145046 119785
rect 145214 119144 145966 119785
rect 146134 119144 146978 119785
rect 147146 119144 147990 119785
rect 148158 119144 148910 119785
rect 149078 119144 149922 119785
rect 150090 119144 150934 119785
rect 151102 119144 151854 119785
rect 152022 119144 152866 119785
rect 153034 119144 153878 119785
rect 154046 119144 154798 119785
rect 154966 119144 155810 119785
rect 155978 119144 156822 119785
rect 156990 119144 157834 119785
rect 158002 119144 158754 119785
rect 158922 119144 159766 119785
rect 159934 119144 160778 119785
rect 160946 119144 161698 119785
rect 161866 119144 162710 119785
rect 162878 119144 163722 119785
rect 163890 119144 164642 119785
rect 164810 119144 165654 119785
rect 165822 119144 166666 119785
rect 166834 119144 167586 119785
rect 167754 119144 168598 119785
rect 168766 119144 169610 119785
rect 169778 119144 170622 119785
rect 170790 119144 171542 119785
rect 171710 119144 172554 119785
rect 172722 119144 173566 119785
rect 173734 119144 174486 119785
rect 174654 119144 175498 119785
rect 175666 119144 176510 119785
rect 176678 119144 177430 119785
rect 177598 119144 178442 119785
rect 178610 119144 179454 119785
rect 480 856 179564 119144
rect 480 167 606 856
rect 774 167 1894 856
rect 2062 167 3274 856
rect 3442 167 4654 856
rect 4822 167 6034 856
rect 6202 167 7414 856
rect 7582 167 8702 856
rect 8870 167 10082 856
rect 10250 167 11462 856
rect 11630 167 12842 856
rect 13010 167 14222 856
rect 14390 167 15602 856
rect 15770 167 16890 856
rect 17058 167 18270 856
rect 18438 167 19650 856
rect 19818 167 21030 856
rect 21198 167 22410 856
rect 22578 167 23790 856
rect 23958 167 25078 856
rect 25246 167 26458 856
rect 26626 167 27838 856
rect 28006 167 29218 856
rect 29386 167 30598 856
rect 30766 167 31886 856
rect 32054 167 33266 856
rect 33434 167 34646 856
rect 34814 167 36026 856
rect 36194 167 37406 856
rect 37574 167 38786 856
rect 38954 167 40074 856
rect 40242 167 41454 856
rect 41622 167 42834 856
rect 43002 167 44214 856
rect 44382 167 45594 856
rect 45762 167 46974 856
rect 47142 167 48262 856
rect 48430 167 49642 856
rect 49810 167 51022 856
rect 51190 167 52402 856
rect 52570 167 53782 856
rect 53950 167 55162 856
rect 55330 167 56450 856
rect 56618 167 57830 856
rect 57998 167 59210 856
rect 59378 167 60590 856
rect 60758 167 61970 856
rect 62138 167 63258 856
rect 63426 167 64638 856
rect 64806 167 66018 856
rect 66186 167 67398 856
rect 67566 167 68778 856
rect 68946 167 70158 856
rect 70326 167 71446 856
rect 71614 167 72826 856
rect 72994 167 74206 856
rect 74374 167 75586 856
rect 75754 167 76966 856
rect 77134 167 78346 856
rect 78514 167 79634 856
rect 79802 167 81014 856
rect 81182 167 82394 856
rect 82562 167 83774 856
rect 83942 167 85154 856
rect 85322 167 86534 856
rect 86702 167 87822 856
rect 87990 167 89202 856
rect 89370 167 90582 856
rect 90750 167 91962 856
rect 92130 167 93342 856
rect 93510 167 94630 856
rect 94798 167 96010 856
rect 96178 167 97390 856
rect 97558 167 98770 856
rect 98938 167 100150 856
rect 100318 167 101530 856
rect 101698 167 102818 856
rect 102986 167 104198 856
rect 104366 167 105578 856
rect 105746 167 106958 856
rect 107126 167 108338 856
rect 108506 167 109718 856
rect 109886 167 111006 856
rect 111174 167 112386 856
rect 112554 167 113766 856
rect 113934 167 115146 856
rect 115314 167 116526 856
rect 116694 167 117906 856
rect 118074 167 119194 856
rect 119362 167 120574 856
rect 120742 167 121954 856
rect 122122 167 123334 856
rect 123502 167 124714 856
rect 124882 167 126002 856
rect 126170 167 127382 856
rect 127550 167 128762 856
rect 128930 167 130142 856
rect 130310 167 131522 856
rect 131690 167 132902 856
rect 133070 167 134190 856
rect 134358 167 135570 856
rect 135738 167 136950 856
rect 137118 167 138330 856
rect 138498 167 139710 856
rect 139878 167 141090 856
rect 141258 167 142378 856
rect 142546 167 143758 856
rect 143926 167 145138 856
rect 145306 167 146518 856
rect 146686 167 147898 856
rect 148066 167 149278 856
rect 149446 167 150566 856
rect 150734 167 151946 856
rect 152114 167 153326 856
rect 153494 167 154706 856
rect 154874 167 156086 856
rect 156254 167 157374 856
rect 157542 167 158754 856
rect 158922 167 160134 856
rect 160302 167 161514 856
rect 161682 167 162894 856
rect 163062 167 164274 856
rect 164442 167 165562 856
rect 165730 167 166942 856
rect 167110 167 168322 856
rect 168490 167 169702 856
rect 169870 167 171082 856
rect 171250 167 172462 856
rect 172630 167 173750 856
rect 173918 167 175130 856
rect 175298 167 176510 856
rect 176678 167 177890 856
rect 178058 167 179270 856
rect 179438 167 179564 856
<< metal3 >>
rect 0 119688 800 119808
rect 0 119416 800 119536
rect 0 119144 800 119264
rect 0 118872 800 118992
rect 0 118600 800 118720
rect 0 118328 800 118448
rect 0 118056 800 118176
rect 179200 118056 180000 118176
rect 0 117784 800 117904
rect 0 117376 800 117496
rect 0 117104 800 117224
rect 0 116832 800 116952
rect 0 116560 800 116680
rect 0 116288 800 116408
rect 0 116016 800 116136
rect 0 115744 800 115864
rect 0 115472 800 115592
rect 0 115064 800 115184
rect 0 114792 800 114912
rect 0 114520 800 114640
rect 179200 114520 180000 114640
rect 0 114248 800 114368
rect 0 113976 800 114096
rect 0 113704 800 113824
rect 0 113432 800 113552
rect 0 113160 800 113280
rect 0 112752 800 112872
rect 0 112480 800 112600
rect 0 112208 800 112328
rect 0 111936 800 112056
rect 0 111664 800 111784
rect 0 111392 800 111512
rect 0 111120 800 111240
rect 0 110848 800 110968
rect 179200 110984 180000 111104
rect 0 110576 800 110696
rect 0 110168 800 110288
rect 0 109896 800 110016
rect 0 109624 800 109744
rect 0 109352 800 109472
rect 0 109080 800 109200
rect 0 108808 800 108928
rect 0 108536 800 108656
rect 0 108264 800 108384
rect 0 107856 800 107976
rect 0 107584 800 107704
rect 0 107312 800 107432
rect 179200 107448 180000 107568
rect 0 107040 800 107160
rect 0 106768 800 106888
rect 0 106496 800 106616
rect 0 106224 800 106344
rect 0 105952 800 106072
rect 0 105544 800 105664
rect 0 105272 800 105392
rect 0 105000 800 105120
rect 0 104728 800 104848
rect 0 104456 800 104576
rect 0 104184 800 104304
rect 0 103912 800 104032
rect 179200 103912 180000 104032
rect 0 103640 800 103760
rect 0 103368 800 103488
rect 0 102960 800 103080
rect 0 102688 800 102808
rect 0 102416 800 102536
rect 0 102144 800 102264
rect 0 101872 800 101992
rect 0 101600 800 101720
rect 0 101328 800 101448
rect 0 101056 800 101176
rect 0 100648 800 100768
rect 0 100376 800 100496
rect 179200 100376 180000 100496
rect 0 100104 800 100224
rect 0 99832 800 99952
rect 0 99560 800 99680
rect 0 99288 800 99408
rect 0 99016 800 99136
rect 0 98744 800 98864
rect 0 98336 800 98456
rect 0 98064 800 98184
rect 0 97792 800 97912
rect 0 97520 800 97640
rect 0 97248 800 97368
rect 0 96976 800 97096
rect 0 96704 800 96824
rect 179200 96840 180000 96960
rect 0 96432 800 96552
rect 0 96160 800 96280
rect 0 95752 800 95872
rect 0 95480 800 95600
rect 0 95208 800 95328
rect 0 94936 800 95056
rect 0 94664 800 94784
rect 0 94392 800 94512
rect 0 94120 800 94240
rect 0 93848 800 93968
rect 0 93440 800 93560
rect 0 93168 800 93288
rect 179200 93304 180000 93424
rect 0 92896 800 93016
rect 0 92624 800 92744
rect 0 92352 800 92472
rect 0 92080 800 92200
rect 0 91808 800 91928
rect 0 91536 800 91656
rect 0 91128 800 91248
rect 0 90856 800 90976
rect 0 90584 800 90704
rect 0 90312 800 90432
rect 0 90040 800 90160
rect 0 89768 800 89888
rect 179200 89768 180000 89888
rect 0 89496 800 89616
rect 0 89224 800 89344
rect 0 88952 800 89072
rect 0 88544 800 88664
rect 0 88272 800 88392
rect 0 88000 800 88120
rect 0 87728 800 87848
rect 0 87456 800 87576
rect 0 87184 800 87304
rect 0 86912 800 87032
rect 0 86640 800 86760
rect 0 86232 800 86352
rect 179200 86232 180000 86352
rect 0 85960 800 86080
rect 0 85688 800 85808
rect 0 85416 800 85536
rect 0 85144 800 85264
rect 0 84872 800 84992
rect 0 84600 800 84720
rect 0 84328 800 84448
rect 0 83920 800 84040
rect 0 83648 800 83768
rect 0 83376 800 83496
rect 0 83104 800 83224
rect 0 82832 800 82952
rect 0 82560 800 82680
rect 179200 82696 180000 82816
rect 0 82288 800 82408
rect 0 82016 800 82136
rect 0 81744 800 81864
rect 0 81336 800 81456
rect 0 81064 800 81184
rect 0 80792 800 80912
rect 0 80520 800 80640
rect 0 80248 800 80368
rect 0 79976 800 80096
rect 0 79704 800 79824
rect 0 79432 800 79552
rect 0 79024 800 79144
rect 179200 79160 180000 79280
rect 0 78752 800 78872
rect 0 78480 800 78600
rect 0 78208 800 78328
rect 0 77936 800 78056
rect 0 77664 800 77784
rect 0 77392 800 77512
rect 0 77120 800 77240
rect 0 76712 800 76832
rect 0 76440 800 76560
rect 0 76168 800 76288
rect 0 75896 800 76016
rect 0 75624 800 75744
rect 179200 75624 180000 75744
rect 0 75352 800 75472
rect 0 75080 800 75200
rect 0 74808 800 74928
rect 0 74536 800 74656
rect 0 74128 800 74248
rect 0 73856 800 73976
rect 0 73584 800 73704
rect 0 73312 800 73432
rect 0 73040 800 73160
rect 0 72768 800 72888
rect 0 72496 800 72616
rect 0 72224 800 72344
rect 179200 72088 180000 72208
rect 0 71816 800 71936
rect 0 71544 800 71664
rect 0 71272 800 71392
rect 0 71000 800 71120
rect 0 70728 800 70848
rect 0 70456 800 70576
rect 0 70184 800 70304
rect 0 69912 800 70032
rect 0 69504 800 69624
rect 0 69232 800 69352
rect 0 68960 800 69080
rect 0 68688 800 68808
rect 0 68416 800 68536
rect 179200 68552 180000 68672
rect 0 68144 800 68264
rect 0 67872 800 67992
rect 0 67600 800 67720
rect 0 67328 800 67448
rect 0 66920 800 67040
rect 0 66648 800 66768
rect 0 66376 800 66496
rect 0 66104 800 66224
rect 0 65832 800 65952
rect 0 65560 800 65680
rect 0 65288 800 65408
rect 0 65016 800 65136
rect 179200 65016 180000 65136
rect 0 64608 800 64728
rect 0 64336 800 64456
rect 0 64064 800 64184
rect 0 63792 800 63912
rect 0 63520 800 63640
rect 0 63248 800 63368
rect 0 62976 800 63096
rect 0 62704 800 62824
rect 0 62296 800 62416
rect 0 62024 800 62144
rect 0 61752 800 61872
rect 0 61480 800 61600
rect 179200 61616 180000 61736
rect 0 61208 800 61328
rect 0 60936 800 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 0 59712 800 59832
rect 0 59440 800 59560
rect 0 59168 800 59288
rect 0 58896 800 59016
rect 0 58624 800 58744
rect 0 58352 800 58472
rect 0 58080 800 58200
rect 179200 58080 180000 58200
rect 0 57808 800 57928
rect 0 57400 800 57520
rect 0 57128 800 57248
rect 0 56856 800 56976
rect 0 56584 800 56704
rect 0 56312 800 56432
rect 0 56040 800 56160
rect 0 55768 800 55888
rect 0 55496 800 55616
rect 0 55088 800 55208
rect 0 54816 800 54936
rect 0 54544 800 54664
rect 179200 54544 180000 54664
rect 0 54272 800 54392
rect 0 54000 800 54120
rect 0 53728 800 53848
rect 0 53456 800 53576
rect 0 53184 800 53304
rect 0 52776 800 52896
rect 0 52504 800 52624
rect 0 52232 800 52352
rect 0 51960 800 52080
rect 0 51688 800 51808
rect 0 51416 800 51536
rect 0 51144 800 51264
rect 0 50872 800 50992
rect 179200 51008 180000 51128
rect 0 50600 800 50720
rect 0 50192 800 50312
rect 0 49920 800 50040
rect 0 49648 800 49768
rect 0 49376 800 49496
rect 0 49104 800 49224
rect 0 48832 800 48952
rect 0 48560 800 48680
rect 0 48288 800 48408
rect 0 47880 800 48000
rect 0 47608 800 47728
rect 0 47336 800 47456
rect 179200 47472 180000 47592
rect 0 47064 800 47184
rect 0 46792 800 46912
rect 0 46520 800 46640
rect 0 46248 800 46368
rect 0 45976 800 46096
rect 0 45568 800 45688
rect 0 45296 800 45416
rect 0 45024 800 45144
rect 0 44752 800 44872
rect 0 44480 800 44600
rect 0 44208 800 44328
rect 0 43936 800 44056
rect 179200 43936 180000 44056
rect 0 43664 800 43784
rect 0 43392 800 43512
rect 0 42984 800 43104
rect 0 42712 800 42832
rect 0 42440 800 42560
rect 0 42168 800 42288
rect 0 41896 800 42016
rect 0 41624 800 41744
rect 0 41352 800 41472
rect 0 41080 800 41200
rect 0 40672 800 40792
rect 0 40400 800 40520
rect 179200 40400 180000 40520
rect 0 40128 800 40248
rect 0 39856 800 39976
rect 0 39584 800 39704
rect 0 39312 800 39432
rect 0 39040 800 39160
rect 0 38768 800 38888
rect 0 38360 800 38480
rect 0 38088 800 38208
rect 0 37816 800 37936
rect 0 37544 800 37664
rect 0 37272 800 37392
rect 0 37000 800 37120
rect 0 36728 800 36848
rect 179200 36864 180000 36984
rect 0 36456 800 36576
rect 0 36184 800 36304
rect 0 35776 800 35896
rect 0 35504 800 35624
rect 0 35232 800 35352
rect 0 34960 800 35080
rect 0 34688 800 34808
rect 0 34416 800 34536
rect 0 34144 800 34264
rect 0 33872 800 33992
rect 0 33464 800 33584
rect 0 33192 800 33312
rect 179200 33328 180000 33448
rect 0 32920 800 33040
rect 0 32648 800 32768
rect 0 32376 800 32496
rect 0 32104 800 32224
rect 0 31832 800 31952
rect 0 31560 800 31680
rect 0 31152 800 31272
rect 0 30880 800 31000
rect 0 30608 800 30728
rect 0 30336 800 30456
rect 0 30064 800 30184
rect 0 29792 800 29912
rect 179200 29792 180000 29912
rect 0 29520 800 29640
rect 0 29248 800 29368
rect 0 28976 800 29096
rect 0 28568 800 28688
rect 0 28296 800 28416
rect 0 28024 800 28144
rect 0 27752 800 27872
rect 0 27480 800 27600
rect 0 27208 800 27328
rect 0 26936 800 27056
rect 0 26664 800 26784
rect 0 26256 800 26376
rect 179200 26256 180000 26376
rect 0 25984 800 26104
rect 0 25712 800 25832
rect 0 25440 800 25560
rect 0 25168 800 25288
rect 0 24896 800 25016
rect 0 24624 800 24744
rect 0 24352 800 24472
rect 0 23944 800 24064
rect 0 23672 800 23792
rect 0 23400 800 23520
rect 0 23128 800 23248
rect 0 22856 800 22976
rect 0 22584 800 22704
rect 179200 22720 180000 22840
rect 0 22312 800 22432
rect 0 22040 800 22160
rect 0 21768 800 21888
rect 0 21360 800 21480
rect 0 21088 800 21208
rect 0 20816 800 20936
rect 0 20544 800 20664
rect 0 20272 800 20392
rect 0 20000 800 20120
rect 0 19728 800 19848
rect 0 19456 800 19576
rect 0 19048 800 19168
rect 179200 19184 180000 19304
rect 0 18776 800 18896
rect 0 18504 800 18624
rect 0 18232 800 18352
rect 0 17960 800 18080
rect 0 17688 800 17808
rect 0 17416 800 17536
rect 0 17144 800 17264
rect 0 16736 800 16856
rect 0 16464 800 16584
rect 0 16192 800 16312
rect 0 15920 800 16040
rect 0 15648 800 15768
rect 179200 15648 180000 15768
rect 0 15376 800 15496
rect 0 15104 800 15224
rect 0 14832 800 14952
rect 0 14560 800 14680
rect 0 14152 800 14272
rect 0 13880 800 14000
rect 0 13608 800 13728
rect 0 13336 800 13456
rect 0 13064 800 13184
rect 0 12792 800 12912
rect 0 12520 800 12640
rect 0 12248 800 12368
rect 179200 12112 180000 12232
rect 0 11840 800 11960
rect 0 11568 800 11688
rect 0 11296 800 11416
rect 0 11024 800 11144
rect 0 10752 800 10872
rect 0 10480 800 10600
rect 0 10208 800 10328
rect 0 9936 800 10056
rect 0 9528 800 9648
rect 0 9256 800 9376
rect 0 8984 800 9104
rect 0 8712 800 8832
rect 0 8440 800 8560
rect 179200 8576 180000 8696
rect 0 8168 800 8288
rect 0 7896 800 8016
rect 0 7624 800 7744
rect 0 7352 800 7472
rect 0 6944 800 7064
rect 0 6672 800 6792
rect 0 6400 800 6520
rect 0 6128 800 6248
rect 0 5856 800 5976
rect 0 5584 800 5704
rect 0 5312 800 5432
rect 0 5040 800 5160
rect 179200 5040 180000 5160
rect 0 4632 800 4752
rect 0 4360 800 4480
rect 0 4088 800 4208
rect 0 3816 800 3936
rect 0 3544 800 3664
rect 0 3272 800 3392
rect 0 3000 800 3120
rect 0 2728 800 2848
rect 0 2320 800 2440
rect 0 2048 800 2168
rect 0 1776 800 1896
rect 0 1504 800 1624
rect 179200 1640 180000 1760
rect 0 1232 800 1352
rect 0 960 800 1080
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
<< obsm3 >>
rect 880 118256 179200 119781
rect 880 117976 179120 118256
rect 880 117704 179200 117976
rect 800 117576 179200 117704
rect 880 115392 179200 117576
rect 800 115264 179200 115392
rect 880 114720 179200 115264
rect 880 114440 179120 114720
rect 880 113080 179200 114440
rect 800 112952 179200 113080
rect 880 111184 179200 112952
rect 880 110904 179120 111184
rect 880 110496 179200 110904
rect 800 110368 179200 110496
rect 880 108184 179200 110368
rect 800 108056 179200 108184
rect 880 107648 179200 108056
rect 880 107368 179120 107648
rect 880 105872 179200 107368
rect 800 105744 179200 105872
rect 880 104112 179200 105744
rect 880 103832 179120 104112
rect 880 103288 179200 103832
rect 800 103160 179200 103288
rect 880 100976 179200 103160
rect 800 100848 179200 100976
rect 880 100576 179200 100848
rect 880 100296 179120 100576
rect 880 98664 179200 100296
rect 800 98536 179200 98664
rect 880 97040 179200 98536
rect 880 96760 179120 97040
rect 880 96080 179200 96760
rect 800 95952 179200 96080
rect 880 93768 179200 95952
rect 800 93640 179200 93768
rect 880 93504 179200 93640
rect 880 93224 179120 93504
rect 880 91456 179200 93224
rect 800 91328 179200 91456
rect 880 89968 179200 91328
rect 880 89688 179120 89968
rect 880 88872 179200 89688
rect 800 88744 179200 88872
rect 880 86560 179200 88744
rect 800 86432 179200 86560
rect 880 86152 179120 86432
rect 880 84248 179200 86152
rect 800 84120 179200 84248
rect 880 82896 179200 84120
rect 880 82616 179120 82896
rect 880 81664 179200 82616
rect 800 81536 179200 81664
rect 880 79360 179200 81536
rect 880 79352 179120 79360
rect 800 79224 179120 79352
rect 880 79080 179120 79224
rect 880 77040 179200 79080
rect 800 76912 179200 77040
rect 880 75824 179200 76912
rect 880 75544 179120 75824
rect 880 74456 179200 75544
rect 800 74328 179200 74456
rect 880 72288 179200 74328
rect 880 72144 179120 72288
rect 800 72016 179120 72144
rect 880 72008 179120 72016
rect 880 69832 179200 72008
rect 800 69704 179200 69832
rect 880 68752 179200 69704
rect 880 68472 179120 68752
rect 880 67248 179200 68472
rect 800 67120 179200 67248
rect 880 65216 179200 67120
rect 880 64936 179120 65216
rect 800 64808 179200 64936
rect 880 62624 179200 64808
rect 800 62496 179200 62624
rect 880 61816 179200 62496
rect 880 61536 179120 61816
rect 880 60040 179200 61536
rect 800 59912 179200 60040
rect 880 58280 179200 59912
rect 880 58000 179120 58280
rect 880 57728 179200 58000
rect 800 57600 179200 57728
rect 880 55416 179200 57600
rect 800 55288 179200 55416
rect 880 54744 179200 55288
rect 880 54464 179120 54744
rect 880 53104 179200 54464
rect 800 52976 179200 53104
rect 880 51208 179200 52976
rect 880 50928 179120 51208
rect 880 50520 179200 50928
rect 800 50392 179200 50520
rect 880 48208 179200 50392
rect 800 48080 179200 48208
rect 880 47672 179200 48080
rect 880 47392 179120 47672
rect 880 45896 179200 47392
rect 800 45768 179200 45896
rect 880 44136 179200 45768
rect 880 43856 179120 44136
rect 880 43312 179200 43856
rect 800 43184 179200 43312
rect 880 41000 179200 43184
rect 800 40872 179200 41000
rect 880 40600 179200 40872
rect 880 40320 179120 40600
rect 880 38688 179200 40320
rect 800 38560 179200 38688
rect 880 37064 179200 38560
rect 880 36784 179120 37064
rect 880 36104 179200 36784
rect 800 35976 179200 36104
rect 880 33792 179200 35976
rect 800 33664 179200 33792
rect 880 33528 179200 33664
rect 880 33248 179120 33528
rect 880 31480 179200 33248
rect 800 31352 179200 31480
rect 880 29992 179200 31352
rect 880 29712 179120 29992
rect 880 28896 179200 29712
rect 800 28768 179200 28896
rect 880 26584 179200 28768
rect 800 26456 179200 26584
rect 880 26176 179120 26456
rect 880 24272 179200 26176
rect 800 24144 179200 24272
rect 880 22920 179200 24144
rect 880 22640 179120 22920
rect 880 21688 179200 22640
rect 800 21560 179200 21688
rect 880 19384 179200 21560
rect 880 19376 179120 19384
rect 800 19248 179120 19376
rect 880 19104 179120 19248
rect 880 17064 179200 19104
rect 800 16936 179200 17064
rect 880 15848 179200 16936
rect 880 15568 179120 15848
rect 880 14480 179200 15568
rect 800 14352 179200 14480
rect 880 12312 179200 14352
rect 880 12168 179120 12312
rect 800 12040 179120 12168
rect 880 12032 179120 12040
rect 880 9856 179200 12032
rect 800 9728 179200 9856
rect 880 8776 179200 9728
rect 880 8496 179120 8776
rect 880 7272 179200 8496
rect 800 7144 179200 7272
rect 880 5240 179200 7144
rect 880 4960 179120 5240
rect 800 4832 179200 4960
rect 880 2648 179200 4832
rect 800 2520 179200 2648
rect 880 1840 179200 2520
rect 880 1560 179120 1840
rect 880 171 179200 1560
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 106227 46683 106293 48245
<< labels >>
rlabel metal2 s 478 119200 534 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 29918 119200 29974 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 32862 119200 32918 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 35806 119200 35862 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 38842 119200 38898 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 41786 119200 41842 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 44730 119200 44786 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 47674 119200 47730 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 50618 119200 50674 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 53562 119200 53618 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 56506 119200 56562 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 3422 119200 3478 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 59450 119200 59506 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 62394 119200 62450 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 65338 119200 65394 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 68282 119200 68338 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 71226 119200 71282 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 74262 119200 74318 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 77206 119200 77262 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 80150 119200 80206 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 83094 119200 83150 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 86038 119200 86094 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 6366 119200 6422 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 88982 119200 89038 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 91926 119200 91982 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 94870 119200 94926 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 97814 119200 97870 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 100758 119200 100814 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 103702 119200 103758 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 106646 119200 106702 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 109682 119200 109738 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 9310 119200 9366 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 12254 119200 12310 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 15198 119200 15254 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 18142 119200 18198 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 21086 119200 21142 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 24030 119200 24086 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 26974 119200 27030 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 1398 119200 1454 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 30930 119200 30986 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 33874 119200 33930 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 36818 119200 36874 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 39762 119200 39818 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 42706 119200 42762 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 45650 119200 45706 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 48686 119200 48742 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 51630 119200 51686 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 54574 119200 54630 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 57518 119200 57574 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 4342 119200 4398 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 60462 119200 60518 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 63406 119200 63462 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 66350 119200 66406 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 69294 119200 69350 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 72238 119200 72294 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 75182 119200 75238 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 78126 119200 78182 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 81070 119200 81126 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 84014 119200 84070 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 7286 119200 7342 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 89994 119200 90050 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 92938 119200 92994 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 95882 119200 95938 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 98826 119200 98882 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 101770 119200 101826 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 104714 119200 104770 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 107658 119200 107714 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 110602 119200 110658 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 10230 119200 10286 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 13266 119200 13322 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 16210 119200 16266 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 19154 119200 19210 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 22098 119200 22154 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 25042 119200 25098 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 27986 119200 28042 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 2410 119200 2466 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 31942 119200 31998 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 34886 119200 34942 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 37830 119200 37886 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 40774 119200 40830 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 43718 119200 43774 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 46662 119200 46718 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 49606 119200 49662 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 52550 119200 52606 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 55494 119200 55550 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 58438 119200 58494 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 5354 119200 5410 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 61474 119200 61530 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 64418 119200 64474 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 67362 119200 67418 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 70306 119200 70362 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 73250 119200 73306 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 76194 119200 76250 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 79138 119200 79194 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 82082 119200 82138 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 85026 119200 85082 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 87970 119200 88026 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 8298 119200 8354 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 90914 119200 90970 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 93858 119200 93914 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 96894 119200 96950 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 99838 119200 99894 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 102782 119200 102838 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 105726 119200 105782 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 108670 119200 108726 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 111614 119200 111670 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 11242 119200 11298 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 14186 119200 14242 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 17130 119200 17186 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 20074 119200 20130 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 23018 119200 23074 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 26054 119200 26110 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 145102 119200 145158 120000 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 150622 0 150678 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 149978 119200 150034 120000 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 0 144 800 264 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 la_data_in[100]
port 119 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 la_data_in[101]
port 120 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 0 89224 800 89344 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 la_data_in[106]
port 125 nsew signal input
rlabel metal3 s 0 92624 800 92744 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 0 93440 800 93560 6 la_data_in[108]
port 127 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 8712 800 8832 6 la_data_in[10]
port 129 nsew signal input
rlabel metal3 s 0 95208 800 95328 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 0 96160 800 96280 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 96976 800 97096 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 0 97792 800 97912 6 la_data_in[113]
port 133 nsew signal input
rlabel metal3 s 0 98744 800 98864 6 la_data_in[114]
port 134 nsew signal input
rlabel metal3 s 0 99560 800 99680 6 la_data_in[115]
port 135 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 la_data_in[116]
port 136 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 la_data_in[117]
port 137 nsew signal input
rlabel metal3 s 0 102144 800 102264 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 0 102960 800 103080 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 9528 800 9648 6 la_data_in[11]
port 140 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 la_data_in[120]
port 141 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_data_in[121]
port 142 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 la_data_in[122]
port 143 nsew signal input
rlabel metal3 s 0 106496 800 106616 6 la_data_in[123]
port 144 nsew signal input
rlabel metal3 s 0 107312 800 107432 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 la_data_in[125]
port 146 nsew signal input
rlabel metal3 s 0 109080 800 109200 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 10480 800 10600 6 la_data_in[12]
port 149 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 13064 800 13184 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 14832 800 14952 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_data_in[18]
port 155 nsew signal input
rlabel metal3 s 0 16464 800 16584 6 la_data_in[19]
port 156 nsew signal input
rlabel metal3 s 0 960 800 1080 6 la_data_in[1]
port 157 nsew signal input
rlabel metal3 s 0 17416 800 17536 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 18232 800 18352 6 la_data_in[21]
port 159 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 0 20000 800 20120 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 0 20816 800 20936 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 0 24352 800 24472 6 la_data_in[28]
port 166 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 la_data_in[29]
port 167 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 la_data_in[2]
port 168 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 la_data_in[30]
port 169 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 la_data_in[31]
port 170 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 la_data_in[32]
port 171 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 la_data_in[33]
port 172 nsew signal input
rlabel metal3 s 0 29520 800 29640 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 0 30336 800 30456 6 la_data_in[35]
port 174 nsew signal input
rlabel metal3 s 0 31152 800 31272 6 la_data_in[36]
port 175 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 la_data_in[38]
port 177 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 la_data_in[3]
port 179 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 la_data_in[40]
port 180 nsew signal input
rlabel metal3 s 0 35504 800 35624 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 la_data_in[43]
port 183 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 39040 800 39160 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 39856 800 39976 6 la_data_in[46]
port 186 nsew signal input
rlabel metal3 s 0 40672 800 40792 6 la_data_in[47]
port 187 nsew signal input
rlabel metal3 s 0 41624 800 41744 6 la_data_in[48]
port 188 nsew signal input
rlabel metal3 s 0 42440 800 42560 6 la_data_in[49]
port 189 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 43392 800 43512 6 la_data_in[50]
port 191 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 la_data_in[51]
port 192 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 la_data_in[53]
port 194 nsew signal input
rlabel metal3 s 0 46792 800 46912 6 la_data_in[54]
port 195 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 la_data_in[55]
port 196 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 la_data_in[56]
port 197 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 la_data_in[57]
port 198 nsew signal input
rlabel metal3 s 0 50192 800 50312 6 la_data_in[58]
port 199 nsew signal input
rlabel metal3 s 0 51144 800 51264 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 4360 800 4480 6 la_data_in[5]
port 201 nsew signal input
rlabel metal3 s 0 51960 800 52080 6 la_data_in[60]
port 202 nsew signal input
rlabel metal3 s 0 52776 800 52896 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 0 53728 800 53848 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 54544 800 54664 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 0 55496 800 55616 6 la_data_in[64]
port 206 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 0 57128 800 57248 6 la_data_in[66]
port 208 nsew signal input
rlabel metal3 s 0 58080 800 58200 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 58896 800 59016 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 0 5312 800 5432 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 la_data_in[71]
port 214 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 la_data_in[72]
port 215 nsew signal input
rlabel metal3 s 0 63248 800 63368 6 la_data_in[73]
port 216 nsew signal input
rlabel metal3 s 0 64064 800 64184 6 la_data_in[74]
port 217 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 la_data_in[75]
port 218 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 0 68416 800 68536 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 la_data_in[7]
port 223 nsew signal input
rlabel metal3 s 0 69232 800 69352 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 la_data_in[82]
port 226 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 72768 800 72888 6 la_data_in[84]
port 228 nsew signal input
rlabel metal3 s 0 73584 800 73704 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 la_data_in[88]
port 232 nsew signal input
rlabel metal3 s 0 77120 800 77240 6 la_data_in[89]
port 233 nsew signal input
rlabel metal3 s 0 6944 800 7064 6 la_data_in[8]
port 234 nsew signal input
rlabel metal3 s 0 77936 800 78056 6 la_data_in[90]
port 235 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 la_data_in[92]
port 237 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 la_data_in[93]
port 238 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 0 84872 800 84992 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 85688 800 85808 6 la_data_in[99]
port 244 nsew signal input
rlabel metal3 s 0 7896 800 8016 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 416 800 536 6 la_data_out[0]
port 246 nsew signal output
rlabel metal3 s 0 86912 800 87032 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 0 87728 800 87848 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 0 89496 800 89616 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 91128 800 91248 6 la_data_out[105]
port 252 nsew signal output
rlabel metal3 s 0 92080 800 92200 6 la_data_out[106]
port 253 nsew signal output
rlabel metal3 s 0 92896 800 93016 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 0 93848 800 93968 6 la_data_out[108]
port 255 nsew signal output
rlabel metal3 s 0 94664 800 94784 6 la_data_out[109]
port 256 nsew signal output
rlabel metal3 s 0 8984 800 9104 6 la_data_out[10]
port 257 nsew signal output
rlabel metal3 s 0 95480 800 95600 6 la_data_out[110]
port 258 nsew signal output
rlabel metal3 s 0 96432 800 96552 6 la_data_out[111]
port 259 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 la_data_out[113]
port 261 nsew signal output
rlabel metal3 s 0 99016 800 99136 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 0 99832 800 99952 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 la_data_out[117]
port 265 nsew signal output
rlabel metal3 s 0 102416 800 102536 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 103368 800 103488 6 la_data_out[119]
port 267 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 0 104184 800 104304 6 la_data_out[120]
port 269 nsew signal output
rlabel metal3 s 0 105000 800 105120 6 la_data_out[121]
port 270 nsew signal output
rlabel metal3 s 0 105952 800 106072 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 0 106768 800 106888 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 107584 800 107704 6 la_data_out[124]
port 273 nsew signal output
rlabel metal3 s 0 108536 800 108656 6 la_data_out[125]
port 274 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 110168 800 110288 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 0 13336 800 13456 6 la_data_out[15]
port 280 nsew signal output
rlabel metal3 s 0 14152 800 14272 6 la_data_out[16]
port 281 nsew signal output
rlabel metal3 s 0 15104 800 15224 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 0 15920 800 16040 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 16736 800 16856 6 la_data_out[19]
port 284 nsew signal output
rlabel metal3 s 0 1232 800 1352 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 0 17688 800 17808 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 18504 800 18624 6 la_data_out[21]
port 287 nsew signal output
rlabel metal3 s 0 19456 800 19576 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 0 20272 800 20392 6 la_data_out[23]
port 289 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 la_data_out[24]
port 290 nsew signal output
rlabel metal3 s 0 22040 800 22160 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 0 23672 800 23792 6 la_data_out[27]
port 293 nsew signal output
rlabel metal3 s 0 24624 800 24744 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 0 25440 800 25560 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 0 2048 800 2168 6 la_data_out[2]
port 296 nsew signal output
rlabel metal3 s 0 26256 800 26376 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 la_data_out[31]
port 298 nsew signal output
rlabel metal3 s 0 28024 800 28144 6 la_data_out[32]
port 299 nsew signal output
rlabel metal3 s 0 28976 800 29096 6 la_data_out[33]
port 300 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 la_data_out[34]
port 301 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 31560 800 31680 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 la_data_out[37]
port 304 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 la_data_out[39]
port 306 nsew signal output
rlabel metal3 s 0 3000 800 3120 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 34960 800 35080 6 la_data_out[40]
port 308 nsew signal output
rlabel metal3 s 0 35776 800 35896 6 la_data_out[41]
port 309 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 la_data_out[42]
port 310 nsew signal output
rlabel metal3 s 0 37544 800 37664 6 la_data_out[43]
port 311 nsew signal output
rlabel metal3 s 0 38360 800 38480 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 0 39312 800 39432 6 la_data_out[45]
port 313 nsew signal output
rlabel metal3 s 0 40128 800 40248 6 la_data_out[46]
port 314 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 la_data_out[48]
port 316 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 3816 800 3936 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 43664 800 43784 6 la_data_out[50]
port 319 nsew signal output
rlabel metal3 s 0 44480 800 44600 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 45296 800 45416 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 48832 800 48952 6 la_data_out[56]
port 325 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 la_data_out[57]
port 326 nsew signal output
rlabel metal3 s 0 50600 800 50720 6 la_data_out[58]
port 327 nsew signal output
rlabel metal3 s 0 51416 800 51536 6 la_data_out[59]
port 328 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 la_data_out[5]
port 329 nsew signal output
rlabel metal3 s 0 52232 800 52352 6 la_data_out[60]
port 330 nsew signal output
rlabel metal3 s 0 53184 800 53304 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 0 54000 800 54120 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 0 54816 800 54936 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 la_data_out[65]
port 335 nsew signal output
rlabel metal3 s 0 57400 800 57520 6 la_data_out[66]
port 336 nsew signal output
rlabel metal3 s 0 58352 800 58472 6 la_data_out[67]
port 337 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 la_data_out[68]
port 338 nsew signal output
rlabel metal3 s 0 60120 800 60240 6 la_data_out[69]
port 339 nsew signal output
rlabel metal3 s 0 5584 800 5704 6 la_data_out[6]
port 340 nsew signal output
rlabel metal3 s 0 60936 800 61056 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 0 61752 800 61872 6 la_data_out[71]
port 342 nsew signal output
rlabel metal3 s 0 62704 800 62824 6 la_data_out[72]
port 343 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 la_data_out[73]
port 344 nsew signal output
rlabel metal3 s 0 64336 800 64456 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 0 65288 800 65408 6 la_data_out[75]
port 346 nsew signal output
rlabel metal3 s 0 66104 800 66224 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 0 66920 800 67040 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 la_data_out[78]
port 349 nsew signal output
rlabel metal3 s 0 68688 800 68808 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 0 6400 800 6520 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 69504 800 69624 6 la_data_out[80]
port 352 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 la_data_out[81]
port 353 nsew signal output
rlabel metal3 s 0 71272 800 71392 6 la_data_out[82]
port 354 nsew signal output
rlabel metal3 s 0 72224 800 72344 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 73040 800 73160 6 la_data_out[84]
port 356 nsew signal output
rlabel metal3 s 0 73856 800 73976 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 0 74808 800 74928 6 la_data_out[86]
port 358 nsew signal output
rlabel metal3 s 0 75624 800 75744 6 la_data_out[87]
port 359 nsew signal output
rlabel metal3 s 0 76440 800 76560 6 la_data_out[88]
port 360 nsew signal output
rlabel metal3 s 0 77392 800 77512 6 la_data_out[89]
port 361 nsew signal output
rlabel metal3 s 0 7352 800 7472 6 la_data_out[8]
port 362 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 la_data_out[90]
port 363 nsew signal output
rlabel metal3 s 0 79024 800 79144 6 la_data_out[91]
port 364 nsew signal output
rlabel metal3 s 0 79976 800 80096 6 la_data_out[92]
port 365 nsew signal output
rlabel metal3 s 0 80792 800 80912 6 la_data_out[93]
port 366 nsew signal output
rlabel metal3 s 0 81744 800 81864 6 la_data_out[94]
port 367 nsew signal output
rlabel metal3 s 0 82560 800 82680 6 la_data_out[95]
port 368 nsew signal output
rlabel metal3 s 0 83376 800 83496 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 la_data_out[97]
port 370 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 la_data_out[98]
port 371 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 la_data_out[99]
port 372 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 la_data_out[9]
port 373 nsew signal output
rlabel metal3 s 0 688 800 808 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 la_oenb[101]
port 376 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 la_oenb[102]
port 377 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 0 90584 800 90704 6 la_oenb[104]
port 379 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 la_oenb[105]
port 380 nsew signal input
rlabel metal3 s 0 92352 800 92472 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 la_oenb[107]
port 382 nsew signal input
rlabel metal3 s 0 94120 800 94240 6 la_oenb[108]
port 383 nsew signal input
rlabel metal3 s 0 94936 800 95056 6 la_oenb[109]
port 384 nsew signal input
rlabel metal3 s 0 9256 800 9376 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 0 95752 800 95872 6 la_oenb[110]
port 386 nsew signal input
rlabel metal3 s 0 96704 800 96824 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 la_oenb[112]
port 388 nsew signal input
rlabel metal3 s 0 98336 800 98456 6 la_oenb[113]
port 389 nsew signal input
rlabel metal3 s 0 99288 800 99408 6 la_oenb[114]
port 390 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 la_oenb[115]
port 391 nsew signal input
rlabel metal3 s 0 101056 800 101176 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 0 101872 800 101992 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 0 102688 800 102808 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 la_oenb[11]
port 396 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 la_oenb[120]
port 397 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 106224 800 106344 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 0 107040 800 107160 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 107856 800 107976 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 la_oenb[125]
port 402 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 0 110576 800 110696 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 11840 800 11960 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 12792 800 12912 6 la_oenb[14]
port 407 nsew signal input
rlabel metal3 s 0 13608 800 13728 6 la_oenb[15]
port 408 nsew signal input
rlabel metal3 s 0 14560 800 14680 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 la_oenb[17]
port 410 nsew signal input
rlabel metal3 s 0 16192 800 16312 6 la_oenb[18]
port 411 nsew signal input
rlabel metal3 s 0 17144 800 17264 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 0 17960 800 18080 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 la_oenb[21]
port 415 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 20544 800 20664 6 la_oenb[23]
port 417 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 la_oenb[24]
port 418 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 la_oenb[25]
port 419 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 la_oenb[27]
port 421 nsew signal input
rlabel metal3 s 0 24896 800 25016 6 la_oenb[28]
port 422 nsew signal input
rlabel metal3 s 0 25712 800 25832 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 2320 800 2440 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 la_oenb[30]
port 425 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 la_oenb[31]
port 426 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 la_oenb[32]
port 427 nsew signal input
rlabel metal3 s 0 29248 800 29368 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 0 30880 800 31000 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 la_oenb[36]
port 431 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 la_oenb[39]
port 434 nsew signal input
rlabel metal3 s 0 3272 800 3392 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 la_oenb[40]
port 436 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 la_oenb[41]
port 437 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 la_oenb[44]
port 440 nsew signal input
rlabel metal3 s 0 39584 800 39704 6 la_oenb[45]
port 441 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 la_oenb[46]
port 442 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 0 42168 800 42288 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 0 42984 800 43104 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 la_oenb[4]
port 446 nsew signal input
rlabel metal3 s 0 43936 800 44056 6 la_oenb[50]
port 447 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 0 46520 800 46640 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 47336 800 47456 6 la_oenb[54]
port 451 nsew signal input
rlabel metal3 s 0 48288 800 48408 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 49104 800 49224 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 0 49920 800 50040 6 la_oenb[57]
port 454 nsew signal input
rlabel metal3 s 0 50872 800 50992 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 la_oenb[59]
port 456 nsew signal input
rlabel metal3 s 0 5040 800 5160 6 la_oenb[5]
port 457 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 la_oenb[60]
port 458 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 la_oenb[61]
port 459 nsew signal input
rlabel metal3 s 0 54272 800 54392 6 la_oenb[62]
port 460 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 la_oenb[63]
port 461 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 la_oenb[64]
port 462 nsew signal input
rlabel metal3 s 0 56856 800 56976 6 la_oenb[65]
port 463 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 58624 800 58744 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 0 59440 800 59560 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 5856 800 5976 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 62976 800 63096 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 la_oenb[73]
port 472 nsew signal input
rlabel metal3 s 0 64608 800 64728 6 la_oenb[74]
port 473 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 la_oenb[75]
port 474 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 0 67328 800 67448 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 0 68960 800 69080 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 la_oenb[82]
port 482 nsew signal input
rlabel metal3 s 0 72496 800 72616 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 0 73312 800 73432 6 la_oenb[84]
port 484 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 la_oenb[87]
port 487 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 la_oenb[8]
port 490 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 la_oenb[91]
port 492 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 la_oenb[93]
port 494 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 0 82832 800 82952 6 la_oenb[95]
port 496 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 la_oenb[96]
port 497 nsew signal input
rlabel metal3 s 0 84600 800 84720 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 la_oenb[99]
port 500 nsew signal input
rlabel metal3 s 0 8440 800 8560 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 mem_data2_i[0]
port 502 nsew signal input
rlabel metal2 s 161754 119200 161810 120000 6 mem_data2_i[10]
port 503 nsew signal input
rlabel metal3 s 179200 61616 180000 61736 6 mem_data2_i[11]
port 504 nsew signal input
rlabel metal2 s 166998 0 167054 800 6 mem_data2_i[12]
port 505 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 mem_data2_i[13]
port 506 nsew signal input
rlabel metal3 s 179200 68552 180000 68672 6 mem_data2_i[14]
port 507 nsew signal input
rlabel metal3 s 0 116016 800 116136 6 mem_data2_i[15]
port 508 nsew signal input
rlabel metal2 s 171138 0 171194 800 6 mem_data2_i[16]
port 509 nsew signal input
rlabel metal3 s 179200 75624 180000 75744 6 mem_data2_i[17]
port 510 nsew signal input
rlabel metal3 s 179200 82696 180000 82816 6 mem_data2_i[18]
port 511 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 mem_data2_i[19]
port 512 nsew signal input
rlabel metal2 s 148966 119200 149022 120000 6 mem_data2_i[1]
port 513 nsew signal input
rlabel metal3 s 179200 86232 180000 86352 6 mem_data2_i[20]
port 514 nsew signal input
rlabel metal3 s 0 117376 800 117496 6 mem_data2_i[21]
port 515 nsew signal input
rlabel metal2 s 176566 0 176622 800 6 mem_data2_i[22]
port 516 nsew signal input
rlabel metal3 s 179200 89768 180000 89888 6 mem_data2_i[23]
port 517 nsew signal input
rlabel metal3 s 179200 93304 180000 93424 6 mem_data2_i[24]
port 518 nsew signal input
rlabel metal3 s 0 118328 800 118448 6 mem_data2_i[25]
port 519 nsew signal input
rlabel metal2 s 175554 119200 175610 120000 6 mem_data2_i[26]
port 520 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 mem_data2_i[27]
port 521 nsew signal input
rlabel metal3 s 179200 100376 180000 100496 6 mem_data2_i[28]
port 522 nsew signal input
rlabel metal3 s 0 119416 800 119536 6 mem_data2_i[29]
port 523 nsew signal input
rlabel metal2 s 150990 119200 151046 120000 6 mem_data2_i[2]
port 524 nsew signal input
rlabel metal2 s 176566 119200 176622 120000 6 mem_data2_i[30]
port 525 nsew signal input
rlabel metal2 s 178498 119200 178554 120000 6 mem_data2_i[31]
port 526 nsew signal input
rlabel metal3 s 0 111936 800 112056 6 mem_data2_i[3]
port 527 nsew signal input
rlabel metal2 s 153934 119200 153990 120000 6 mem_data2_i[4]
port 528 nsew signal input
rlabel metal3 s 179200 36864 180000 36984 6 mem_data2_i[5]
port 529 nsew signal input
rlabel metal3 s 0 112752 800 112872 6 mem_data2_i[6]
port 530 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 mem_data2_i[7]
port 531 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 mem_data2_i[8]
port 532 nsew signal input
rlabel metal2 s 164330 0 164386 800 6 mem_data2_i[9]
port 533 nsew signal input
rlabel metal2 s 146022 119200 146078 120000 6 mem_data_i[0]
port 534 nsew signal input
rlabel metal3 s 0 114248 800 114368 6 mem_data_i[10]
port 535 nsew signal input
rlabel metal2 s 162766 119200 162822 120000 6 mem_data_i[11]
port 536 nsew signal input
rlabel metal3 s 179200 65016 180000 65136 6 mem_data_i[12]
port 537 nsew signal input
rlabel metal2 s 163778 119200 163834 120000 6 mem_data_i[13]
port 538 nsew signal input
rlabel metal3 s 0 115472 800 115592 6 mem_data_i[14]
port 539 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 mem_data_i[15]
port 540 nsew signal input
rlabel metal3 s 0 116560 800 116680 6 mem_data_i[16]
port 541 nsew signal input
rlabel metal3 s 179200 79160 180000 79280 6 mem_data_i[17]
port 542 nsew signal input
rlabel metal2 s 166722 119200 166778 120000 6 mem_data_i[18]
port 543 nsew signal input
rlabel metal2 s 173806 0 173862 800 6 mem_data_i[19]
port 544 nsew signal input
rlabel metal3 s 0 110848 800 110968 6 mem_data_i[1]
port 545 nsew signal input
rlabel metal3 s 0 116832 800 116952 6 mem_data_i[20]
port 546 nsew signal input
rlabel metal2 s 168654 119200 168710 120000 6 mem_data_i[21]
port 547 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 mem_data_i[22]
port 548 nsew signal input
rlabel metal2 s 171598 119200 171654 120000 6 mem_data_i[23]
port 549 nsew signal input
rlabel metal2 s 172610 119200 172666 120000 6 mem_data_i[24]
port 550 nsew signal input
rlabel metal2 s 174542 119200 174598 120000 6 mem_data_i[25]
port 551 nsew signal input
rlabel metal3 s 0 118600 800 118720 6 mem_data_i[26]
port 552 nsew signal input
rlabel metal3 s 179200 96840 180000 96960 6 mem_data_i[27]
port 553 nsew signal input
rlabel metal3 s 179200 103912 180000 104032 6 mem_data_i[28]
port 554 nsew signal input
rlabel metal3 s 179200 110984 180000 111104 6 mem_data_i[29]
port 555 nsew signal input
rlabel metal3 s 0 111664 800 111784 6 mem_data_i[2]
port 556 nsew signal input
rlabel metal3 s 179200 118056 180000 118176 6 mem_data_i[30]
port 557 nsew signal input
rlabel metal2 s 179510 119200 179566 120000 6 mem_data_i[31]
port 558 nsew signal input
rlabel metal2 s 154762 0 154818 800 6 mem_data_i[3]
port 559 nsew signal input
rlabel metal3 s 179200 29792 180000 29912 6 mem_data_i[4]
port 560 nsew signal input
rlabel metal2 s 155866 119200 155922 120000 6 mem_data_i[5]
port 561 nsew signal input
rlabel metal2 s 160190 0 160246 800 6 mem_data_i[6]
port 562 nsew signal input
rlabel metal3 s 179200 51008 180000 51128 6 mem_data_i[7]
port 563 nsew signal input
rlabel metal2 s 161570 0 161626 800 6 mem_data_i[8]
port 564 nsew signal input
rlabel metal3 s 179200 58080 180000 58200 6 mem_data_i[9]
port 565 nsew signal input
rlabel metal2 s 147034 119200 147090 120000 6 mem_data_o[0]
port 566 nsew signal output
rlabel metal3 s 0 114520 800 114640 6 mem_data_o[10]
port 567 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 mem_data_o[11]
port 568 nsew signal output
rlabel metal2 s 168378 0 168434 800 6 mem_data_o[12]
port 569 nsew signal output
rlabel metal2 s 169758 0 169814 800 6 mem_data_o[13]
port 570 nsew signal output
rlabel metal3 s 0 115744 800 115864 6 mem_data_o[14]
port 571 nsew signal output
rlabel metal3 s 179200 72088 180000 72208 6 mem_data_o[15]
port 572 nsew signal output
rlabel metal2 s 164698 119200 164754 120000 6 mem_data_o[16]
port 573 nsew signal output
rlabel metal2 s 165710 119200 165766 120000 6 mem_data_o[17]
port 574 nsew signal output
rlabel metal2 s 167642 119200 167698 120000 6 mem_data_o[18]
port 575 nsew signal output
rlabel metal2 s 175186 0 175242 800 6 mem_data_o[19]
port 576 nsew signal output
rlabel metal3 s 179200 8576 180000 8696 6 mem_data_o[1]
port 577 nsew signal output
rlabel metal3 s 0 117104 800 117224 6 mem_data_o[20]
port 578 nsew signal output
rlabel metal2 s 169666 119200 169722 120000 6 mem_data_o[21]
port 579 nsew signal output
rlabel metal2 s 170678 119200 170734 120000 6 mem_data_o[22]
port 580 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 mem_data_o[23]
port 581 nsew signal output
rlabel metal2 s 173622 119200 173678 120000 6 mem_data_o[24]
port 582 nsew signal output
rlabel metal2 s 177946 0 178002 800 6 mem_data_o[25]
port 583 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 mem_data_o[26]
port 584 nsew signal output
rlabel metal2 s 179326 0 179382 800 6 mem_data_o[27]
port 585 nsew signal output
rlabel metal3 s 179200 107448 180000 107568 6 mem_data_o[28]
port 586 nsew signal output
rlabel metal3 s 179200 114520 180000 114640 6 mem_data_o[29]
port 587 nsew signal output
rlabel metal2 s 151910 119200 151966 120000 6 mem_data_o[2]
port 588 nsew signal output
rlabel metal2 s 177486 119200 177542 120000 6 mem_data_o[30]
port 589 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 mem_data_o[31]
port 590 nsew signal output
rlabel metal2 s 156142 0 156198 800 6 mem_data_o[3]
port 591 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 mem_data_o[4]
port 592 nsew signal output
rlabel metal2 s 158810 0 158866 800 6 mem_data_o[5]
port 593 nsew signal output
rlabel metal3 s 179200 40400 180000 40520 6 mem_data_o[6]
port 594 nsew signal output
rlabel metal2 s 157890 119200 157946 120000 6 mem_data_o[7]
port 595 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 mem_data_o[8]
port 596 nsew signal output
rlabel metal2 s 160834 119200 160890 120000 6 mem_data_o[9]
port 597 nsew signal output
rlabel metal2 s 148046 119200 148102 120000 6 mem_raddr_o[0]
port 598 nsew signal output
rlabel metal3 s 179200 12112 180000 12232 6 mem_raddr_o[1]
port 599 nsew signal output
rlabel metal3 s 179200 15648 180000 15768 6 mem_raddr_o[2]
port 600 nsew signal output
rlabel metal3 s 179200 22720 180000 22840 6 mem_raddr_o[3]
port 601 nsew signal output
rlabel metal2 s 154854 119200 154910 120000 6 mem_raddr_o[4]
port 602 nsew signal output
rlabel metal3 s 0 112480 800 112600 6 mem_raddr_o[5]
port 603 nsew signal output
rlabel metal3 s 179200 43936 180000 44056 6 mem_raddr_o[6]
port 604 nsew signal output
rlabel metal3 s 179200 54544 180000 54664 6 mem_raddr_o[7]
port 605 nsew signal output
rlabel metal2 s 162950 0 163006 800 6 mem_raddr_o[8]
port 606 nsew signal output
rlabel metal2 s 165618 0 165674 800 6 mem_raddr_o[9]
port 607 nsew signal output
rlabel metal3 s 179200 1640 180000 1760 6 mem_renb_o
port 608 nsew signal output
rlabel metal3 s 179200 5040 180000 5160 6 mem_waddr_o[0]
port 609 nsew signal output
rlabel metal3 s 0 111120 800 111240 6 mem_waddr_o[1]
port 610 nsew signal output
rlabel metal3 s 179200 19184 180000 19304 6 mem_waddr_o[2]
port 611 nsew signal output
rlabel metal3 s 179200 26256 180000 26376 6 mem_waddr_o[3]
port 612 nsew signal output
rlabel metal3 s 179200 33328 180000 33448 6 mem_waddr_o[4]
port 613 nsew signal output
rlabel metal2 s 156878 119200 156934 120000 6 mem_waddr_o[5]
port 614 nsew signal output
rlabel metal3 s 179200 47472 180000 47592 6 mem_waddr_o[6]
port 615 nsew signal output
rlabel metal2 s 158810 119200 158866 120000 6 mem_waddr_o[7]
port 616 nsew signal output
rlabel metal2 s 159822 119200 159878 120000 6 mem_waddr_o[8]
port 617 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 mem_waddr_o[9]
port 618 nsew signal output
rlabel metal2 s 145194 0 145250 800 6 mem_wenb_o
port 619 nsew signal output
rlabel metal2 s 112626 119200 112682 120000 6 phase0_in[0]
port 620 nsew signal input
rlabel metal2 s 142066 119200 142122 120000 6 phase0_in[10]
port 621 nsew signal input
rlabel metal2 s 115570 119200 115626 120000 6 phase0_in[1]
port 622 nsew signal input
rlabel metal2 s 118514 119200 118570 120000 6 phase0_in[2]
port 623 nsew signal input
rlabel metal2 s 121458 119200 121514 120000 6 phase0_in[3]
port 624 nsew signal input
rlabel metal2 s 124402 119200 124458 120000 6 phase0_in[4]
port 625 nsew signal input
rlabel metal2 s 127346 119200 127402 120000 6 phase0_in[5]
port 626 nsew signal input
rlabel metal2 s 130290 119200 130346 120000 6 phase0_in[6]
port 627 nsew signal input
rlabel metal2 s 133234 119200 133290 120000 6 phase0_in[7]
port 628 nsew signal input
rlabel metal2 s 136178 119200 136234 120000 6 phase0_in[8]
port 629 nsew signal input
rlabel metal2 s 139122 119200 139178 120000 6 phase0_in[9]
port 630 nsew signal input
rlabel metal2 s 113546 119200 113602 120000 6 phase1_in[0]
port 631 nsew signal input
rlabel metal2 s 143078 119200 143134 120000 6 phase1_in[10]
port 632 nsew signal input
rlabel metal2 s 116490 119200 116546 120000 6 phase1_in[1]
port 633 nsew signal input
rlabel metal2 s 119434 119200 119490 120000 6 phase1_in[2]
port 634 nsew signal input
rlabel metal2 s 122470 119200 122526 120000 6 phase1_in[3]
port 635 nsew signal input
rlabel metal2 s 125414 119200 125470 120000 6 phase1_in[4]
port 636 nsew signal input
rlabel metal2 s 128358 119200 128414 120000 6 phase1_in[5]
port 637 nsew signal input
rlabel metal2 s 131302 119200 131358 120000 6 phase1_in[6]
port 638 nsew signal input
rlabel metal2 s 134246 119200 134302 120000 6 phase1_in[7]
port 639 nsew signal input
rlabel metal2 s 137190 119200 137246 120000 6 phase1_in[8]
port 640 nsew signal input
rlabel metal2 s 140134 119200 140190 120000 6 phase1_in[9]
port 641 nsew signal input
rlabel metal2 s 114558 119200 114614 120000 6 phase2_in[0]
port 642 nsew signal input
rlabel metal2 s 144090 119200 144146 120000 6 phase2_in[10]
port 643 nsew signal input
rlabel metal2 s 117502 119200 117558 120000 6 phase2_in[1]
port 644 nsew signal input
rlabel metal2 s 120446 119200 120502 120000 6 phase2_in[2]
port 645 nsew signal input
rlabel metal2 s 123390 119200 123446 120000 6 phase2_in[3]
port 646 nsew signal input
rlabel metal2 s 126334 119200 126390 120000 6 phase2_in[4]
port 647 nsew signal input
rlabel metal2 s 129278 119200 129334 120000 6 phase2_in[5]
port 648 nsew signal input
rlabel metal2 s 132222 119200 132278 120000 6 phase2_in[6]
port 649 nsew signal input
rlabel metal2 s 135258 119200 135314 120000 6 phase2_in[7]
port 650 nsew signal input
rlabel metal2 s 138202 119200 138258 120000 6 phase2_in[8]
port 651 nsew signal input
rlabel metal2 s 141146 119200 141202 120000 6 phase2_in[9]
port 652 nsew signal input
rlabel metal2 s 147954 0 148010 800 6 vco_enb_o[0]
port 653 nsew signal output
rlabel metal3 s 0 111392 800 111512 6 vco_enb_o[1]
port 654 nsew signal output
rlabel metal2 s 153382 0 153438 800 6 vco_enb_o[2]
port 655 nsew signal output
rlabel metal2 s 662 0 718 800 6 wb_clk_i
port 656 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wb_rst_i
port 657 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_ack_o
port 658 nsew signal output
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[0]
port 659 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 wbs_adr_i[10]
port 660 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 wbs_adr_i[11]
port 661 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 wbs_adr_i[12]
port 662 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_adr_i[13]
port 663 nsew signal input
rlabel metal2 s 71502 0 71558 800 6 wbs_adr_i[14]
port 664 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 wbs_adr_i[15]
port 665 nsew signal input
rlabel metal2 s 79690 0 79746 800 6 wbs_adr_i[16]
port 666 nsew signal input
rlabel metal2 s 83830 0 83886 800 6 wbs_adr_i[17]
port 667 nsew signal input
rlabel metal2 s 87878 0 87934 800 6 wbs_adr_i[18]
port 668 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 wbs_adr_i[19]
port 669 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 wbs_adr_i[1]
port 670 nsew signal input
rlabel metal2 s 96066 0 96122 800 6 wbs_adr_i[20]
port 671 nsew signal input
rlabel metal2 s 100206 0 100262 800 6 wbs_adr_i[21]
port 672 nsew signal input
rlabel metal2 s 104254 0 104310 800 6 wbs_adr_i[22]
port 673 nsew signal input
rlabel metal2 s 108394 0 108450 800 6 wbs_adr_i[23]
port 674 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 wbs_adr_i[24]
port 675 nsew signal input
rlabel metal2 s 116582 0 116638 800 6 wbs_adr_i[25]
port 676 nsew signal input
rlabel metal2 s 120630 0 120686 800 6 wbs_adr_i[26]
port 677 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 wbs_adr_i[27]
port 678 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 wbs_adr_i[28]
port 679 nsew signal input
rlabel metal2 s 132958 0 133014 800 6 wbs_adr_i[29]
port 680 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 wbs_adr_i[2]
port 681 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 wbs_adr_i[30]
port 682 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 wbs_adr_i[31]
port 683 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[3]
port 684 nsew signal input
rlabel metal2 s 30654 0 30710 800 6 wbs_adr_i[4]
port 685 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 wbs_adr_i[5]
port 686 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 wbs_adr_i[6]
port 687 nsew signal input
rlabel metal2 s 42890 0 42946 800 6 wbs_adr_i[7]
port 688 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 wbs_adr_i[8]
port 689 nsew signal input
rlabel metal2 s 51078 0 51134 800 6 wbs_adr_i[9]
port 690 nsew signal input
rlabel metal2 s 4710 0 4766 800 6 wbs_cyc_i
port 691 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[0]
port 692 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 wbs_dat_i[10]
port 693 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_dat_i[11]
port 694 nsew signal input
rlabel metal2 s 64694 0 64750 800 6 wbs_dat_i[12]
port 695 nsew signal input
rlabel metal2 s 68834 0 68890 800 6 wbs_dat_i[13]
port 696 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_i[14]
port 697 nsew signal input
rlabel metal2 s 77022 0 77078 800 6 wbs_dat_i[15]
port 698 nsew signal input
rlabel metal2 s 81070 0 81126 800 6 wbs_dat_i[16]
port 699 nsew signal input
rlabel metal2 s 85210 0 85266 800 6 wbs_dat_i[17]
port 700 nsew signal input
rlabel metal2 s 89258 0 89314 800 6 wbs_dat_i[18]
port 701 nsew signal input
rlabel metal2 s 93398 0 93454 800 6 wbs_dat_i[19]
port 702 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_dat_i[1]
port 703 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_dat_i[20]
port 704 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 wbs_dat_i[21]
port 705 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 wbs_dat_i[22]
port 706 nsew signal input
rlabel metal2 s 109774 0 109830 800 6 wbs_dat_i[23]
port 707 nsew signal input
rlabel metal2 s 113822 0 113878 800 6 wbs_dat_i[24]
port 708 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 wbs_dat_i[25]
port 709 nsew signal input
rlabel metal2 s 122010 0 122066 800 6 wbs_dat_i[26]
port 710 nsew signal input
rlabel metal2 s 126058 0 126114 800 6 wbs_dat_i[27]
port 711 nsew signal input
rlabel metal2 s 130198 0 130254 800 6 wbs_dat_i[28]
port 712 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 wbs_dat_i[29]
port 713 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_dat_i[2]
port 714 nsew signal input
rlabel metal2 s 138386 0 138442 800 6 wbs_dat_i[30]
port 715 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 wbs_dat_i[31]
port 716 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 wbs_dat_i[3]
port 717 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 wbs_dat_i[4]
port 718 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_dat_i[5]
port 719 nsew signal input
rlabel metal2 s 40130 0 40186 800 6 wbs_dat_i[6]
port 720 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 wbs_dat_i[7]
port 721 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_dat_i[8]
port 722 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_dat_i[9]
port 723 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_dat_o[0]
port 724 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 wbs_dat_o[10]
port 725 nsew signal output
rlabel metal2 s 62026 0 62082 800 6 wbs_dat_o[11]
port 726 nsew signal output
rlabel metal2 s 66074 0 66130 800 6 wbs_dat_o[12]
port 727 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 wbs_dat_o[13]
port 728 nsew signal output
rlabel metal2 s 74262 0 74318 800 6 wbs_dat_o[14]
port 729 nsew signal output
rlabel metal2 s 78402 0 78458 800 6 wbs_dat_o[15]
port 730 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 wbs_dat_o[16]
port 731 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 wbs_dat_o[17]
port 732 nsew signal output
rlabel metal2 s 90638 0 90694 800 6 wbs_dat_o[18]
port 733 nsew signal output
rlabel metal2 s 94686 0 94742 800 6 wbs_dat_o[19]
port 734 nsew signal output
rlabel metal2 s 16946 0 17002 800 6 wbs_dat_o[1]
port 735 nsew signal output
rlabel metal2 s 98826 0 98882 800 6 wbs_dat_o[20]
port 736 nsew signal output
rlabel metal2 s 102874 0 102930 800 6 wbs_dat_o[21]
port 737 nsew signal output
rlabel metal2 s 107014 0 107070 800 6 wbs_dat_o[22]
port 738 nsew signal output
rlabel metal2 s 111062 0 111118 800 6 wbs_dat_o[23]
port 739 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 wbs_dat_o[24]
port 740 nsew signal output
rlabel metal2 s 119250 0 119306 800 6 wbs_dat_o[25]
port 741 nsew signal output
rlabel metal2 s 123390 0 123446 800 6 wbs_dat_o[26]
port 742 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 wbs_dat_o[27]
port 743 nsew signal output
rlabel metal2 s 131578 0 131634 800 6 wbs_dat_o[28]
port 744 nsew signal output
rlabel metal2 s 135626 0 135682 800 6 wbs_dat_o[29]
port 745 nsew signal output
rlabel metal2 s 22466 0 22522 800 6 wbs_dat_o[2]
port 746 nsew signal output
rlabel metal2 s 139766 0 139822 800 6 wbs_dat_o[30]
port 747 nsew signal output
rlabel metal2 s 143814 0 143870 800 6 wbs_dat_o[31]
port 748 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[3]
port 749 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_o[4]
port 750 nsew signal output
rlabel metal2 s 37462 0 37518 800 6 wbs_dat_o[5]
port 751 nsew signal output
rlabel metal2 s 41510 0 41566 800 6 wbs_dat_o[6]
port 752 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 wbs_dat_o[7]
port 753 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 wbs_dat_o[8]
port 754 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 wbs_dat_o[9]
port 755 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 wbs_sel_i[0]
port 756 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_sel_i[1]
port 757 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 wbs_sel_i[2]
port 758 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 wbs_sel_i[3]
port 759 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 wbs_stb_i
port 760 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_we_i
port 761 nsew signal input
rlabel metal2 s 149334 0 149390 800 6 wmask_o[0]
port 762 nsew signal output
rlabel metal2 s 152002 0 152058 800 6 wmask_o[1]
port 763 nsew signal output
rlabel metal2 s 152922 119200 152978 120000 6 wmask_o[2]
port 764 nsew signal output
rlabel metal2 s 157430 0 157486 800 6 wmask_o[3]
port 765 nsew signal output
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 766 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 767 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 768 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 769 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 770 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 771 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 772 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 773 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 775 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 776 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 777 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 778 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 779 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 780 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 781 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 782 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 783 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 784 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 785 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 786 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 787 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 788 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 789 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 790 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 791 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 792 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 793 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 794 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 795 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 796 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 797 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 798 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 799 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 800 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 801 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 802 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 803 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 804 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 805 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 806 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 807 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 808 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 809 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 810 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 811 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 812 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 813 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 14779026
string GDS_START 980350
<< end >>

