magic
tech sky130A
magscale 1 2
timestamp 1637924323
<< obsli1 >>
rect 1104 2159 52808 51697
<< obsm1 >>
rect 750 2048 53162 51728
<< metal2 >>
rect 2410 53200 2466 54000
rect 7286 53200 7342 54000
rect 12162 53200 12218 54000
rect 17130 53200 17186 54000
rect 22006 53200 22062 54000
rect 26882 53200 26938 54000
rect 31850 53200 31906 54000
rect 36726 53200 36782 54000
rect 41602 53200 41658 54000
rect 46570 53200 46626 54000
rect 51446 53200 51502 54000
rect 754 0 810 800
rect 2318 0 2374 800
rect 3974 0 4030 800
rect 5630 0 5686 800
rect 7286 0 7342 800
rect 8850 0 8906 800
rect 10506 0 10562 800
rect 12162 0 12218 800
rect 13818 0 13874 800
rect 15474 0 15530 800
rect 17038 0 17094 800
rect 18694 0 18750 800
rect 20350 0 20406 800
rect 22006 0 22062 800
rect 23662 0 23718 800
rect 25226 0 25282 800
rect 26882 0 26938 800
rect 28538 0 28594 800
rect 30194 0 30250 800
rect 31758 0 31814 800
rect 33414 0 33470 800
rect 35070 0 35126 800
rect 36726 0 36782 800
rect 38382 0 38438 800
rect 39946 0 40002 800
rect 41602 0 41658 800
rect 43258 0 43314 800
rect 44914 0 44970 800
rect 46570 0 46626 800
rect 48134 0 48190 800
rect 49790 0 49846 800
rect 51446 0 51502 800
rect 53102 0 53158 800
<< obsm2 >>
rect 756 53144 2354 53258
rect 2522 53144 7230 53258
rect 7398 53144 12106 53258
rect 12274 53144 17074 53258
rect 17242 53144 21950 53258
rect 22118 53144 26826 53258
rect 26994 53144 31794 53258
rect 31962 53144 36670 53258
rect 36838 53144 41546 53258
rect 41714 53144 46514 53258
rect 46682 53144 51390 53258
rect 51558 53144 53156 53258
rect 756 856 53156 53144
rect 866 800 2262 856
rect 2430 800 3918 856
rect 4086 800 5574 856
rect 5742 800 7230 856
rect 7398 800 8794 856
rect 8962 800 10450 856
rect 10618 800 12106 856
rect 12274 800 13762 856
rect 13930 800 15418 856
rect 15586 800 16982 856
rect 17150 800 18638 856
rect 18806 800 20294 856
rect 20462 800 21950 856
rect 22118 800 23606 856
rect 23774 800 25170 856
rect 25338 800 26826 856
rect 26994 800 28482 856
rect 28650 800 30138 856
rect 30306 800 31702 856
rect 31870 800 33358 856
rect 33526 800 35014 856
rect 35182 800 36670 856
rect 36838 800 38326 856
rect 38494 800 39890 856
rect 40058 800 41546 856
rect 41714 800 43202 856
rect 43370 800 44858 856
rect 45026 800 46514 856
rect 46682 800 48078 856
rect 48246 800 49734 856
rect 49902 800 51390 856
rect 51558 800 53046 856
<< metal3 >>
rect 0 51824 800 51944
rect 0 47608 800 47728
rect 0 43528 800 43648
rect 0 39312 800 39432
rect 0 35232 800 35352
rect 0 31016 800 31136
rect 0 26936 800 27056
rect 0 22720 800 22840
rect 0 18640 800 18760
rect 0 14424 800 14544
rect 0 10344 800 10464
rect 0 6128 800 6248
rect 0 2048 800 2168
<< obsm3 >>
rect 880 51744 50608 51917
rect 800 47808 50608 51744
rect 880 47528 50608 47808
rect 800 43728 50608 47528
rect 880 43448 50608 43728
rect 800 39512 50608 43448
rect 880 39232 50608 39512
rect 800 35432 50608 39232
rect 880 35152 50608 35432
rect 800 31216 50608 35152
rect 880 30936 50608 31216
rect 800 27136 50608 30936
rect 880 26856 50608 27136
rect 800 22920 50608 26856
rect 880 22640 50608 22920
rect 800 18840 50608 22640
rect 880 18560 50608 18840
rect 800 14624 50608 18560
rect 880 14344 50608 14624
rect 800 10544 50608 14344
rect 880 10264 50608 10544
rect 800 6328 50608 10264
rect 880 6048 50608 6328
rect 800 2248 50608 6048
rect 880 2075 50608 2248
<< metal4 >>
rect 4208 2128 4528 51728
rect 19568 2128 19888 51728
rect 34928 2128 35248 51728
rect 50288 2128 50608 51728
<< obsm4 >>
rect 15147 11867 19488 38317
rect 19968 11867 20181 38317
<< labels >>
rlabel metal3 s 0 2048 800 2168 6 clk
port 1 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 data_out[0]
port 2 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 data_out[10]
port 3 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 data_out[11]
port 4 nsew signal output
rlabel metal2 s 22006 0 22062 800 6 data_out[12]
port 5 nsew signal output
rlabel metal2 s 23662 0 23718 800 6 data_out[13]
port 6 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 data_out[14]
port 7 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 data_out[15]
port 8 nsew signal output
rlabel metal2 s 28538 0 28594 800 6 data_out[16]
port 9 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 data_out[17]
port 10 nsew signal output
rlabel metal2 s 31758 0 31814 800 6 data_out[18]
port 11 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 data_out[19]
port 12 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 data_out[1]
port 13 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 data_out[20]
port 14 nsew signal output
rlabel metal2 s 36726 0 36782 800 6 data_out[21]
port 15 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 data_out[22]
port 16 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 data_out[23]
port 17 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 data_out[24]
port 18 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 data_out[25]
port 19 nsew signal output
rlabel metal2 s 44914 0 44970 800 6 data_out[26]
port 20 nsew signal output
rlabel metal2 s 46570 0 46626 800 6 data_out[27]
port 21 nsew signal output
rlabel metal2 s 48134 0 48190 800 6 data_out[28]
port 22 nsew signal output
rlabel metal2 s 49790 0 49846 800 6 data_out[29]
port 23 nsew signal output
rlabel metal2 s 5630 0 5686 800 6 data_out[2]
port 24 nsew signal output
rlabel metal2 s 51446 0 51502 800 6 data_out[30]
port 25 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 data_out[31]
port 26 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 data_out[3]
port 27 nsew signal output
rlabel metal2 s 8850 0 8906 800 6 data_out[4]
port 28 nsew signal output
rlabel metal2 s 10506 0 10562 800 6 data_out[5]
port 29 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 data_out[6]
port 30 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 data_out[7]
port 31 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 data_out[8]
port 32 nsew signal output
rlabel metal2 s 17038 0 17094 800 6 data_out[9]
port 33 nsew signal output
rlabel metal2 s 754 0 810 800 6 data_valid_out
port 34 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 enable_in
port 35 nsew signal input
rlabel metal3 s 0 14424 800 14544 6 oversample_in[0]
port 36 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 oversample_in[1]
port 37 nsew signal input
rlabel metal3 s 0 22720 800 22840 6 oversample_in[2]
port 38 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 oversample_in[3]
port 39 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 oversample_in[4]
port 40 nsew signal input
rlabel metal3 s 0 35232 800 35352 6 oversample_in[5]
port 41 nsew signal input
rlabel metal3 s 0 39312 800 39432 6 oversample_in[6]
port 42 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 oversample_in[7]
port 43 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 oversample_in[8]
port 44 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 oversample_in[9]
port 45 nsew signal input
rlabel metal2 s 2410 53200 2466 54000 6 phase_in[0]
port 46 nsew signal input
rlabel metal2 s 51446 53200 51502 54000 6 phase_in[10]
port 47 nsew signal input
rlabel metal2 s 7286 53200 7342 54000 6 phase_in[1]
port 48 nsew signal input
rlabel metal2 s 12162 53200 12218 54000 6 phase_in[2]
port 49 nsew signal input
rlabel metal2 s 17130 53200 17186 54000 6 phase_in[3]
port 50 nsew signal input
rlabel metal2 s 22006 53200 22062 54000 6 phase_in[4]
port 51 nsew signal input
rlabel metal2 s 26882 53200 26938 54000 6 phase_in[5]
port 52 nsew signal input
rlabel metal2 s 31850 53200 31906 54000 6 phase_in[6]
port 53 nsew signal input
rlabel metal2 s 36726 53200 36782 54000 6 phase_in[7]
port 54 nsew signal input
rlabel metal2 s 41602 53200 41658 54000 6 phase_in[8]
port 55 nsew signal input
rlabel metal2 s 46570 53200 46626 54000 6 phase_in[9]
port 56 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 rst
port 57 nsew signal input
rlabel metal4 s 4208 2128 4528 51728 6 vccd1
port 58 nsew power input
rlabel metal4 s 34928 2128 35248 51728 6 vccd1
port 58 nsew power input
rlabel metal4 s 19568 2128 19888 51728 6 vssd1
port 59 nsew ground input
rlabel metal4 s 50288 2128 50608 51728 6 vssd1
port 59 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 54000 54000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc/runs/vco_adc/results/magic/vco_adc.gds
string GDS_END 7841906
string GDS_START 693900
<< end >>

