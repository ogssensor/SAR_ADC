* NGSPICE file created from vco_adc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_4 abstract view
.subckt sky130_fd_sc_hd__o2111ai_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_1 abstract view
.subckt sky130_fd_sc_hd__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2ai_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_4 abstract view
.subckt sky130_fd_sc_hd__o41ai_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_2 abstract view
.subckt sky130_fd_sc_hd__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt vco_adc clk data_out[0] data_out[10] data_out[11] data_out[12] data_out[13]
+ data_out[14] data_out[15] data_out[16] data_out[17] data_out[18] data_out[19] data_out[1]
+ data_out[20] data_out[21] data_out[22] data_out[23] data_out[24] data_out[25] data_out[26]
+ data_out[27] data_out[28] data_out[29] data_out[2] data_out[30] data_out[31] data_out[3]
+ data_out[4] data_out[5] data_out[6] data_out[7] data_out[8] data_out[9] data_valid_out
+ enable_in oversample_in[0] oversample_in[1] oversample_in[2] oversample_in[3] oversample_in[4]
+ oversample_in[5] oversample_in[6] oversample_in[7] oversample_in[8] oversample_in[9]
+ phase_in[0] phase_in[10] phase_in[1] phase_in[2] phase_in[3] phase_in[4] phase_in[5]
+ phase_in[6] phase_in[7] phase_in[8] phase_in[9] rst vccd1 vssd1
XFILLER_79_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3155_ _5277_/Q vssd1 vssd1 vccd1 vccd1 _3730_/B sky130_fd_sc_hd__inv_2
XFILLER_82_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3086_ _3787_/B _5160_/Q _3351_/A _3359_/B vssd1 vssd1 vccd1 vccd1 _3346_/B sky130_fd_sc_hd__a22oi_4
XFILLER_54_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3988_ _5002_/Q _5002_/D vssd1 vssd1 vccd1 vccd1 _3990_/B sky130_fd_sc_hd__and2_1
XFILLER_22_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2939_ _3613_/A vssd1 vssd1 vccd1 vccd1 _2939_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4609_ _5034_/Q _5066_/Q vssd1 vssd1 vccd1 vccd1 _4671_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_89_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4960_ _4966_/B _4962_/B _4960_/C vssd1 vssd1 vccd1 vccd1 _4960_/X sky130_fd_sc_hd__and3_1
X_3911_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3911_/X sky130_fd_sc_hd__clkbuf_2
X_4891_ _4891_/A _5018_/Q vssd1 vssd1 vccd1 vccd1 _4891_/X sky130_fd_sc_hd__and2_1
X_3842_ _5139_/Q _3835_/X _3830_/X _3841_/Y vssd1 vssd1 vccd1 vccd1 _5139_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3773_ _3781_/A _3773_/B vssd1 vssd1 vccd1 vccd1 _3773_/Y sky130_fd_sc_hd__nand2_1
X_2724_ _2962_/A _2958_/A vssd1 vssd1 vccd1 vccd1 _2724_/Y sky130_fd_sc_hd__nand2_1
X_2655_ _2655_/A vssd1 vssd1 vccd1 vccd1 _2776_/A sky130_fd_sc_hd__inv_2
X_2586_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2586_/X sky130_fd_sc_hd__clkbuf_2
X_4325_ _5063_/Q vssd1 vssd1 vccd1 vccd1 _4661_/B sky130_fd_sc_hd__inv_2
XFILLER_59_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4256_ _4460_/A _4462_/A vssd1 vssd1 vccd1 vccd1 _4367_/A sky130_fd_sc_hd__nor2_1
X_4187_ _4185_/Y _4321_/A _4186_/X vssd1 vssd1 vccd1 vccd1 _5093_/D sky130_fd_sc_hd__a21oi_1
X_3207_ _3180_/Y _3183_/Y _3204_/Y _3206_/X vssd1 vssd1 vccd1 vccd1 _3207_/X sky130_fd_sc_hd__a31o_1
X_3138_ _5172_/Q _3752_/B vssd1 vssd1 vccd1 vccd1 _3138_/Y sky130_fd_sc_hd__nor2_1
X_3069_ _3756_/B _5171_/Q vssd1 vssd1 vccd1 vccd1 _3123_/A sky130_fd_sc_hd__nand2_1
XPHY_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5090_ _5118_/CLK _5090_/D vssd1 vssd1 vccd1 vccd1 _5090_/Q sky130_fd_sc_hd__dfxtp_1
X_4110_ _4110_/A _4110_/B vssd1 vssd1 vccd1 vccd1 _5112_/D sky130_fd_sc_hd__nor2_1
X_4041_ _4041_/A _4045_/C _4041_/C vssd1 vssd1 vccd1 vccd1 _4056_/B sky130_fd_sc_hd__nand3_4
XFILLER_83_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4943_ _5120_/Q _4944_/A vssd1 vssd1 vccd1 vccd1 _4946_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4874_ _4878_/C _4878_/B vssd1 vssd1 vccd1 vccd1 _4874_/Y sky130_fd_sc_hd__nand2_1
X_3825_ _5146_/Q _3822_/X _3817_/X _3824_/Y vssd1 vssd1 vccd1 vccd1 _5146_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3756_ _3765_/A _3756_/B vssd1 vssd1 vccd1 vccd1 _3756_/Y sky130_fd_sc_hd__nand2_1
X_2707_ _2799_/A _2981_/A vssd1 vssd1 vccd1 vccd1 _2707_/Y sky130_fd_sc_hd__nor2_1
X_3687_ _3687_/A _3687_/B vssd1 vssd1 vccd1 vccd1 _3687_/Y sky130_fd_sc_hd__nor2_1
X_2638_ _5287_/Q vssd1 vssd1 vccd1 vccd1 _3017_/B sky130_fd_sc_hd__inv_2
XFILLER_87_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2569_ _5036_/Q vssd1 vssd1 vccd1 vccd1 _4682_/A sky130_fd_sc_hd__inv_2
X_4308_ _4546_/A _4546_/B _4307_/Y vssd1 vssd1 vccd1 vccd1 _4534_/B sky130_fd_sc_hd__a21oi_2
XFILLER_58_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5288_ _5288_/CLK _5288_/D vssd1 vssd1 vccd1 vccd1 _5288_/Q sky130_fd_sc_hd__dfxtp_2
X_4239_ _5113_/Q vssd1 vssd1 vccd1 vccd1 _4405_/B sky130_fd_sc_hd__inv_2
XFILLER_74_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4590_ _4588_/B _4587_/Y _4588_/Y _4587_/B _4906_/A vssd1 vssd1 vccd1 vccd1 _5051_/D
+ sky130_fd_sc_hd__a221oi_2
X_3610_ _3610_/A _3610_/B vssd1 vssd1 vccd1 vccd1 _3611_/B sky130_fd_sc_hd__and2_1
X_3541_ _3541_/A _3541_/B _3563_/B vssd1 vssd1 vccd1 vccd1 _3541_/Y sky130_fd_sc_hd__nand3_1
XFILLER_6_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3472_ _3472_/A _3472_/B vssd1 vssd1 vccd1 vccd1 _3635_/B sky130_fd_sc_hd__or2_1
X_5211_ _5228_/CLK _5211_/D vssd1 vssd1 vccd1 vccd1 _5211_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5142_ _5228_/CLK _5142_/D vssd1 vssd1 vccd1 vccd1 _5142_/Q sky130_fd_sc_hd__dfxtp_1
X_5073_ _5076_/CLK _5073_/D vssd1 vssd1 vccd1 vccd1 _5073_/Q sky130_fd_sc_hd__dfxtp_1
X_4024_ _4055_/B vssd1 vssd1 vccd1 vccd1 _4048_/B sky130_fd_sc_hd__inv_2
XFILLER_56_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4926_ _4921_/Y _4922_/Y _4923_/Y _4924_/Y _4925_/X vssd1 vssd1 vccd1 vccd1 _4927_/B
+ sky130_fd_sc_hd__o2111a_1
X_4857_ _5025_/Q _4217_/X _4197_/B _4856_/X vssd1 vssd1 vccd1 vccd1 _5025_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3808_ _5152_/Q _3796_/X _3804_/X _3807_/Y vssd1 vssd1 vccd1 vccd1 _5152_/D sky130_fd_sc_hd__o211a_1
X_4788_ _4788_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4788_/Y sky130_fd_sc_hd__nand2_1
X_3739_ _3739_/A _3739_/B vssd1 vssd1 vccd1 vccd1 _3739_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2972_ _5263_/Q _2924_/X _2968_/Y _2970_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _5263_/D
+ sky130_fd_sc_hd__o221a_1
X_4711_ _4720_/B _4711_/B vssd1 vssd1 vccd1 vccd1 _4757_/B sky130_fd_sc_hd__nand2_2
X_4642_ _4627_/A _4862_/C _4627_/B vssd1 vssd1 vccd1 vccd1 _4849_/B sky130_fd_sc_hd__o21ba_1
X_4573_ _4567_/X _4570_/Y _4571_/X _4550_/X _4572_/Y vssd1 vssd1 vccd1 vccd1 _5054_/D
+ sky130_fd_sc_hd__o311a_1
X_3524_ _3550_/A vssd1 vssd1 vccd1 vccd1 _3524_/Y sky130_fd_sc_hd__inv_2
X_3455_ _3455_/A _3455_/B vssd1 vssd1 vccd1 vccd1 _3651_/A sky130_fd_sc_hd__nand2_1
X_3386_ _3566_/A _3568_/A _3566_/B vssd1 vssd1 vccd1 vccd1 _3386_/X sky130_fd_sc_hd__o21ba_1
XFILLER_84_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5125_ _5125_/CLK _5125_/D vssd1 vssd1 vccd1 vccd1 _5125_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5056_ _5124_/CLK _5056_/D vssd1 vssd1 vccd1 vccd1 _5056_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4007_ _4984_/D vssd1 vssd1 vccd1 vccd1 _4009_/B sky130_fd_sc_hd__inv_2
XFILLER_84_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4909_ _4910_/A hold36/X vssd1 vssd1 vccd1 vccd1 hold37/A sky130_fd_sc_hd__or2_1
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold41 hold41/A vssd1 vssd1 vccd1 vccd1 hold41/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 oversample_in[8] vssd1 vssd1 vccd1 vccd1 hold30/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_5 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3240_ _3247_/B _3247_/A vssd1 vssd1 vccd1 vccd1 _3243_/A sky130_fd_sc_hd__or2_1
XFILLER_66_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3171_ _3241_/B _3167_/Y _3170_/Y _3164_/C vssd1 vssd1 vccd1 vccd1 _3231_/C sky130_fd_sc_hd__o22a_2
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2955_ _2962_/B _2962_/A vssd1 vssd1 vccd1 vccd1 _2957_/A sky130_fd_sc_hd__nand2_1
X_2886_ _2884_/X _2760_/A _2885_/Y vssd1 vssd1 vccd1 vccd1 _2886_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4625_ _5024_/Q _5056_/Q vssd1 vssd1 vccd1 vccd1 _4627_/A sky130_fd_sc_hd__nor2_2
X_4556_ _4556_/A vssd1 vssd1 vccd1 vccd1 _4561_/A sky130_fd_sc_hd__inv_2
X_3507_ _3820_/B _5147_/Q vssd1 vssd1 vccd1 vccd1 _3508_/B sky130_fd_sc_hd__and2_1
XFILLER_89_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4487_ _4487_/A _4487_/B vssd1 vssd1 vccd1 vccd1 _4488_/B sky130_fd_sc_hd__nor2_1
X_3438_ _3677_/B _3438_/B vssd1 vssd1 vccd1 vccd1 _3681_/B sky130_fd_sc_hd__nand2_2
X_3369_ _5252_/Q vssd1 vssd1 vccd1 vccd1 _3798_/B sky130_fd_sc_hd__inv_2
X_5108_ _5108_/CLK _5108_/D vssd1 vssd1 vccd1 vccd1 _5108_/Q sky130_fd_sc_hd__dfxtp_1
X_5039_ _5311_/CLK _5039_/D vssd1 vssd1 vccd1 vccd1 _5039_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput31 _5206_/Q vssd1 vssd1 vccd1 vccd1 data_out[16] sky130_fd_sc_hd__clkbuf_2
Xoutput42 _5216_/Q vssd1 vssd1 vccd1 vccd1 data_out[26] sky130_fd_sc_hd__clkbuf_2
Xoutput53 _5197_/Q vssd1 vssd1 vccd1 vccd1 data_out[7] sky130_fd_sc_hd__clkbuf_2
XFILLER_76_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2740_ _4818_/A _5300_/Q vssd1 vssd1 vccd1 vccd1 _2741_/B sky130_fd_sc_hd__nand2_1
X_2671_ _5302_/Q _4808_/A vssd1 vssd1 vccd1 vccd1 _2926_/B sky130_fd_sc_hd__or2_2
XFILLER_8_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4410_ _4403_/Y _4416_/A _4406_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4411_/B sky130_fd_sc_hd__o2bb2ai_1
X_4341_ _5069_/Q vssd1 vssd1 vccd1 vccd1 _4691_/B sky130_fd_sc_hd__inv_2
X_4272_ _5098_/Q _5066_/Q vssd1 vssd1 vccd1 vccd1 _4504_/B sky130_fd_sc_hd__and2_1
X_3223_ _3223_/A _3223_/B _3223_/C vssd1 vssd1 vccd1 vccd1 _3224_/A sky130_fd_sc_hd__or3_1
X_3154_ _3154_/A _3154_/B vssd1 vssd1 vccd1 vccd1 _3237_/A sky130_fd_sc_hd__nand2_1
X_3085_ _5159_/Q _5255_/Q vssd1 vssd1 vccd1 vccd1 _3359_/B sky130_fd_sc_hd__or2b_2
XFILLER_35_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3987_ _5002_/Q _5002_/D vssd1 vssd1 vccd1 vccd1 _3990_/A sky130_fd_sc_hd__nor2_2
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2938_ _5269_/Q _2924_/X _2935_/X _2937_/Y _2899_/X vssd1 vssd1 vccd1 vccd1 _5269_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2869_ _3262_/A vssd1 vssd1 vccd1 vccd1 _2869_/X sky130_fd_sc_hd__buf_2
X_4608_ _4608_/A vssd1 vssd1 vccd1 vccd1 _4767_/A sky130_fd_sc_hd__inv_2
X_4539_ _4492_/X _5060_/Q _4537_/Y _4538_/X _4508_/X vssd1 vssd1 vccd1 vccd1 _5060_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_2_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3910_ _3907_/X _4976_/X _3893_/X _3909_/Y vssd1 vssd1 vccd1 vccd1 _5119_/D sky130_fd_sc_hd__o211a_1
X_4890_ _5018_/Q _4891_/A vssd1 vssd1 vccd1 vccd1 _4890_/Y sky130_fd_sc_hd__nor2_1
XFILLER_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3841_ _3847_/A _3841_/B vssd1 vssd1 vccd1 vccd1 _3841_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3772_ _5166_/Q _3768_/X _3762_/X _3771_/Y vssd1 vssd1 vccd1 vccd1 _5166_/D sky130_fd_sc_hd__o211a_1
X_2723_ _2726_/A _2723_/B vssd1 vssd1 vccd1 vccd1 _2958_/A sky130_fd_sc_hd__nor2_2
XFILLER_8_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2654_ _2865_/A _2857_/B vssd1 vssd1 vccd1 vccd1 _2655_/A sky130_fd_sc_hd__nand2_1
X_2585_ _5299_/Q _2567_/X _2582_/X _2584_/Y vssd1 vssd1 vccd1 vccd1 _5299_/D sky130_fd_sc_hd__o211a_1
X_4324_ _4523_/A _4523_/B _4323_/X vssd1 vssd1 vccd1 vccd1 _4513_/B sky130_fd_sc_hd__a21oi_2
XFILLER_86_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4255_ _4255_/A vssd1 vssd1 vccd1 vccd1 _4462_/A sky130_fd_sc_hd__inv_2
X_4186_ _4202_/B _4181_/B _4180_/C _4214_/A vssd1 vssd1 vccd1 vccd1 _4186_/X sky130_fd_sc_hd__a31o_1
X_3206_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3206_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_27_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3137_ _5268_/Q vssd1 vssd1 vccd1 vccd1 _3752_/B sky130_fd_sc_hd__inv_2
X_3068_ _5267_/Q vssd1 vssd1 vccd1 vccd1 _3756_/B sky130_fd_sc_hd__inv_2
XPHY_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_77_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4040_ _4040_/A _4040_/B vssd1 vssd1 vccd1 vccd1 _4041_/C sky130_fd_sc_hd__nor2_2
XFILLER_64_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4942_ _4951_/A _4942_/B vssd1 vssd1 vccd1 vccd1 _4942_/X sky130_fd_sc_hd__and2_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4873_ _4528_/A _4870_/Y _4871_/X _2510_/X _4872_/Y vssd1 vssd1 vccd1 vccd1 _5022_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_20_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3824_ _3833_/A _3824_/B vssd1 vssd1 vccd1 vccd1 _3824_/Y sky130_fd_sc_hd__nand2_1
X_3755_ _3755_/A vssd1 vssd1 vccd1 vccd1 _3765_/A sky130_fd_sc_hd__clkbuf_2
X_2706_ _2709_/A _2966_/B vssd1 vssd1 vccd1 vccd1 _2981_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3686_ _3691_/A _3686_/B vssd1 vssd1 vccd1 vccd1 _3687_/B sky130_fd_sc_hd__or2_1
X_2637_ _3604_/A vssd1 vssd1 vccd1 vccd1 _2995_/A sky130_fd_sc_hd__clkbuf_2
X_2568_ _2605_/A vssd1 vssd1 vccd1 vccd1 _2584_/A sky130_fd_sc_hd__buf_1
XFILLER_87_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4307_ _4545_/A _4549_/B vssd1 vssd1 vccd1 vccd1 _4307_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5287_ _5288_/CLK _5287_/D vssd1 vssd1 vccd1 vccd1 _5287_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4238_ _4238_/A _4238_/B _4238_/C vssd1 vssd1 vccd1 vccd1 _5083_/D sky130_fd_sc_hd__and3_1
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4169_ _4169_/A _4169_/B vssd1 vssd1 vccd1 vccd1 _4169_/Y sky130_fd_sc_hd__nor2_1
XFILLER_70_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3540_ _3544_/A _3540_/B _3540_/C vssd1 vssd1 vccd1 vccd1 _3541_/A sky130_fd_sc_hd__nand3b_1
XFILLER_6_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3471_ _3845_/B _5138_/Q vssd1 vssd1 vccd1 vccd1 _3472_/B sky130_fd_sc_hd__and2_1
X_5210_ _5228_/CLK _5210_/D vssd1 vssd1 vccd1 vccd1 _5210_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5141_ _5285_/CLK _5141_/D vssd1 vssd1 vccd1 vccd1 _5141_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5072_ _5076_/CLK _5072_/D vssd1 vssd1 vccd1 vccd1 _5072_/Q sky130_fd_sc_hd__dfxtp_1
X_4023_ _4023_/A _4023_/B vssd1 vssd1 vccd1 vccd1 _4055_/B sky130_fd_sc_hd__or2_1
XFILLER_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4925_ _5005_/Q _4930_/B _4930_/A _5006_/Q vssd1 vssd1 vccd1 vccd1 _4925_/X sky130_fd_sc_hd__o2bb2a_1
X_4856_ _4852_/A _4855_/Y _4588_/A vssd1 vssd1 vccd1 vccd1 _4856_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3807_ _3807_/A _3807_/B vssd1 vssd1 vccd1 vccd1 _3807_/Y sky130_fd_sc_hd__nand2_1
X_4787_ _4787_/A _4787_/B vssd1 vssd1 vccd1 vccd1 _4787_/Y sky130_fd_sc_hd__xnor2_1
X_3738_ _5178_/Q _3728_/X _3736_/X _3737_/Y vssd1 vssd1 vccd1 vccd1 _5178_/D sky130_fd_sc_hd__o211a_1
X_3669_ _3670_/B _3670_/A vssd1 vssd1 vccd1 vccd1 _3669_/X sky130_fd_sc_hd__or2_1
XFILLER_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2971_ _3262_/A vssd1 vssd1 vccd1 vccd1 _2971_/X sky130_fd_sc_hd__clkbuf_2
X_4710_ _4710_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4711_/B sky130_fd_sc_hd__nand2_1
X_4641_ _3000_/A _5054_/Q _4862_/B _4865_/A _4859_/A vssd1 vssd1 vccd1 vccd1 _4849_/A
+ sky130_fd_sc_hd__o2111ai_4
X_4572_ _4572_/A _4858_/B vssd1 vssd1 vccd1 vccd1 _4572_/Y sky130_fd_sc_hd__nand2_1
X_3523_ _5154_/Q _3802_/B vssd1 vssd1 vccd1 vccd1 _3550_/A sky130_fd_sc_hd__nor2_1
X_3454_ _5230_/Q _5134_/Q vssd1 vssd1 vccd1 vccd1 _3658_/B sky130_fd_sc_hd__xor2_2
X_3385_ _3811_/B _5151_/Q vssd1 vssd1 vccd1 vccd1 _3566_/B sky130_fd_sc_hd__and2_1
X_5124_ _5124_/CLK _5124_/D vssd1 vssd1 vccd1 vccd1 _5124_/Q sky130_fd_sc_hd__dfxtp_1
X_5055_ _5062_/CLK _5055_/D vssd1 vssd1 vccd1 vccd1 _5055_/Q sky130_fd_sc_hd__dfxtp_2
X_4006_ _4029_/A _4029_/B _4004_/Y _4005_/X vssd1 vssd1 vccd1 vccd1 _4022_/A sky130_fd_sc_hd__o22ai_4
XFILLER_72_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4908_ _4910_/A hold31/X vssd1 vssd1 vccd1 vccd1 hold33/A sky130_fd_sc_hd__or2_1
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4839_ _5029_/Q _4217_/X _4807_/X _4838_/X vssd1 vssd1 vccd1 vccd1 _5029_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold20 oversample_in[7] vssd1 vssd1 vccd1 vccd1 input9/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold31 input4/X vssd1 vssd1 vccd1 vccd1 hold31/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 hold42/A vssd1 vssd1 vccd1 vccd1 hold42/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_6 _4197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3170_ _3170_/A vssd1 vssd1 vccd1 vccd1 _3170_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2954_ _2954_/A _2954_/B vssd1 vssd1 vccd1 vccd1 _2962_/B sky130_fd_sc_hd__nand2_1
X_2885_ _2885_/A _2885_/B vssd1 vssd1 vccd1 vccd1 _2885_/Y sky130_fd_sc_hd__nor2_1
X_4624_ _4645_/A _4852_/C _4645_/B vssd1 vssd1 vccd1 vccd1 _4840_/A sky130_fd_sc_hd__o21bai_1
X_4555_ _4530_/X _5057_/Q _4540_/X _4554_/X vssd1 vssd1 vccd1 vccd1 _5057_/D sky130_fd_sc_hd__o211a_1
X_3506_ _5147_/Q _3820_/B vssd1 vssd1 vccd1 vccd1 _3512_/A sky130_fd_sc_hd__nor2_1
XFILLER_89_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4486_ _4420_/X _5070_/Q _4483_/Y _4485_/X _4432_/X vssd1 vssd1 vccd1 vccd1 _5070_/D
+ sky130_fd_sc_hd__o221a_1
X_3437_ _3866_/B _5130_/Q vssd1 vssd1 vccd1 vccd1 _3438_/B sky130_fd_sc_hd__nand2_1
X_3368_ _5222_/Q _3365_/X _3366_/Y _3367_/Y _3363_/X vssd1 vssd1 vccd1 vccd1 _5222_/D
+ sky130_fd_sc_hd__o221a_1
X_5107_ _5109_/CLK _5107_/D vssd1 vssd1 vccd1 vccd1 _5107_/Q sky130_fd_sc_hd__dfxtp_1
X_3299_ _3305_/B _3305_/A vssd1 vssd1 vccd1 vccd1 _3300_/A sky130_fd_sc_hd__or2_1
X_5038_ _5040_/CLK _5038_/D vssd1 vssd1 vccd1 vccd1 _5038_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_82_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput32 _5207_/Q vssd1 vssd1 vccd1 vccd1 data_out[17] sky130_fd_sc_hd__clkbuf_2
Xoutput43 _5217_/Q vssd1 vssd1 vccd1 vccd1 data_out[27] sky130_fd_sc_hd__clkbuf_2
Xoutput54 _5198_/Q vssd1 vssd1 vccd1 vccd1 data_out[8] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2670_ _2747_/A vssd1 vssd1 vccd1 vccd1 _2670_/Y sky130_fd_sc_hd__inv_2
X_4340_ _4502_/A _4502_/B _4339_/X vssd1 vssd1 vccd1 vccd1 _4479_/B sky130_fd_sc_hd__a21oi_4
X_4271_ _4271_/A vssd1 vssd1 vccd1 vccd1 _4506_/B sky130_fd_sc_hd__inv_2
X_3222_ _5249_/Q _3210_/X _3220_/Y _3221_/X _3208_/X vssd1 vssd1 vccd1 vccd1 _5249_/D
+ sky130_fd_sc_hd__o221a_1
X_3153_ _3737_/B _5178_/Q vssd1 vssd1 vccd1 vccd1 _3154_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3084_ _5159_/Q _3789_/B _5254_/Q _3083_/Y vssd1 vssd1 vccd1 vccd1 _3351_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3986_ _4998_/Q _4998_/D vssd1 vssd1 vccd1 vccd1 _4031_/C sky130_fd_sc_hd__xor2_4
X_2937_ _2937_/A _2937_/B vssd1 vssd1 vccd1 vccd1 _2937_/Y sky130_fd_sc_hd__nor2_1
X_4607_ _4600_/Y _4604_/X _4598_/B _4606_/Y vssd1 vssd1 vccd1 vccd1 _4608_/A sky130_fd_sc_hd__a211oi_4
X_2868_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3262_/A sky130_fd_sc_hd__clkbuf_2
X_2799_ _2799_/A _2991_/B vssd1 vssd1 vccd1 vccd1 _2799_/X sky130_fd_sc_hd__or2_1
X_4538_ _4537_/B _4537_/A _4484_/X vssd1 vssd1 vccd1 vccd1 _4538_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4469_ _4470_/B _4470_/A vssd1 vssd1 vccd1 vccd1 _4469_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3840_ _5140_/Q _3835_/X _3830_/X _3839_/Y vssd1 vssd1 vccd1 vccd1 _5140_/D sky130_fd_sc_hd__o211a_1
XFILLER_44_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3771_ _3781_/A _3771_/B vssd1 vssd1 vccd1 vccd1 _3771_/Y sky130_fd_sc_hd__nand2_1
X_2722_ _4835_/A _5297_/Q vssd1 vssd1 vccd1 vccd1 _2723_/B sky130_fd_sc_hd__and2_1
XFILLER_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2653_ _2661_/A _2653_/B vssd1 vssd1 vccd1 vccd1 _2857_/B sky130_fd_sc_hd__nor2_1
X_2584_ _2584_/A _4666_/A vssd1 vssd1 vccd1 vccd1 _2584_/Y sky130_fd_sc_hd__nand2_1
X_4323_ _4525_/B _4525_/A _4531_/B vssd1 vssd1 vccd1 vccd1 _4323_/X sky130_fd_sc_hd__or3_1
X_4254_ _4254_/A _4254_/B vssd1 vssd1 vccd1 vccd1 _4255_/A sky130_fd_sc_hd__nor2_1
X_3205_ _3180_/Y _3183_/Y _3204_/Y vssd1 vssd1 vccd1 vccd1 _3205_/Y sky130_fd_sc_hd__a21oi_1
X_4185_ _4185_/A _5092_/Q vssd1 vssd1 vccd1 vccd1 _4185_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3136_ _3278_/A _3278_/B _3135_/Y vssd1 vssd1 vccd1 vccd1 _3257_/A sky130_fd_sc_hd__o21bai_1
XFILLER_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3067_ _5170_/Q _3758_/B vssd1 vssd1 vccd1 vccd1 _3125_/A sky130_fd_sc_hd__nor2_1
XPHY_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3969_ _3970_/B _4988_/Q vssd1 vssd1 vccd1 vccd1 _4023_/B sky130_fd_sc_hd__and2_1
XFILLER_6_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4941_ _4941_/A _4944_/A vssd1 vssd1 vccd1 vccd1 _4942_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4872_ _4872_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4872_/Y sky130_fd_sc_hd__nand2_1
X_3823_ _3823_/A vssd1 vssd1 vccd1 vccd1 _3833_/A sky130_fd_sc_hd__buf_1
X_3754_ _3754_/A vssd1 vssd1 vccd1 vccd1 _3754_/X sky130_fd_sc_hd__clkbuf_2
X_2705_ _4853_/A _5293_/Q vssd1 vssd1 vccd1 vccd1 _2966_/B sky130_fd_sc_hd__nand2_2
X_3685_ _3685_/A _3685_/B vssd1 vssd1 vccd1 vccd1 _3687_/A sky130_fd_sc_hd__nand2_1
X_2636_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3604_/A sky130_fd_sc_hd__clkbuf_2
X_2567_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4306_ _4306_/A _4306_/B vssd1 vssd1 vccd1 vccd1 _4549_/B sky130_fd_sc_hd__nor2_1
X_5286_ _5288_/CLK _5286_/D vssd1 vssd1 vccd1 vccd1 _5286_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4237_ _4237_/A _4587_/B vssd1 vssd1 vccd1 vccd1 _4238_/C sky130_fd_sc_hd__nand2_1
XFILLER_74_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4168_ _4337_/A _4168_/B _4183_/A vssd1 vssd1 vccd1 vccd1 _4172_/C sky130_fd_sc_hd__nor3_4
X_4099_ _5111_/Q vssd1 vssd1 vccd1 vccd1 _4244_/A sky130_fd_sc_hd__inv_2
X_3119_ _3119_/A vssd1 vssd1 vccd1 vccd1 _3301_/A sky130_fd_sc_hd__inv_2
XFILLER_82_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_80_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3470_ _3470_/A vssd1 vssd1 vccd1 vccd1 _3628_/B sky130_fd_sc_hd__inv_2
XFILLER_69_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5140_ _5285_/CLK _5140_/D vssd1 vssd1 vccd1 vccd1 _5140_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5071_ _5076_/CLK _5071_/D vssd1 vssd1 vccd1 vccd1 _5071_/Q sky130_fd_sc_hd__dfxtp_1
X_4022_ _4022_/A _4022_/B _4022_/C vssd1 vssd1 vccd1 vccd1 _4055_/A sky130_fd_sc_hd__nand3_4
XFILLER_49_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4924_ _5118_/Q _5007_/Q vssd1 vssd1 vccd1 vccd1 _4924_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_64_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4855_ _4855_/A _4855_/B vssd1 vssd1 vccd1 vccd1 _4855_/Y sky130_fd_sc_hd__nand2_1
X_3806_ _5153_/Q _3796_/X _3804_/X _3805_/Y vssd1 vssd1 vccd1 vccd1 _5153_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4786_ _5040_/Q _4770_/X _4783_/Y _4784_/X _4785_/X vssd1 vssd1 vccd1 vccd1 _5040_/D
+ sky130_fd_sc_hd__o221a_1
X_3737_ _3739_/A _3737_/B vssd1 vssd1 vccd1 vccd1 _3737_/Y sky130_fd_sc_hd__nand2_1
X_3668_ _3754_/A vssd1 vssd1 vccd1 vccd1 _3668_/X sky130_fd_sc_hd__buf_2
X_2619_ _2892_/A vssd1 vssd1 vccd1 vccd1 _2619_/X sky130_fd_sc_hd__clkbuf_2
X_3599_ _3599_/A _3599_/B vssd1 vssd1 vccd1 vccd1 _3599_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5269_ _5288_/CLK _5269_/D vssd1 vssd1 vccd1 vccd1 _5269_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_43_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2970_ _2968_/B _2968_/A _2969_/X vssd1 vssd1 vccd1 vccd1 _2970_/X sky130_fd_sc_hd__a21o_1
XFILLER_30_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4640_ _4868_/A _4871_/B _4878_/B vssd1 vssd1 vccd1 vccd1 _4859_/A sky130_fd_sc_hd__nand3_2
X_4571_ _4571_/A _4571_/B _4571_/C vssd1 vssd1 vccd1 vccd1 _4571_/X sky130_fd_sc_hd__and3_1
X_3522_ _5250_/Q vssd1 vssd1 vccd1 vccd1 _3802_/B sky130_fd_sc_hd__inv_2
X_3453_ _3450_/B _3663_/B _3450_/A vssd1 vssd1 vccd1 vccd1 _3652_/B sky130_fd_sc_hd__o21ba_1
XFILLER_69_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5123_ _5124_/CLK _5123_/D vssd1 vssd1 vccd1 vccd1 _5123_/Q sky130_fd_sc_hd__dfxtp_1
X_3384_ _5150_/Q _3813_/B vssd1 vssd1 vccd1 vccd1 _3568_/A sky130_fd_sc_hd__nor2_2
XFILLER_69_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5054_ _5062_/CLK _5054_/D vssd1 vssd1 vccd1 vccd1 _5054_/Q sky130_fd_sc_hd__dfxtp_4
X_4005_ _4003_/A _4003_/B _4030_/A _4011_/A vssd1 vssd1 vccd1 vccd1 _4005_/X sky130_fd_sc_hd__o211a_1
XFILLER_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4907_ _4910_/A hold26/X vssd1 vssd1 vccd1 vccd1 hold28/A sky130_fd_sc_hd__or2_1
X_4838_ _4834_/A _4837_/Y _4542_/X vssd1 vssd1 vccd1 vccd1 _4838_/X sky130_fd_sc_hd__a21o_1
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4769_ _5043_/Q _4530_/X _4540_/X _4768_/X vssd1 vssd1 vccd1 vccd1 _5043_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold21 hold21/A vssd1 vssd1 vccd1 vccd1 hold21/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 phase_in[4] vssd1 vssd1 vccd1 vccd1 hold10/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 oversample_in[2] vssd1 vssd1 vccd1 vccd1 input4/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 hold43/A vssd1 vssd1 vccd1 vccd1 hold43/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_7 _4827_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2953_ _5266_/Q _2939_/X _2892_/X _2952_/Y vssd1 vssd1 vccd1 vccd1 _5266_/D sky130_fd_sc_hd__o211a_1
X_2884_ _2893_/B _2893_/A vssd1 vssd1 vccd1 vccd1 _2884_/X sky130_fd_sc_hd__or2_1
XFILLER_30_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4623_ _4853_/A _4623_/B vssd1 vssd1 vccd1 vccd1 _4645_/B sky130_fd_sc_hd__nor2_1
X_4554_ _4549_/A _4553_/Y _4542_/X vssd1 vssd1 vccd1 vccd1 _4554_/X sky130_fd_sc_hd__a21o_1
X_3505_ _5243_/Q vssd1 vssd1 vccd1 vccd1 _3820_/B sky130_fd_sc_hd__inv_2
X_4485_ _4483_/B _4483_/A _4484_/X vssd1 vssd1 vccd1 vccd1 _4485_/X sky130_fd_sc_hd__a21o_1
X_3436_ _3436_/A vssd1 vssd1 vccd1 vccd1 _3685_/A sky130_fd_sc_hd__inv_2
X_3367_ _3705_/A _3367_/B vssd1 vssd1 vccd1 vccd1 _3367_/Y sky130_fd_sc_hd__nand2_1
X_5106_ _5109_/CLK _5106_/D vssd1 vssd1 vccd1 vccd1 _5106_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5037_ _5040_/CLK _5037_/D vssd1 vssd1 vccd1 vccd1 _5037_/Q sky130_fd_sc_hd__dfxtp_1
X_3298_ _3298_/A _3298_/B vssd1 vssd1 vccd1 vccd1 _3305_/A sky130_fd_sc_hd__nor2_1
XFILLER_72_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput33 _5208_/Q vssd1 vssd1 vccd1 vccd1 data_out[18] sky130_fd_sc_hd__clkbuf_2
Xoutput55 _5199_/Q vssd1 vssd1 vccd1 vccd1 data_out[9] sky130_fd_sc_hd__clkbuf_2
Xoutput44 _5218_/Q vssd1 vssd1 vccd1 vccd1 data_out[28] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4270_ _4337_/A _4610_/B vssd1 vssd1 vccd1 vccd1 _4271_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3221_ _3224_/C _3172_/B _3047_/B _3206_/X vssd1 vssd1 vccd1 vccd1 _3221_/X sky130_fd_sc_hd__a31o_1
X_3152_ _5178_/Q _3737_/B vssd1 vssd1 vccd1 vccd1 _3154_/A sky130_fd_sc_hd__or2_1
XFILLER_39_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3083_ _5158_/Q vssd1 vssd1 vccd1 vccd1 _3083_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3985_ _3985_/A _4039_/B vssd1 vssd1 vccd1 vccd1 _4029_/B sky130_fd_sc_hd__and2_1
XFILLER_22_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2936_ _2936_/A _2936_/B vssd1 vssd1 vccd1 vccd1 _2937_/B sky130_fd_sc_hd__and2_1
X_2867_ _2867_/A _3862_/A _2867_/C vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__and3_1
X_4606_ _4606_/A _4774_/B vssd1 vssd1 vccd1 vccd1 _4606_/Y sky130_fd_sc_hd__nor2_2
X_2798_ _2798_/A vssd1 vssd1 vccd1 vccd1 _2991_/B sky130_fd_sc_hd__inv_2
X_4537_ _4537_/A _4537_/B vssd1 vssd1 vccd1 vccd1 _4537_/Y sky130_fd_sc_hd__nor2_1
X_4468_ _4468_/A _4468_/B vssd1 vssd1 vccd1 vccd1 _4470_/A sky130_fd_sc_hd__nor2_1
X_3419_ _5135_/Q _3853_/B vssd1 vssd1 vccd1 vccd1 _3455_/A sky130_fd_sc_hd__or2_1
XFILLER_58_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4399_ _4428_/A _4427_/A _4429_/A vssd1 vssd1 vccd1 vccd1 _4423_/D sky130_fd_sc_hd__a21oi_4
XFILLER_73_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3770_ _3823_/A vssd1 vssd1 vccd1 vccd1 _3781_/A sky130_fd_sc_hd__clkbuf_2
X_2721_ _5297_/Q _4835_/A vssd1 vssd1 vccd1 vccd1 _2726_/A sky130_fd_sc_hd__nor2_2
XFILLER_8_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2652_ _2652_/A vssd1 vssd1 vccd1 vccd1 _2865_/A sky130_fd_sc_hd__inv_2
X_2583_ _5032_/Q vssd1 vssd1 vccd1 vccd1 _4666_/A sky130_fd_sc_hd__inv_2
X_4322_ _4322_/A _4527_/C vssd1 vssd1 vccd1 vccd1 _4531_/B sky130_fd_sc_hd__nand2_1
X_4253_ _4253_/A _4253_/B vssd1 vssd1 vccd1 vccd1 _4460_/A sky130_fd_sc_hd__nand2_1
X_3204_ _3204_/A _3204_/B vssd1 vssd1 vccd1 vccd1 _3204_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4184_ _4181_/Y _4277_/A _4183_/Y vssd1 vssd1 vccd1 vccd1 _5094_/D sky130_fd_sc_hd__a21oi_1
XFILLER_55_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3135_ _3135_/A vssd1 vssd1 vccd1 vccd1 _3135_/Y sky130_fd_sc_hd__inv_2
XFILLER_82_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3066_ _5266_/Q vssd1 vssd1 vccd1 vccd1 _3758_/B sky130_fd_sc_hd__inv_2
XPHY_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3968_ hold46/A vssd1 vssd1 vccd1 vccd1 _3970_/B sky130_fd_sc_hd__inv_2
XFILLER_10_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2919_ _2919_/A _3011_/A vssd1 vssd1 vccd1 vccd1 _2919_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3899_ _3887_/X _4973_/X _3893_/X _3898_/Y vssd1 vssd1 vccd1 vccd1 _5122_/D sky130_fd_sc_hd__o211a_1
XFILLER_12_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_77_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4940_ _4940_/A _4940_/B vssd1 vssd1 vccd1 vccd1 _4944_/A sky130_fd_sc_hd__nor2_2
X_4871_ _4871_/A _4871_/B _4871_/C vssd1 vssd1 vccd1 vccd1 _4871_/X sky130_fd_sc_hd__and3_1
XFILLER_17_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3822_ _3822_/A vssd1 vssd1 vccd1 vccd1 _3822_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3753_ _5172_/Q _3741_/X _3749_/X _3752_/Y vssd1 vssd1 vccd1 vccd1 _5172_/D sky130_fd_sc_hd__o211a_1
X_2704_ _2704_/A _5026_/Q vssd1 vssd1 vccd1 vccd1 _2709_/A sky130_fd_sc_hd__nand2_1
X_3684_ _3868_/B _5129_/Q vssd1 vssd1 vccd1 vccd1 _3685_/B sky130_fd_sc_hd__nand2_1
X_2635_ _2847_/A vssd1 vssd1 vccd1 vccd1 _3642_/A sky130_fd_sc_hd__clkbuf_2
X_4305_ _4305_/A _4549_/C vssd1 vssd1 vccd1 vccd1 _4545_/A sky130_fd_sc_hd__and2_1
X_2566_ _5304_/Q _2548_/X _2563_/X _2565_/Y vssd1 vssd1 vccd1 vccd1 _5304_/D sky130_fd_sc_hd__o211a_1
X_5285_ _5285_/CLK _5285_/D vssd1 vssd1 vccd1 vccd1 _5285_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4236_ _4587_/B _4237_/A vssd1 vssd1 vccd1 vccd1 _4238_/A sky130_fd_sc_hd__or2_1
X_4167_ _4180_/A _4180_/B _4173_/C vssd1 vssd1 vccd1 vccd1 _4183_/A sky130_fd_sc_hd__nand3_4
XFILLER_74_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3118_ _3118_/A _3118_/B vssd1 vssd1 vccd1 vccd1 _3119_/A sky130_fd_sc_hd__nor2_1
X_4098_ _5112_/Q vssd1 vssd1 vccd1 vccd1 _4402_/A sky130_fd_sc_hd__inv_2
XFILLER_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3049_ _5272_/Q vssd1 vssd1 vccd1 vccd1 _3743_/B sky130_fd_sc_hd__inv_2
XPHY_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5070_ _5098_/CLK _5070_/D vssd1 vssd1 vccd1 vccd1 _5070_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4021_ _4022_/C _4022_/A _4017_/A _4017_/B vssd1 vssd1 vccd1 vccd1 _4056_/C sky130_fd_sc_hd__o2bb2ai_2
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4923_ _5121_/Q _5010_/Q vssd1 vssd1 vccd1 vccd1 _4923_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_33_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4854_ _4567_/X _4851_/Y _4852_/X _2510_/X _4853_/Y vssd1 vssd1 vccd1 vccd1 _5026_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_60_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3805_ _3807_/A _3805_/B vssd1 vssd1 vccd1 vccd1 _3805_/Y sky130_fd_sc_hd__nand2_1
X_4785_ _4785_/A vssd1 vssd1 vccd1 vccd1 _4785_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3736_ _3762_/A vssd1 vssd1 vccd1 vccd1 _3736_/X sky130_fd_sc_hd__buf_1
X_3667_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3754_/A sky130_fd_sc_hd__clkbuf_2
X_2618_ _5290_/Q _2604_/X _2600_/X _2617_/Y vssd1 vssd1 vccd1 vccd1 _5290_/D sky130_fd_sc_hd__o211a_1
X_3598_ _3603_/B _3603_/A _3406_/B vssd1 vssd1 vccd1 vccd1 _3599_/B sky130_fd_sc_hd__o21a_1
X_2549_ _2605_/A vssd1 vssd1 vccd1 vccd1 _2565_/A sky130_fd_sc_hd__buf_1
X_5268_ _5268_/CLK _5268_/D vssd1 vssd1 vccd1 vccd1 _5268_/Q sky130_fd_sc_hd__dfxtp_1
X_4219_ _4580_/A _4219_/B vssd1 vssd1 vccd1 vccd1 _4226_/A sky130_fd_sc_hd__or2_1
X_5199_ _5199_/CLK _5199_/D vssd1 vssd1 vccd1 vccd1 _5199_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4570_ _4571_/B _4571_/C _4571_/A vssd1 vssd1 vccd1 vccd1 _4570_/Y sky130_fd_sc_hd__a21oi_1
X_3521_ _5250_/Q _3549_/B _3551_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3521_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_6_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3452_ _3424_/Y _3673_/A _3442_/Y _3451_/Y vssd1 vssd1 vccd1 vccd1 _3652_/A sky130_fd_sc_hd__o211ai_2
X_3383_ _5151_/Q _3811_/B vssd1 vssd1 vccd1 vccd1 _3566_/A sky130_fd_sc_hd__nor2_1
X_5122_ _5125_/CLK _5122_/D vssd1 vssd1 vccd1 vccd1 _5122_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5053_ _5085_/CLK _5053_/D vssd1 vssd1 vccd1 vccd1 _5053_/Q sky130_fd_sc_hd__dfxtp_2
X_4004_ _4011_/A _4030_/A _4011_/C vssd1 vssd1 vccd1 vccd1 _4004_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4906_ _4906_/A hold13/X vssd1 vssd1 vccd1 vccd1 hold15/A sky130_fd_sc_hd__or2_1
X_4837_ _4837_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4837_/Y sky130_fd_sc_hd__nand2_1
X_4768_ _4762_/A _4767_/X _4542_/X vssd1 vssd1 vccd1 vccd1 _4768_/X sky130_fd_sc_hd__a21o_1
X_3719_ _3726_/A _3719_/B vssd1 vssd1 vccd1 vccd1 _3719_/Y sky130_fd_sc_hd__nand2_1
X_4699_ _4699_/A _4701_/B vssd1 vssd1 vccd1 vccd1 _4700_/A sky130_fd_sc_hd__nor2_2
XFILLER_88_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold22 phase_in[9] vssd1 vssd1 vccd1 vccd1 hold22/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 hold11/A vssd1 vssd1 vccd1 vccd1 hold11/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_29_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold44 hold44/A vssd1 vssd1 vccd1 vccd1 hold44/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 hold33/A vssd1 vssd1 vccd1 vccd1 hold33/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_8 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2952_ _2949_/Y _2950_/Y _2951_/X vssd1 vssd1 vccd1 vccd1 _2952_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2883_ _2762_/Y _2882_/Y _2764_/B vssd1 vssd1 vccd1 vccd1 _2893_/A sky130_fd_sc_hd__o21ai_1
X_4622_ _5025_/Q _5057_/Q vssd1 vssd1 vccd1 vccd1 _4852_/C sky130_fd_sc_hd__nand2_1
X_4553_ _4553_/A _4553_/B vssd1 vssd1 vccd1 vccd1 _4553_/Y sky130_fd_sc_hd__nand2_1
X_3504_ _3586_/B _3504_/B vssd1 vssd1 vccd1 vccd1 _3509_/B sky130_fd_sc_hd__or2_1
X_4484_ _4764_/A vssd1 vssd1 vccd1 vccd1 _4484_/X sky130_fd_sc_hd__buf_2
X_3435_ _5129_/Q _3868_/B vssd1 vssd1 vccd1 vccd1 _3436_/A sky130_fd_sc_hd__nor2_1
X_3366_ _5158_/Q _3792_/B vssd1 vssd1 vccd1 vccd1 _3366_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3297_ _5234_/Q _3253_/X _3246_/X _3296_/X vssd1 vssd1 vccd1 vccd1 _5234_/D sky130_fd_sc_hd__o211a_1
X_5105_ _5109_/CLK _5105_/D vssd1 vssd1 vccd1 vccd1 _5105_/Q sky130_fd_sc_hd__dfxtp_1
X_5036_ _5040_/CLK _5036_/D vssd1 vssd1 vccd1 vccd1 _5036_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput34 _5209_/Q vssd1 vssd1 vccd1 vccd1 data_out[19] sky130_fd_sc_hd__clkbuf_2
Xoutput56 _4967_/X vssd1 vssd1 vccd1 vccd1 data_valid_out sky130_fd_sc_hd__clkbuf_2
Xoutput45 _5219_/Q vssd1 vssd1 vccd1 vccd1 data_out[29] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3220_ _3224_/C _3047_/B _3172_/B vssd1 vssd1 vccd1 vccd1 _3220_/Y sky130_fd_sc_hd__a21oi_1
X_3151_ _3151_/A vssd1 vssd1 vccd1 vccd1 _3164_/A sky130_fd_sc_hd__inv_2
XFILLER_39_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3082_ _5160_/Q _3787_/B vssd1 vssd1 vccd1 vccd1 _3346_/A sky130_fd_sc_hd__nor2_4
XFILLER_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3984_ _4039_/B _3985_/A vssd1 vssd1 vccd1 vccd1 _4029_/A sky130_fd_sc_hd__nor2_4
XFILLER_50_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2935_ _2936_/A _2937_/A _2936_/B _2901_/A vssd1 vssd1 vccd1 vccd1 _2935_/X sky130_fd_sc_hd__a31o_1
XFILLER_50_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2866_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3862_/A sky130_fd_sc_hd__buf_2
XFILLER_30_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4605_ _4605_/A vssd1 vssd1 vccd1 vccd1 _4774_/B sky130_fd_sc_hd__inv_2
X_2797_ _2943_/B vssd1 vssd1 vccd1 vccd1 _2797_/Y sky130_fd_sc_hd__inv_2
X_4536_ _4536_/A _4536_/B vssd1 vssd1 vccd1 vccd1 _4537_/B sky130_fd_sc_hd__nand2_1
XFILLER_89_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4467_ _4913_/A _4467_/B vssd1 vssd1 vccd1 vccd1 _5073_/D sky130_fd_sc_hd__nor2_1
X_3418_ _3855_/B _5134_/Q _3455_/B vssd1 vssd1 vccd1 vccd1 _3420_/A sky130_fd_sc_hd__or3b_2
X_4398_ _5111_/Q _5079_/Q vssd1 vssd1 vccd1 vccd1 _4429_/A sky130_fd_sc_hd__nor2_2
X_3349_ _5225_/Q _3321_/X _3347_/Y _3348_/X _3316_/X vssd1 vssd1 vccd1 vccd1 _5225_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5019_ _5027_/CLK _5019_/D vssd1 vssd1 vccd1 vccd1 _5019_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_45_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2720_ _2720_/A vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__inv_2
X_2651_ _2857_/C _2651_/B vssd1 vssd1 vccd1 vccd1 _2652_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2582_ _2892_/A vssd1 vssd1 vccd1 vccd1 _2582_/X sky130_fd_sc_hd__clkbuf_2
X_4321_ _4321_/A _4657_/B vssd1 vssd1 vccd1 vccd1 _4322_/A sky130_fd_sc_hd__nand2_1
X_4252_ _4252_/A _4594_/B vssd1 vssd1 vccd1 vccd1 _4253_/B sky130_fd_sc_hd__nand2_1
X_3203_ _3199_/Y _3200_/Y _3202_/X vssd1 vssd1 vccd1 vccd1 _5252_/D sky130_fd_sc_hd__a21oi_1
XFILLER_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4183_ _4183_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4183_/Y sky130_fd_sc_hd__nand2_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3134_ _3284_/B _3281_/A vssd1 vssd1 vccd1 vccd1 _3135_/A sky130_fd_sc_hd__and2b_1
XFILLER_55_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3065_ _3057_/Y _3063_/X _3055_/A _3064_/Y vssd1 vssd1 vccd1 vccd1 _3236_/A sky130_fd_sc_hd__a211o_1
XPHY_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3967_ _3967_/A _5114_/Q vssd1 vssd1 vccd1 vccd1 _4090_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2918_ _2634_/X _2913_/Y _2914_/X _2915_/X _2917_/Y vssd1 vssd1 vccd1 vccd1 _5273_/D
+ sky130_fd_sc_hd__o311a_1
X_3898_ _4572_/A _3898_/B vssd1 vssd1 vccd1 vccd1 _3898_/Y sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_30_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5250_/CLK sky130_fd_sc_hd__clkbuf_16
X_2849_ _2846_/B _2846_/A _2848_/X vssd1 vssd1 vccd1 vccd1 _2849_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4519_ _4520_/B _4520_/A vssd1 vssd1 vccd1 vccd1 _4519_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 _4987_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_68_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4870_ _4871_/B _4871_/C _4871_/A vssd1 vssd1 vccd1 vccd1 _4870_/Y sky130_fd_sc_hd__a21oi_1
X_3821_ _5147_/Q _3809_/X _3817_/X _3820_/Y vssd1 vssd1 vccd1 vccd1 _5147_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_12_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5001_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3752_ _3752_/A _3752_/B vssd1 vssd1 vccd1 vccd1 _3752_/Y sky130_fd_sc_hd__nand2_1
X_2703_ _5293_/Q vssd1 vssd1 vccd1 vccd1 _2704_/A sky130_fd_sc_hd__inv_2
X_3683_ _5194_/Q _3668_/X _3646_/X _3682_/Y vssd1 vssd1 vccd1 vccd1 _5194_/D sky130_fd_sc_hd__o211a_1
X_2634_ _3615_/A vssd1 vssd1 vccd1 vccd1 _2634_/X sky130_fd_sc_hd__clkbuf_2
X_2565_ _2565_/A _4691_/A vssd1 vssd1 vccd1 vccd1 _2565_/Y sky130_fd_sc_hd__nand2_1
X_4304_ _4304_/A _4643_/B vssd1 vssd1 vccd1 vccd1 _4305_/A sky130_fd_sc_hd__nand2_1
X_5284_ _5285_/CLK _5284_/D vssd1 vssd1 vccd1 vccd1 _5284_/Q sky130_fd_sc_hd__dfxtp_1
X_4235_ _4542_/A _4235_/B vssd1 vssd1 vccd1 vccd1 _4237_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4166_ _4166_/A vssd1 vssd1 vccd1 vccd1 _4173_/C sky130_fd_sc_hd__inv_2
XFILLER_28_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3117_ _3760_/B _5169_/Q vssd1 vssd1 vccd1 vccd1 _3118_/B sky130_fd_sc_hd__and2_1
X_4097_ _4116_/A _4097_/B _4097_/C vssd1 vssd1 vccd1 vccd1 _5114_/D sky130_fd_sc_hd__nor3_1
XFILLER_70_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3048_ _3223_/B _3172_/B _3223_/A _3042_/A _3047_/Y vssd1 vssd1 vccd1 vccd1 _3048_/X
+ sky130_fd_sc_hd__a311o_2
XPHY_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4999_ _5001_/CLK hold1/X vssd1 vssd1 vccd1 vccd1 _5000_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_11_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4020_ _4996_/Q _4996_/D vssd1 vssd1 vccd1 vccd1 _4064_/A sky130_fd_sc_hd__xnor2_4
Xclkbuf_leaf_1_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5109_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_77_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4922_ _4962_/A _4922_/B vssd1 vssd1 vccd1 vccd1 _4922_/Y sky130_fd_sc_hd__nor2_1
XFILLER_33_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4853_ _4853_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4853_/Y sky130_fd_sc_hd__nand2_1
X_3804_ _3830_/A vssd1 vssd1 vccd1 vccd1 _3804_/X sky130_fd_sc_hd__clkbuf_2
X_4784_ _4783_/B _4783_/A _4764_/X vssd1 vssd1 vccd1 vccd1 _4784_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3735_ _5179_/Q _3728_/X _3723_/X _3734_/Y vssd1 vssd1 vccd1 vccd1 _5179_/D sky130_fd_sc_hd__o211a_1
X_3666_ _5197_/Q _3650_/X _3664_/Y _3665_/X _3644_/X vssd1 vssd1 vccd1 vccd1 _5197_/D
+ sky130_fd_sc_hd__o221a_1
X_2617_ _2622_/A _4628_/A vssd1 vssd1 vccd1 vccd1 _2617_/Y sky130_fd_sc_hd__nand2_1
X_3597_ _3608_/B _3405_/Y _3489_/C _3614_/A vssd1 vssd1 vccd1 vccd1 _3603_/A sky130_fd_sc_hd__o22a_1
X_2548_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2548_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5267_ _5267_/CLK _5267_/D vssd1 vssd1 vccd1 vccd1 _5267_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4218_ _4057_/Y _4052_/A _4060_/Y vssd1 vssd1 vccd1 vccd1 _4219_/B sky130_fd_sc_hd__o21a_1
X_5198_ _5199_/CLK _5198_/D vssd1 vssd1 vccd1 vccd1 _5198_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4149_ _4149_/A _4149_/B vssd1 vssd1 vccd1 vccd1 _4154_/A sky130_fd_sc_hd__nand2_1
XFILLER_55_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3520_ _3572_/A _3572_/C _3519_/X vssd1 vssd1 vccd1 vccd1 _3551_/B sky130_fd_sc_hd__a21oi_4
XFILLER_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3451_ _3670_/B _3664_/A vssd1 vssd1 vccd1 vccd1 _3451_/Y sky130_fd_sc_hd__nor2_1
X_3382_ _5247_/Q vssd1 vssd1 vccd1 vccd1 _3811_/B sky130_fd_sc_hd__inv_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5121_ _5124_/CLK _5121_/D vssd1 vssd1 vccd1 vccd1 _5121_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5052_ _5085_/CLK _5052_/D vssd1 vssd1 vccd1 vccd1 _5052_/Q sky130_fd_sc_hd__dfxtp_1
X_4003_ _4003_/A _4003_/B vssd1 vssd1 vccd1 vccd1 _4011_/C sky130_fd_sc_hd__or2_2
XFILLER_84_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4905_ _4906_/A hold16/X vssd1 vssd1 vccd1 vccd1 hold18/A sky130_fd_sc_hd__or2_1
XFILLER_21_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4836_ _4567_/X _4833_/Y _4834_/X _4550_/X _4835_/Y vssd1 vssd1 vccd1 vccd1 _5030_/D
+ sky130_fd_sc_hd__o311a_1
X_4767_ _4767_/A _4767_/B _4761_/A vssd1 vssd1 vccd1 vccd1 _4767_/X sky130_fd_sc_hd__or3b_1
XFILLER_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3718_ _5186_/Q _3715_/X _3710_/X _3717_/Y vssd1 vssd1 vccd1 vccd1 _5186_/D sky130_fd_sc_hd__o211a_1
X_4698_ _4771_/A _4771_/B _4697_/X vssd1 vssd1 vccd1 vccd1 _4767_/B sky130_fd_sc_hd__a21oi_2
X_3649_ _5200_/Q _3613_/X _3646_/X _3648_/X vssd1 vssd1 vccd1 vccd1 _5200_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold12 phase_in[0] vssd1 vssd1 vccd1 vccd1 hold12/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_88_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold23 input8/X vssd1 vssd1 vccd1 vccd1 hold23/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_48_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold45 hold45/A vssd1 vssd1 vccd1 vccd1 hold45/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 hold34/A vssd1 vssd1 vccd1 vccd1 hold34/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_9 _4667_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2951_ _3650_/A vssd1 vssd1 vccd1 vccd1 _2951_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_34_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4621_ _5026_/Q _5058_/Q vssd1 vssd1 vccd1 vccd1 _4645_/A sky130_fd_sc_hd__nor2_1
X_2882_ _2903_/B _2882_/B vssd1 vssd1 vccd1 vccd1 _2882_/Y sky130_fd_sc_hd__nand2_1
X_4552_ _4434_/X _4548_/Y _4549_/X _4550_/X _4551_/Y vssd1 vssd1 vccd1 vccd1 _5058_/D
+ sky130_fd_sc_hd__o311a_1
X_3503_ _3511_/B _3503_/B vssd1 vssd1 vccd1 vccd1 _3504_/B sky130_fd_sc_hd__or2_1
X_4483_ _4483_/A _4483_/B vssd1 vssd1 vccd1 vccd1 _4483_/Y sky130_fd_sc_hd__nor2_1
X_3434_ _5225_/Q vssd1 vssd1 vccd1 vccd1 _3868_/B sky130_fd_sc_hd__inv_2
X_3365_ _3650_/A vssd1 vssd1 vccd1 vccd1 _3365_/X sky130_fd_sc_hd__buf_2
XFILLER_85_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5104_ _5109_/CLK _5104_/D vssd1 vssd1 vccd1 vccd1 _5104_/Q sky130_fd_sc_hd__dfxtp_1
X_3296_ _3289_/X _3295_/Y _2963_/X vssd1 vssd1 vccd1 vccd1 _3296_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5035_ _5040_/CLK _5035_/D vssd1 vssd1 vccd1 vccd1 _5035_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4819_ _3879_/X _4817_/Y _4807_/X _4818_/Y vssd1 vssd1 vccd1 vccd1 _5033_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput24 _5190_/Q vssd1 vssd1 vccd1 vccd1 data_out[0] sky130_fd_sc_hd__clkbuf_2
Xoutput46 _5192_/Q vssd1 vssd1 vccd1 vccd1 data_out[2] sky130_fd_sc_hd__clkbuf_2
Xoutput35 _5191_/Q vssd1 vssd1 vccd1 vccd1 data_out[1] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3150_ _3150_/A _3150_/B vssd1 vssd1 vccd1 vccd1 _3151_/A sky130_fd_sc_hd__nor2_2
XFILLER_67_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3081_ _5256_/Q vssd1 vssd1 vccd1 vccd1 _3787_/B sky130_fd_sc_hd__inv_2
XFILLER_39_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3983_ _4039_/A _4038_/A vssd1 vssd1 vccd1 vccd1 _3985_/A sky130_fd_sc_hd__nand2_1
X_2934_ _2940_/B _2940_/A vssd1 vssd1 vccd1 vccd1 _2936_/A sky130_fd_sc_hd__nand2_1
X_2865_ _2865_/A _2865_/B _2865_/C vssd1 vssd1 vccd1 vccd1 _2867_/A sky130_fd_sc_hd__or3_2
X_4604_ _4693_/B _4695_/B _4693_/A vssd1 vssd1 vccd1 vccd1 _4604_/X sky130_fd_sc_hd__o21ba_1
X_4535_ _4541_/B _4541_/A vssd1 vssd1 vccd1 vccd1 _4536_/A sky130_fd_sc_hd__or2_1
X_2796_ _2853_/B vssd1 vssd1 vccd1 vccd1 _2796_/Y sky130_fd_sc_hd__inv_2
X_4466_ _4742_/B _4594_/B _4462_/C _4465_/X vssd1 vssd1 vccd1 vccd1 _4467_/B sky130_fd_sc_hd__o22a_1
X_3417_ _3853_/B _5135_/Q vssd1 vssd1 vccd1 vccd1 _3455_/B sky130_fd_sc_hd__nand2_1
X_4397_ _4387_/A _4383_/A _4392_/Y _4396_/X vssd1 vssd1 vccd1 vccd1 _4427_/A sky130_fd_sc_hd__o211a_1
X_3348_ _3347_/B _3347_/A _3292_/X vssd1 vssd1 vccd1 vccd1 _3348_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3279_ _3284_/B _3284_/A vssd1 vssd1 vccd1 vccd1 _3279_/X sky130_fd_sc_hd__or2_1
X_5018_ _5114_/CLK _5018_/D vssd1 vssd1 vccd1 vccd1 _5018_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2650_ _4710_/A _5312_/Q vssd1 vssd1 vccd1 vccd1 _2651_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2581_ _5300_/Q _2567_/X _2563_/X _2580_/Y vssd1 vssd1 vccd1 vccd1 _5300_/D sky130_fd_sc_hd__o211a_1
X_4320_ _5061_/Q vssd1 vssd1 vccd1 vccd1 _4657_/B sky130_fd_sc_hd__inv_2
XFILLER_4_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4251_ _4254_/B vssd1 vssd1 vccd1 vccd1 _4251_/Y sky130_fd_sc_hd__inv_2
X_3202_ _4214_/A vssd1 vssd1 vccd1 vccd1 _3202_/X sky130_fd_sc_hd__clkbuf_4
X_4182_ _5094_/Q vssd1 vssd1 vccd1 vccd1 _4277_/A sky130_fd_sc_hd__inv_2
XFILLER_67_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3133_ _3133_/A _3133_/B vssd1 vssd1 vccd1 vccd1 _3281_/A sky130_fd_sc_hd__nor2_2
XFILLER_27_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3064_ _3064_/A _3064_/B vssd1 vssd1 vccd1 vccd1 _3064_/Y sky130_fd_sc_hd__nor2_1
XFILLER_63_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3966_ _5113_/Q _5112_/Q _5111_/Q vssd1 vssd1 vccd1 vccd1 _3967_/A sky130_fd_sc_hd__and3_1
XFILLER_10_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2917_ _2995_/A _3739_/B vssd1 vssd1 vccd1 vccd1 _2917_/Y sky130_fd_sc_hd__nand2_1
X_3897_ _5122_/Q vssd1 vssd1 vccd1 vccd1 _3898_/B sky130_fd_sc_hd__inv_2
XFILLER_12_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2848_ _3361_/A vssd1 vssd1 vccd1 vccd1 _2848_/X sky130_fd_sc_hd__buf_2
X_2779_ _5314_/Q _4592_/A vssd1 vssd1 vccd1 vccd1 _2843_/A sky130_fd_sc_hd__nor2_2
X_4518_ _4492_/X _5064_/Q _4516_/Y _4517_/X _4508_/X vssd1 vssd1 vccd1 vccd1 _5064_/D
+ sky130_fd_sc_hd__o221a_1
X_4449_ _4449_/A _4449_/B vssd1 vssd1 vccd1 vccd1 _4450_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3820_ _3820_/A _3820_/B vssd1 vssd1 vccd1 vccd1 _3820_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3751_ _5173_/Q _3741_/X _3749_/X _3750_/Y vssd1 vssd1 vccd1 vccd1 _5173_/D sky130_fd_sc_hd__o211a_1
X_2702_ _2801_/A _2702_/B vssd1 vssd1 vccd1 vccd1 _2799_/A sky130_fd_sc_hd__nand2_1
XFILLER_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3682_ _3673_/A _3681_/X _2951_/X vssd1 vssd1 vccd1 vccd1 _3682_/Y sky130_fd_sc_hd__o21ai_1
X_2633_ _2847_/A vssd1 vssd1 vccd1 vccd1 _3615_/A sky130_fd_sc_hd__clkbuf_2
X_2564_ _5037_/Q vssd1 vssd1 vccd1 vccd1 _4691_/A sky130_fd_sc_hd__inv_2
X_4303_ _5057_/Q vssd1 vssd1 vccd1 vccd1 _4643_/B sky130_fd_sc_hd__inv_2
X_5283_ _5283_/CLK _5283_/D vssd1 vssd1 vccd1 vccd1 _5283_/Q sky130_fd_sc_hd__dfxtp_1
X_4234_ _4234_/A _4234_/B vssd1 vssd1 vccd1 vccd1 _4235_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4165_ _4165_/A _4190_/B vssd1 vssd1 vccd1 vccd1 _4166_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3116_ _5169_/Q _3760_/B vssd1 vssd1 vccd1 vccd1 _3118_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4096_ _4202_/B _4094_/X _4095_/X _3967_/A _5114_/Q vssd1 vssd1 vccd1 vccd1 _4097_/C
+ sky130_fd_sc_hd__a41oi_1
X_3047_ _3047_/A _3047_/B vssd1 vssd1 vccd1 vccd1 _3047_/Y sky130_fd_sc_hd__nor2_1
XFILLER_82_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4998_ _5002_/CLK _4998_/D vssd1 vssd1 vccd1 vccd1 _4998_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3949_ _5107_/Q vssd1 vssd1 vccd1 vccd1 _4370_/A sky130_fd_sc_hd__inv_2
XFILLER_2_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4921_ _5124_/Q _5013_/Q vssd1 vssd1 vccd1 vccd1 _4921_/Y sky130_fd_sc_hd__nor2_1
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4852_ _4852_/A _4852_/B _4852_/C vssd1 vssd1 vccd1 vccd1 _4852_/X sky130_fd_sc_hd__and3_1
XFILLER_60_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3803_ _5154_/Q _3796_/X _3791_/X _3802_/Y vssd1 vssd1 vccd1 vccd1 _5154_/D sky130_fd_sc_hd__o211a_1
X_4783_ _4783_/A _4783_/B vssd1 vssd1 vccd1 vccd1 _4783_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3734_ _3739_/A _3734_/B vssd1 vssd1 vccd1 vccd1 _3734_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3665_ _3664_/B _3664_/A _3642_/X vssd1 vssd1 vccd1 vccd1 _3665_/X sky130_fd_sc_hd__a21o_1
X_2616_ _5023_/Q vssd1 vssd1 vccd1 vccd1 _4628_/A sky130_fd_sc_hd__inv_2
X_3596_ _3650_/A vssd1 vssd1 vccd1 vccd1 _3596_/X sky130_fd_sc_hd__clkbuf_2
X_2547_ _5309_/Q _2528_/X _2544_/X _2546_/Y vssd1 vssd1 vccd1 vccd1 _5309_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5266_ _5267_/CLK _5266_/D vssd1 vssd1 vccd1 vccd1 _5266_/Q sky130_fd_sc_hd__dfxtp_1
X_4217_ _4780_/B vssd1 vssd1 vccd1 vccd1 _4217_/X sky130_fd_sc_hd__clkbuf_2
X_5197_ _5197_/CLK _5197_/D vssd1 vssd1 vccd1 vccd1 _5197_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_18_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4148_ _4150_/A _4258_/A _4147_/Y vssd1 vssd1 vccd1 vccd1 _5104_/D sky130_fd_sc_hd__a21oi_1
X_4079_ _4181_/B _5094_/Q _5091_/Q vssd1 vssd1 vccd1 vccd1 _4165_/A sky130_fd_sc_hd__and3_1
XFILLER_43_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3450_ _3450_/A _3450_/B vssd1 vssd1 vccd1 vccd1 _3664_/A sky130_fd_sc_hd__or2_1
X_3381_ _3562_/B vssd1 vssd1 vccd1 vccd1 _3381_/Y sky130_fd_sc_hd__inv_2
X_5120_ _5120_/CLK _5120_/D vssd1 vssd1 vccd1 vccd1 _5120_/Q sky130_fd_sc_hd__dfxtp_1
X_5051_ _5085_/CLK _5051_/D vssd1 vssd1 vccd1 vccd1 _5051_/Q sky130_fd_sc_hd__dfxtp_1
X_4002_ _4984_/Q _4984_/D vssd1 vssd1 vccd1 vccd1 _4003_/B sky130_fd_sc_hd__and2_1
XFILLER_52_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4904_ _4906_/A hold23/X vssd1 vssd1 vccd1 vccd1 hold25/A sky130_fd_sc_hd__or2_1
XFILLER_60_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4835_ _4835_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4835_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4766_ _5044_/Q _4574_/X _4763_/Y _4765_/X _4584_/X vssd1 vssd1 vccd1 vccd1 _5044_/D
+ sky130_fd_sc_hd__o221a_1
X_3717_ _3726_/A _3717_/B vssd1 vssd1 vccd1 vccd1 _3717_/Y sky130_fd_sc_hd__nand2_1
X_4697_ _4779_/B _4697_/B _4775_/A vssd1 vssd1 vccd1 vccd1 _4697_/X sky130_fd_sc_hd__or3_1
X_3648_ _3640_/A _3647_/Y _3615_/X vssd1 vssd1 vccd1 vccd1 _3648_/X sky130_fd_sc_hd__a21o_1
X_3579_ _3578_/Y _3512_/Y _3494_/A _3508_/B vssd1 vssd1 vccd1 vccd1 _3586_/A sky130_fd_sc_hd__a31o_1
XFILLER_88_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold13 input6/X vssd1 vssd1 vccd1 vccd1 hold13/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 oversample_in[9] vssd1 vssd1 vccd1 vccd1 hold35/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 hold46/A vssd1 vssd1 vccd1 vccd1 hold46/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 oversample_in[6] vssd1 vssd1 vccd1 vccd1 input8/A sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _5250_/CLK _5249_/D vssd1 vssd1 vccd1 vccd1 _5249_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2950_ _2950_/A _2950_/B vssd1 vssd1 vccd1 vccd1 _2950_/Y sky130_fd_sc_hd__nor2_1
X_2881_ _2902_/A _2902_/B _2902_/C vssd1 vssd1 vccd1 vccd1 _2903_/B sky130_fd_sc_hd__a21o_1
XPHY_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4620_ _4620_/A vssd1 vssd1 vccd1 vccd1 _4821_/A sky130_fd_sc_hd__inv_2
X_4551_ _4572_/A _4623_/B vssd1 vssd1 vccd1 vccd1 _4551_/Y sky130_fd_sc_hd__nand2_1
X_3502_ _3815_/B _5149_/Q vssd1 vssd1 vccd1 vccd1 _3503_/B sky130_fd_sc_hd__and2_1
X_4482_ _4482_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _4483_/B sky130_fd_sc_hd__nand2_1
X_3433_ _5225_/Q _3425_/Y _3691_/A _3686_/B vssd1 vssd1 vccd1 vccd1 _3681_/A sky130_fd_sc_hd__o22ai_4
X_3364_ _5223_/Q _3321_/X _3360_/Y _3362_/X _3363_/X vssd1 vssd1 vccd1 vccd1 _5223_/D
+ sky130_fd_sc_hd__o221a_1
X_5103_ _5109_/CLK _5103_/D vssd1 vssd1 vccd1 vccd1 _5103_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3295_ _3295_/A _3295_/B vssd1 vssd1 vccd1 vccd1 _3295_/Y sky130_fd_sc_hd__nand2_1
X_5034_ _5303_/CLK _5034_/D vssd1 vssd1 vccd1 vccd1 _5034_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4818_ _4818_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4818_/Y sky130_fd_sc_hd__nand2_1
X_4749_ _5047_/Q _4574_/X _4747_/Y _4748_/X _4584_/X vssd1 vssd1 vccd1 vccd1 _5047_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_31_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput25 _5200_/Q vssd1 vssd1 vccd1 vccd1 data_out[10] sky130_fd_sc_hd__clkbuf_2
Xoutput36 _5210_/Q vssd1 vssd1 vccd1 vccd1 data_out[20] sky130_fd_sc_hd__clkbuf_2
Xoutput47 _5220_/Q vssd1 vssd1 vccd1 vccd1 data_out[30] sky130_fd_sc_hd__clkbuf_2
XFILLER_29_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3080_ _5161_/Q vssd1 vssd1 vccd1 vccd1 _3080_/Y sky130_fd_sc_hd__inv_2
X_3982_ _3981_/A _3981_/B _3981_/C vssd1 vssd1 vccd1 vccd1 _4038_/A sky130_fd_sc_hd__o21ai_2
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2933_ _2933_/A _2933_/B vssd1 vssd1 vccd1 vccd1 _2940_/B sky130_fd_sc_hd__nand2_1
X_2864_ _3721_/B _4968_/A vssd1 vssd1 vccd1 vccd1 _2864_/Y sky130_fd_sc_hd__nor2_1
X_2795_ _2827_/A _2793_/Y _3605_/A vssd1 vssd1 vccd1 vccd1 _2795_/Y sky130_fd_sc_hd__a21oi_1
X_4603_ _5040_/Q _5072_/Q vssd1 vssd1 vccd1 vccd1 _4693_/A sky130_fd_sc_hd__nor2_1
X_4534_ _4534_/A _4534_/B vssd1 vssd1 vccd1 vccd1 _4541_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4465_ _4460_/B _4460_/A _4542_/A vssd1 vssd1 vccd1 vccd1 _4465_/X sky130_fd_sc_hd__a21o_1
X_3416_ _5231_/Q vssd1 vssd1 vccd1 vccd1 _3853_/B sky130_fd_sc_hd__inv_2
X_4396_ _4444_/C _4444_/B _4396_/C vssd1 vssd1 vccd1 vccd1 _4396_/X sky130_fd_sc_hd__or3_2
X_3347_ _3347_/A _3347_/B vssd1 vssd1 vccd1 vccd1 _3347_/Y sky130_fd_sc_hd__nor2_1
XFILLER_85_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5017_ _5114_/CLK _5017_/D vssd1 vssd1 vccd1 vccd1 _5017_/Q sky130_fd_sc_hd__dfxtp_1
X_3278_ _3278_/A _3278_/B vssd1 vssd1 vccd1 vccd1 _3284_/A sky130_fd_sc_hd__nor2_1
XFILLER_26_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_83_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2580_ _2584_/A _4818_/A vssd1 vssd1 vccd1 vccd1 _2580_/Y sky130_fd_sc_hd__nand2_1
X_4250_ _4250_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _4254_/B sky130_fd_sc_hd__nor2_1
X_3201_ hold44/X vssd1 vssd1 vccd1 vccd1 _4214_/A sky130_fd_sc_hd__buf_2
X_4181_ _4185_/A _4181_/B vssd1 vssd1 vccd1 vccd1 _4181_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3132_ _3132_/A vssd1 vssd1 vccd1 vccd1 _3133_/B sky130_fd_sc_hd__inv_2
XFILLER_67_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3063_ _3143_/A _3142_/A _3143_/B vssd1 vssd1 vccd1 vccd1 _3063_/X sky130_fd_sc_hd__o21ba_1
XFILLER_23_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3965_ _4095_/A vssd1 vssd1 vccd1 vccd1 _4115_/B sky130_fd_sc_hd__inv_2
XFILLER_50_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3896_ _3887_/X _4972_/X _3893_/X _3895_/Y vssd1 vssd1 vccd1 vccd1 _5123_/D sky130_fd_sc_hd__o211a_1
X_2916_ _5273_/Q vssd1 vssd1 vccd1 vccd1 _3739_/B sky130_fd_sc_hd__inv_2
XFILLER_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2847_ _2847_/A vssd1 vssd1 vccd1 vccd1 _3361_/A sky130_fd_sc_hd__clkbuf_2
X_2778_ _2842_/B _5047_/Q _2814_/A _2777_/Y vssd1 vssd1 vccd1 vccd1 _2836_/A sky130_fd_sc_hd__o22ai_2
X_4517_ _4516_/B _4516_/A _4484_/X vssd1 vssd1 vccd1 vccd1 _4517_/X sky130_fd_sc_hd__a21o_1
X_4448_ _4454_/A _4454_/B _4378_/A vssd1 vssd1 vccd1 vccd1 _4449_/A sky130_fd_sc_hd__o21bai_1
X_4379_ _5077_/Q vssd1 vssd1 vccd1 vccd1 _4710_/B sky130_fd_sc_hd__inv_2
XFILLER_58_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3750_ _3752_/A _3750_/B vssd1 vssd1 vccd1 vccd1 _3750_/Y sky130_fd_sc_hd__nand2_1
X_2701_ _4643_/A _5292_/Q vssd1 vssd1 vccd1 vccd1 _2702_/B sky130_fd_sc_hd__nand2_1
X_3681_ _3681_/A _3681_/B _3685_/A vssd1 vssd1 vccd1 vccd1 _3681_/X sky130_fd_sc_hd__and3_1
XFILLER_64_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2632_ _2632_/A vssd1 vssd1 vccd1 vccd1 _2847_/A sky130_fd_sc_hd__inv_2
X_2563_ _2892_/A vssd1 vssd1 vccd1 vccd1 _2563_/X sky130_fd_sc_hd__clkbuf_2
X_4302_ _4302_/A _4302_/B vssd1 vssd1 vccd1 vccd1 _4546_/B sky130_fd_sc_hd__nor2_1
X_5282_ _5285_/CLK _5282_/D vssd1 vssd1 vccd1 vccd1 _5282_/Q sky130_fd_sc_hd__dfxtp_2
X_4233_ _4233_/A _4233_/B vssd1 vssd1 vccd1 vccd1 _4234_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4164_ _4164_/A vssd1 vssd1 vccd1 vccd1 _4168_/B sky130_fd_sc_hd__inv_2
XFILLER_55_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3115_ _5265_/Q vssd1 vssd1 vccd1 vccd1 _3760_/B sky130_fd_sc_hd__inv_2
X_4095_ _4095_/A vssd1 vssd1 vccd1 vccd1 _4095_/X sky130_fd_sc_hd__buf_1
XFILLER_82_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3046_ _3046_/A vssd1 vssd1 vccd1 vccd1 _3223_/A sky130_fd_sc_hd__inv_2
XFILLER_82_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4997_ _5001_/CLK hold3/X vssd1 vssd1 vccd1 vccd1 _4998_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_11_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3948_ _5108_/Q vssd1 vssd1 vccd1 vccd1 _4375_/A sky130_fd_sc_hd__inv_2
X_3879_ _3879_/A vssd1 vssd1 vccd1 vccd1 _3879_/X sky130_fd_sc_hd__buf_2
XFILLER_78_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4920_ _4920_/A _4920_/B _4920_/C vssd1 vssd1 vccd1 vccd1 _4927_/A sky130_fd_sc_hd__and3_1
XFILLER_64_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4851_ _4852_/A _4852_/C _4852_/B vssd1 vssd1 vccd1 vccd1 _4851_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3802_ _3807_/A _3802_/B vssd1 vssd1 vccd1 vccd1 _3802_/Y sky130_fd_sc_hd__nand2_1
X_4782_ _4695_/A _4787_/B _4695_/B vssd1 vssd1 vccd1 vccd1 _4783_/B sky130_fd_sc_hd__o21ba_1
X_3733_ _5180_/Q _3728_/X _3723_/X _3732_/Y vssd1 vssd1 vccd1 vccd1 _5180_/D sky130_fd_sc_hd__o211a_1
X_3664_ _3664_/A _3664_/B vssd1 vssd1 vccd1 vccd1 _3664_/Y sky130_fd_sc_hd__nor2_1
X_2615_ _5291_/Q _2604_/X _2600_/X _2614_/Y vssd1 vssd1 vccd1 vccd1 _5291_/D sky130_fd_sc_hd__o211a_1
X_3595_ _5210_/Q _3328_/X _3585_/X _3594_/X vssd1 vssd1 vccd1 vccd1 _5210_/D sky130_fd_sc_hd__o211a_1
X_2546_ _2546_/A _4597_/A vssd1 vssd1 vccd1 vccd1 _2546_/Y sky130_fd_sc_hd__nand2_1
X_5265_ _5267_/CLK _5265_/D vssd1 vssd1 vccd1 vccd1 _5265_/Q sky130_fd_sc_hd__dfxtp_1
X_5196_ _5196_/CLK _5196_/D vssd1 vssd1 vccd1 vccd1 _5196_/Q sky130_fd_sc_hd__dfxtp_1
X_4216_ _4417_/A vssd1 vssd1 vccd1 vccd1 _4780_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_28_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4147_ _4137_/A _4115_/C _3533_/X vssd1 vssd1 vccd1 vccd1 _4147_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_55_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4078_ _4321_/A _4315_/A vssd1 vssd1 vccd1 vccd1 _4181_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3029_ _5284_/Q _5188_/Q vssd1 vssd1 vccd1 vccd1 _3197_/A sky130_fd_sc_hd__nor2_2
XFILLER_24_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3380_ _3391_/B _3380_/B vssd1 vssd1 vccd1 vccd1 _3562_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5050_ _5112_/CLK _5050_/D vssd1 vssd1 vccd1 vccd1 _5050_/Q sky130_fd_sc_hd__dfxtp_1
X_4001_ _4984_/Q _4984_/D vssd1 vssd1 vccd1 vccd1 _4003_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4903_ _4906_/A hold19/X vssd1 vssd1 vccd1 vccd1 _5012_/D sky130_fd_sc_hd__or2_1
XFILLER_33_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4834_ _4834_/A _4834_/B _4834_/C vssd1 vssd1 vccd1 vccd1 _4834_/X sky130_fd_sc_hd__and3_1
X_4765_ _4763_/B _4763_/A _4764_/X vssd1 vssd1 vccd1 vccd1 _4765_/X sky130_fd_sc_hd__a21o_1
X_3716_ _3755_/A vssd1 vssd1 vccd1 vccd1 _3726_/A sky130_fd_sc_hd__clkbuf_2
X_4696_ _4783_/A _4787_/A vssd1 vssd1 vccd1 vccd1 _4697_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3647_ _3647_/A _3647_/B vssd1 vssd1 vccd1 vccd1 _3647_/Y sky130_fd_sc_hd__nand2_1
X_3578_ _3593_/B _3593_/A vssd1 vssd1 vccd1 vccd1 _3578_/Y sky130_fd_sc_hd__nand2_2
XFILLER_0_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5317_ _5317_/CLK _5317_/D vssd1 vssd1 vccd1 vccd1 _5317_/Q sky130_fd_sc_hd__dfxtp_1
X_2529_ _3769_/A vssd1 vssd1 vccd1 vccd1 _2605_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold14 oversample_in[4] vssd1 vssd1 vccd1 vccd1 input6/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold25 hold25/A vssd1 vssd1 vccd1 vccd1 hold25/X sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _5250_/CLK _5248_/D vssd1 vssd1 vccd1 vccd1 _5248_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold36 input3/X vssd1 vssd1 vccd1 vccd1 hold36/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_75_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5179_ _5179_/CLK _5179_/D vssd1 vssd1 vccd1 vccd1 _5179_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2880_ _5278_/Q _2625_/X _2619_/X _2879_/X vssd1 vssd1 vccd1 vccd1 _5278_/D sky130_fd_sc_hd__o211a_1
XPHY_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4550_ _4550_/A vssd1 vssd1 vccd1 vccd1 _4550_/X sky130_fd_sc_hd__buf_2
X_3501_ _5149_/Q _3815_/B vssd1 vssd1 vccd1 vccd1 _3511_/B sky130_fd_sc_hd__nor2_1
X_4481_ _4487_/B _4487_/A vssd1 vssd1 vccd1 vccd1 _4482_/A sky130_fd_sc_hd__nand2_1
X_3432_ _3871_/B _5128_/Q _3693_/A _3700_/B vssd1 vssd1 vccd1 vccd1 _3686_/B sky130_fd_sc_hd__a22oi_4
X_3363_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3363_/X sky130_fd_sc_hd__buf_2
X_5102_ _5109_/CLK _5102_/D vssd1 vssd1 vccd1 vccd1 _5102_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_85_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3294_ _5235_/Q _3269_/X _3291_/Y _3293_/X _3262_/X vssd1 vssd1 vccd1 vccd1 _5235_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5033_ _5303_/CLK _5033_/D vssd1 vssd1 vccd1 vccd1 _5033_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_25_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4817_ _4817_/A _4817_/B vssd1 vssd1 vccd1 vccd1 _4817_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_21_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4748_ _4747_/B _4747_/A _4484_/X vssd1 vssd1 vccd1 vccd1 _4748_/X sky130_fd_sc_hd__a21o_1
X_4679_ _5037_/Q _5069_/Q vssd1 vssd1 vccd1 vccd1 _4797_/A sky130_fd_sc_hd__xor2_2
Xoutput26 _5201_/Q vssd1 vssd1 vccd1 vccd1 data_out[11] sky130_fd_sc_hd__clkbuf_2
Xoutput37 _5211_/Q vssd1 vssd1 vccd1 vccd1 data_out[21] sky130_fd_sc_hd__clkbuf_2
Xoutput48 _5221_/Q vssd1 vssd1 vccd1 vccd1 data_out[31] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_71_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3981_ _3981_/A _3981_/B _3981_/C vssd1 vssd1 vccd1 vccd1 _4039_/A sky130_fd_sc_hd__or3_1
XFILLER_62_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2932_ _5270_/Q _2625_/X _2892_/X _2931_/X vssd1 vssd1 vccd1 vccd1 _5270_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5204_/CLK sky130_fd_sc_hd__clkbuf_16
X_2863_ _3650_/A vssd1 vssd1 vccd1 vccd1 _4968_/A sky130_fd_sc_hd__buf_2
X_2794_ _3615_/A vssd1 vssd1 vccd1 vccd1 _3605_/A sky130_fd_sc_hd__buf_2
X_4602_ _4788_/A _4602_/B vssd1 vssd1 vccd1 vccd1 _4695_/B sky130_fd_sc_hd__nor2_1
X_4533_ _4530_/X _5061_/Q _4473_/X _4532_/X vssd1 vssd1 vccd1 vccd1 _5061_/D sky130_fd_sc_hd__o211a_1
X_4464_ _4420_/X _5074_/Q _4461_/X _4463_/Y _4432_/X vssd1 vssd1 vccd1 vccd1 _5074_/D
+ sky130_fd_sc_hd__o221a_1
X_3415_ _5230_/Q vssd1 vssd1 vccd1 vccd1 _3855_/B sky130_fd_sc_hd__inv_2
X_4395_ _4395_/A _4395_/B vssd1 vssd1 vccd1 vccd1 _4444_/C sky130_fd_sc_hd__nand2_1
X_3346_ _3346_/A _3346_/B vssd1 vssd1 vccd1 vccd1 _3347_/B sky130_fd_sc_hd__or2_1
XFILLER_85_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5016_ _5114_/CLK _5016_/D vssd1 vssd1 vccd1 vccd1 _5016_/Q sky130_fd_sc_hd__dfxtp_1
X_3277_ _2901_/X _3274_/Y _3246_/X _3276_/Y vssd1 vssd1 vccd1 vccd1 _5238_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_33_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5236_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_0_clk/A sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_24_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 _5288_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_8_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4180_ _4180_/A _4180_/B _4180_/C vssd1 vssd1 vccd1 vccd1 _4185_/A sky130_fd_sc_hd__and3_1
X_3200_ _3542_/A _5252_/Q vssd1 vssd1 vccd1 vccd1 _3200_/Y sky130_fd_sc_hd__nand2_1
XFILLER_67_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3131_ _3750_/B _5173_/Q vssd1 vssd1 vccd1 vccd1 _3132_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3062_ _3745_/B _5175_/Q vssd1 vssd1 vccd1 vccd1 _3143_/B sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_15_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _4992_/CLK sky130_fd_sc_hd__clkbuf_16
X_3964_ _4100_/C _4127_/B vssd1 vssd1 vccd1 vccd1 _4095_/A sky130_fd_sc_hd__nor2_1
X_3895_ _4572_/A _4958_/B vssd1 vssd1 vccd1 vccd1 _3895_/Y sky130_fd_sc_hd__nand2_1
X_2915_ _4550_/A vssd1 vssd1 vccd1 vccd1 _2915_/X sky130_fd_sc_hd__buf_2
X_2846_ _2846_/A _2846_/B vssd1 vssd1 vccd1 vccd1 _2846_/Y sky130_fd_sc_hd__nor2_1
XFILLER_12_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2777_ _2853_/A _2853_/B _2776_/Y vssd1 vssd1 vccd1 vccd1 _2777_/Y sky130_fd_sc_hd__a21oi_2
X_4516_ _4516_/A _4516_/B vssd1 vssd1 vccd1 vccd1 _4516_/Y sky130_fd_sc_hd__nor2_1
X_4447_ _4445_/X _4446_/Y _4214_/X vssd1 vssd1 vccd1 vccd1 _5077_/D sky130_fd_sc_hd__a21oi_1
XFILLER_58_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4378_ _4378_/A _4450_/A vssd1 vssd1 vccd1 vccd1 _4390_/A sky130_fd_sc_hd__nor2_1
X_3329_ _3330_/B _3330_/A vssd1 vssd1 vccd1 vccd1 _3329_/X sky130_fd_sc_hd__or2_1
XFILLER_85_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2700_ _2700_/A _5025_/Q vssd1 vssd1 vccd1 vccd1 _2801_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3680_ _5195_/Q _3650_/X _3676_/X _3679_/Y _3644_/X vssd1 vssd1 vccd1 vccd1 _5195_/D
+ sky130_fd_sc_hd__o221a_1
X_2631_ _5020_/Q vssd1 vssd1 vccd1 vccd1 _4631_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2562_ _3315_/A vssd1 vssd1 vccd1 vccd1 _2892_/A sky130_fd_sc_hd__clkbuf_2
X_4301_ _4301_/A _4301_/B vssd1 vssd1 vccd1 vccd1 _4302_/B sky130_fd_sc_hd__nor2_1
X_5281_ _5283_/CLK _5281_/D vssd1 vssd1 vccd1 vccd1 _5281_/Q sky130_fd_sc_hd__dfxtp_1
X_4232_ _5083_/Q vssd1 vssd1 vccd1 vccd1 _4587_/B sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_4_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5040_/CLK sky130_fd_sc_hd__clkbuf_16
X_4163_ _5097_/Q vssd1 vssd1 vccd1 vccd1 _4337_/A sky130_fd_sc_hd__inv_2
XFILLER_28_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4094_ _4105_/A vssd1 vssd1 vccd1 vccd1 _4094_/X sky130_fd_sc_hd__clkbuf_2
X_3114_ _3300_/B _3114_/B vssd1 vssd1 vccd1 vccd1 _3305_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3045_ _3047_/B _3045_/B vssd1 vssd1 vccd1 vccd1 _3046_/A sky130_fd_sc_hd__nand2_1
XFILLER_82_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4996_ _5125_/CLK _4996_/D vssd1 vssd1 vccd1 vccd1 _4996_/Q sky130_fd_sc_hd__dfxtp_1
X_3947_ _5109_/Q vssd1 vssd1 vccd1 vccd1 _4382_/A sky130_fd_sc_hd__inv_2
XFILLER_23_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3878_ _4893_/A vssd1 vssd1 vccd1 vccd1 _3879_/A sky130_fd_sc_hd__buf_2
XFILLER_31_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2829_ _3542_/A _5284_/Q vssd1 vssd1 vccd1 vccd1 _2829_/Y sky130_fd_sc_hd__nand2_1
XFILLER_78_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4850_ _4855_/B _4855_/A vssd1 vssd1 vccd1 vccd1 _4852_/A sky130_fd_sc_hd__or2_1
XFILLER_45_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3801_ _5155_/Q _3796_/X _3791_/X _3800_/Y vssd1 vssd1 vccd1 vccd1 _5155_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4781_ _4778_/Y _4780_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _5041_/D sky130_fd_sc_hd__o21a_1
X_3732_ _3739_/A _3732_/B vssd1 vssd1 vccd1 vccd1 _3732_/Y sky130_fd_sc_hd__nand2_1
XFILLER_9_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3663_ _3663_/A _3663_/B vssd1 vssd1 vccd1 vccd1 _3664_/B sky130_fd_sc_hd__nand2_1
X_2614_ _2622_/A _4863_/A vssd1 vssd1 vccd1 vccd1 _2614_/Y sky130_fd_sc_hd__nand2_1
X_3594_ _3593_/X _3578_/Y _3306_/X vssd1 vssd1 vccd1 vccd1 _3594_/X sky130_fd_sc_hd__a21o_1
X_2545_ _5042_/Q vssd1 vssd1 vccd1 vccd1 _4597_/A sky130_fd_sc_hd__inv_2
X_5264_ _5267_/CLK _5264_/D vssd1 vssd1 vccd1 vccd1 _5264_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4215_ _4212_/Y _4213_/Y _4214_/X vssd1 vssd1 vccd1 vccd1 _5086_/D sky130_fd_sc_hd__a21oi_1
XFILLER_68_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5195_ _5195_/CLK _5195_/D vssd1 vssd1 vccd1 vccd1 _5195_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4146_ _4149_/A _4146_/B vssd1 vssd1 vccd1 vccd1 _4150_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4077_ _5092_/Q vssd1 vssd1 vccd1 vccd1 _4315_/A sky130_fd_sc_hd__inv_2
XFILLER_70_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3028_ _5284_/Q _5188_/Q vssd1 vssd1 vccd1 vccd1 _3197_/B sky130_fd_sc_hd__and2_1
XPHY_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4979_ _4928_/Y _4930_/B _4979_/S vssd1 vssd1 vccd1 vccd1 _4979_/X sky130_fd_sc_hd__mux2_1
XFILLER_3_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4000_ _4000_/A _4000_/B _4032_/A vssd1 vssd1 vccd1 vccd1 _4030_/A sky130_fd_sc_hd__nand3_4
XFILLER_65_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4902_ _4902_/A hold29/X vssd1 vssd1 vccd1 vccd1 _5013_/D sky130_fd_sc_hd__and2_1
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4833_ _4834_/A _4834_/C _4834_/B vssd1 vssd1 vccd1 vccd1 _4833_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_21_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4764_ _4764_/A vssd1 vssd1 vccd1 vccd1 _4764_/X sky130_fd_sc_hd__clkbuf_2
X_3715_ _3754_/A vssd1 vssd1 vccd1 vccd1 _3715_/X sky130_fd_sc_hd__clkbuf_2
X_4695_ _4695_/A _4695_/B vssd1 vssd1 vccd1 vccd1 _4787_/A sky130_fd_sc_hd__nor2_1
X_3646_ _3646_/A vssd1 vssd1 vccd1 vccd1 _3646_/X sky130_fd_sc_hd__clkbuf_2
X_3577_ _3577_/A vssd1 vssd1 vccd1 vccd1 _3593_/A sky130_fd_sc_hd__inv_2
XFILLER_0_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5316_ _5317_/CLK _5316_/D vssd1 vssd1 vccd1 vccd1 _5316_/Q sky130_fd_sc_hd__dfxtp_1
X_2528_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2528_/X sky130_fd_sc_hd__clkbuf_2
X_5247_ _5247_/CLK _5247_/D vssd1 vssd1 vccd1 vccd1 _5247_/Q sky130_fd_sc_hd__dfxtp_1
Xhold15 hold15/A vssd1 vssd1 vccd1 vccd1 hold15/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 hold37/A vssd1 vssd1 vccd1 vccd1 hold37/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 input5/X vssd1 vssd1 vccd1 vccd1 hold26/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_56_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5178_ _5179_/CLK _5178_/D vssd1 vssd1 vccd1 vccd1 _5178_/Q sky130_fd_sc_hd__dfxtp_1
X_4129_ _4119_/B _4115_/C _3533_/X vssd1 vssd1 vccd1 vccd1 _4129_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3500_ _5245_/Q vssd1 vssd1 vccd1 vccd1 _3815_/B sky130_fd_sc_hd__inv_2
X_4480_ _4359_/B _4499_/A _4361_/Y vssd1 vssd1 vccd1 vccd1 _4487_/B sky130_fd_sc_hd__o21ai_1
X_3431_ _5127_/Q _5223_/Q vssd1 vssd1 vccd1 vccd1 _3700_/B sky130_fd_sc_hd__or2b_2
X_3362_ _3367_/B _3360_/B _3361_/X vssd1 vssd1 vccd1 vccd1 _3362_/X sky130_fd_sc_hd__a21o_1
X_5101_ _5109_/CLK _5101_/D vssd1 vssd1 vccd1 vccd1 _5101_/Q sky130_fd_sc_hd__dfxtp_1
X_3293_ _3291_/B _3291_/A _3292_/X vssd1 vssd1 vccd1 vccd1 _3293_/X sky130_fd_sc_hd__a21o_1
X_5032_ _5062_/CLK _5032_/D vssd1 vssd1 vccd1 vccd1 _5032_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4816_ _4567_/X _4812_/Y _4813_/X _4550_/X _4815_/Y vssd1 vssd1 vccd1 vccd1 _5034_/D
+ sky130_fd_sc_hd__o311a_1
X_4747_ _4747_/A _4747_/B vssd1 vssd1 vccd1 vccd1 _4747_/Y sky130_fd_sc_hd__nor2_1
XFILLER_31_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4678_ _4691_/C _4678_/B vssd1 vssd1 vccd1 vccd1 _4794_/A sky130_fd_sc_hd__nor2_1
X_3629_ _3629_/A _3629_/B vssd1 vssd1 vccd1 vccd1 _3635_/A sky130_fd_sc_hd__and2_1
Xoutput27 _5202_/Q vssd1 vssd1 vccd1 vccd1 data_out[12] sky130_fd_sc_hd__clkbuf_2
Xoutput49 _5193_/Q vssd1 vssd1 vccd1 vccd1 data_out[3] sky130_fd_sc_hd__clkbuf_2
Xoutput38 _5212_/Q vssd1 vssd1 vccd1 vccd1 data_out[22] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_75_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3980_ _3980_/A _3980_/B vssd1 vssd1 vccd1 vccd1 _3981_/C sky130_fd_sc_hd__nor2_1
XFILLER_62_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2931_ _2926_/A _2930_/Y _2878_/X vssd1 vssd1 vccd1 vccd1 _2931_/X sky130_fd_sc_hd__a21o_1
XFILLER_43_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clkbuf_0_clk/X sky130_fd_sc_hd__clkbuf_16
XFILLER_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2862_ _2888_/A vssd1 vssd1 vccd1 vccd1 _3650_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4601_ _4601_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4693_/B sky130_fd_sc_hd__nor2_1
X_2793_ _2793_/A _2793_/B _2793_/C vssd1 vssd1 vccd1 vccd1 _2793_/Y sky130_fd_sc_hd__nor3_2
XFILLER_30_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4532_ _4527_/A _4531_/Y _4204_/X vssd1 vssd1 vccd1 vccd1 _4532_/X sky130_fd_sc_hd__a21o_1
X_4463_ _4463_/A _4912_/B vssd1 vssd1 vccd1 vccd1 _4463_/Y sky130_fd_sc_hd__nand2_1
X_3414_ _3472_/A _3470_/A _3628_/A vssd1 vssd1 vccd1 vccd1 _3618_/A sky130_fd_sc_hd__a21o_1
X_4394_ _4394_/A vssd1 vssd1 vccd1 vccd1 _4395_/B sky130_fd_sc_hd__inv_2
X_3345_ _3345_/A _3345_/B vssd1 vssd1 vccd1 vccd1 _3347_/A sky130_fd_sc_hd__nand2_1
X_3276_ _3276_/A _3833_/B vssd1 vssd1 vccd1 vccd1 _3276_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5015_ _5114_/CLK _5015_/D vssd1 vssd1 vccd1 vccd1 _5015_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3130_ _5173_/Q _3750_/B vssd1 vssd1 vccd1 vccd1 _3133_/A sky130_fd_sc_hd__nor2_2
XFILLER_79_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3061_ _5174_/Q _3747_/B vssd1 vssd1 vccd1 vccd1 _3142_/A sky130_fd_sc_hd__nor2_1
XFILLER_82_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3963_ _4131_/B vssd1 vssd1 vccd1 vccd1 _4127_/B sky130_fd_sc_hd__inv_2
XFILLER_50_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3894_ _5123_/Q vssd1 vssd1 vccd1 vccd1 _4958_/B sky130_fd_sc_hd__inv_2
XFILLER_31_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2914_ _2919_/A _2914_/B _2914_/C vssd1 vssd1 vccd1 vccd1 _2914_/X sky130_fd_sc_hd__and3_1
X_2845_ _2845_/A _2845_/B vssd1 vssd1 vccd1 vccd1 _2846_/B sky130_fd_sc_hd__nand2_1
X_2776_ _2776_/A _2854_/B vssd1 vssd1 vccd1 vccd1 _2776_/Y sky130_fd_sc_hd__nand2_1
X_4515_ _4520_/B _4520_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _4516_/B sky130_fd_sc_hd__o21ai_1
X_4446_ _4446_/A _5077_/Q vssd1 vssd1 vccd1 vccd1 _4446_/Y sky130_fd_sc_hd__nand2_1
X_4377_ _4377_/A vssd1 vssd1 vccd1 vccd1 _4450_/A sky130_fd_sc_hd__inv_2
X_3328_ _3613_/A vssd1 vssd1 vccd1 vccd1 _3328_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3259_ _3266_/B _3266_/A vssd1 vssd1 vccd1 vccd1 _3267_/A sky130_fd_sc_hd__or2_1
XFILLER_39_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2630_ _5288_/Q _2625_/X _2619_/X _2629_/Y vssd1 vssd1 vccd1 vccd1 _5288_/D sky130_fd_sc_hd__o211a_1
X_2561_ _5305_/Q _2548_/X _2544_/X _2560_/Y vssd1 vssd1 vccd1 vccd1 _5305_/D sky130_fd_sc_hd__o211a_1
X_4300_ _5086_/Q _5054_/Q _4556_/A _4559_/C _4559_/A vssd1 vssd1 vccd1 vccd1 _4546_/A
+ sky130_fd_sc_hd__o2111ai_4
X_5280_ _5280_/CLK _5280_/D vssd1 vssd1 vccd1 vccd1 _5280_/Q sky130_fd_sc_hd__dfxtp_1
X_4231_ _4229_/Y _4230_/Y _4214_/X vssd1 vssd1 vccd1 vccd1 _5084_/D sky130_fd_sc_hd__a21oi_1
XFILLER_4_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4162_ _4356_/A _4115_/C _4161_/Y vssd1 vssd1 vccd1 vccd1 _5099_/D sky130_fd_sc_hd__a21oi_1
XFILLER_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4093_ _4106_/A _4201_/C vssd1 vssd1 vccd1 vccd1 _4202_/B sky130_fd_sc_hd__nor2_4
X_3113_ _3763_/B _5168_/Q vssd1 vssd1 vccd1 vccd1 _3114_/B sky130_fd_sc_hd__nand2_1
X_3044_ _3721_/B _5184_/Q vssd1 vssd1 vccd1 vccd1 _3045_/B sky130_fd_sc_hd__nand2_1
XFILLER_63_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4995_ _5002_/CLK hold7/X vssd1 vssd1 vccd1 vccd1 _4996_/D sky130_fd_sc_hd__dfxtp_2
XFILLER_23_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3946_ _5110_/Q vssd1 vssd1 vccd1 vccd1 _4386_/A sky130_fd_sc_hd__inv_2
X_3877_ _4199_/A vssd1 vssd1 vccd1 vccd1 _4893_/A sky130_fd_sc_hd__buf_2
X_2828_ _3604_/A vssd1 vssd1 vccd1 vccd1 _3542_/A sky130_fd_sc_hd__buf_2
X_2759_ _4778_/B _5308_/Q vssd1 vssd1 vccd1 vccd1 _2760_/B sky130_fd_sc_hd__nand2_1
X_4429_ _4429_/A _4429_/B vssd1 vssd1 vccd1 vccd1 _4429_/X sky130_fd_sc_hd__or2_1
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_2_2_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_48_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_86_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3800_ _3807_/A _3800_/B vssd1 vssd1 vccd1 vccd1 _3800_/Y sky130_fd_sc_hd__nand2_1
X_4780_ _4780_/A _4780_/B _4780_/C vssd1 vssd1 vccd1 vccd1 _4780_/X sky130_fd_sc_hd__and3_1
XFILLER_60_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3731_ _5181_/Q _3728_/X _3723_/X _3730_/Y vssd1 vssd1 vccd1 vccd1 _5181_/D sky130_fd_sc_hd__o211a_1
X_3662_ _3860_/B _5132_/Q _3670_/A vssd1 vssd1 vccd1 vccd1 _3663_/A sky130_fd_sc_hd__a21o_1
X_2613_ _2698_/A vssd1 vssd1 vccd1 vccd1 _4863_/A sky130_fd_sc_hd__clkbuf_2
X_3593_ _3593_/A _3593_/B vssd1 vssd1 vccd1 vccd1 _3593_/X sky130_fd_sc_hd__or2_1
X_2544_ _4550_/A vssd1 vssd1 vccd1 vccd1 _2544_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_87_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5263_ _5267_/CLK _5263_/D vssd1 vssd1 vccd1 vccd1 _5263_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5194_ _5196_/CLK _5194_/D vssd1 vssd1 vccd1 vccd1 _5194_/Q sky130_fd_sc_hd__dfxtp_1
X_4214_ _4214_/A vssd1 vssd1 vccd1 vccd1 _4214_/X sky130_fd_sc_hd__buf_2
XFILLER_68_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4145_ _4365_/A _4145_/B vssd1 vssd1 vccd1 vccd1 _4146_/B sky130_fd_sc_hd__nor2_1
XFILLER_83_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4076_ _5093_/Q vssd1 vssd1 vccd1 vccd1 _4321_/A sky130_fd_sc_hd__inv_2
X_3027_ _3190_/A vssd1 vssd1 vccd1 vccd1 _3027_/Y sky130_fd_sc_hd__inv_2
XFILLER_24_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4978_ _4934_/X _4934_/B _4979_/S vssd1 vssd1 vccd1 vccd1 _4978_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3929_ _5123_/Q _4922_/B _5116_/Q _3927_/Y _3928_/X vssd1 vssd1 vccd1 vccd1 _3933_/A
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4901_ _4902_/A hold34/X vssd1 vssd1 vccd1 vccd1 _5014_/D sky130_fd_sc_hd__and2_1
XFILLER_18_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4832_ _4832_/A _4832_/B vssd1 vssd1 vccd1 vccd1 _4834_/B sky130_fd_sc_hd__nor2_1
XFILLER_60_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4763_ _4763_/A _4763_/B vssd1 vssd1 vccd1 vccd1 _4763_/Y sky130_fd_sc_hd__nor2_1
X_3714_ _5187_/Q _3668_/X _3710_/X _3713_/Y vssd1 vssd1 vccd1 vccd1 _5187_/D sky130_fd_sc_hd__o211a_1
X_4694_ _5039_/Q _5071_/Q vssd1 vssd1 vccd1 vccd1 _4695_/A sky130_fd_sc_hd__nor2_1
X_3645_ _5201_/Q _3596_/X _3641_/Y _3643_/X _3644_/X vssd1 vssd1 vccd1 vccd1 _5201_/D
+ sky130_fd_sc_hd__o221a_1
X_3576_ _3489_/X _3614_/A _3408_/Y vssd1 vssd1 vccd1 vccd1 _3593_/B sky130_fd_sc_hd__o21bai_1
XFILLER_0_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5315_ _5317_/CLK _5315_/D vssd1 vssd1 vccd1 vccd1 _5315_/Q sky130_fd_sc_hd__dfxtp_1
X_2527_ _3767_/A vssd1 vssd1 vccd1 vccd1 _2604_/A sky130_fd_sc_hd__buf_2
X_5246_ _5252_/CLK _5246_/D vssd1 vssd1 vccd1 vccd1 _5246_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold16 input7/X vssd1 vssd1 vccd1 vccd1 hold16/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 input2/X vssd1 vssd1 vccd1 vccd1 hold38/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 oversample_in[3] vssd1 vssd1 vccd1 vccd1 input5/A sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_68_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5177_ _5179_/CLK _5177_/D vssd1 vssd1 vccd1 vccd1 _5177_/Q sky130_fd_sc_hd__dfxtp_1
X_4128_ _4149_/A _4128_/B vssd1 vssd1 vccd1 vccd1 _4133_/A sky130_fd_sc_hd__nand2_1
X_4059_ _4059_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4060_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3430_ _5127_/Q _3873_/B _5222_/Q _3429_/Y vssd1 vssd1 vccd1 vccd1 _3693_/A sky130_fd_sc_hd__o2bb2ai_2
X_3361_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3361_/X sky130_fd_sc_hd__buf_2
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5100_ _5109_/CLK _5100_/D vssd1 vssd1 vccd1 vccd1 _5100_/Q sky130_fd_sc_hd__dfxtp_1
X_3292_ _3361_/A vssd1 vssd1 vccd1 vccd1 _3292_/X sky130_fd_sc_hd__clkbuf_2
X_5031_ _5303_/CLK _5031_/D vssd1 vssd1 vccd1 vccd1 _5031_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_80_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4815_ _4815_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4746_ _4746_/A _4746_/B vssd1 vssd1 vccd1 vccd1 _4747_/B sky130_fd_sc_hd__nand2_1
X_4677_ _4677_/A _4677_/B vssd1 vssd1 vccd1 vccd1 _4678_/B sky130_fd_sc_hd__nor2_1
X_3628_ _3628_/A _3628_/B vssd1 vssd1 vccd1 vccd1 _3632_/A sky130_fd_sc_hd__nor2_1
Xoutput28 _5203_/Q vssd1 vssd1 vccd1 vccd1 data_out[13] sky130_fd_sc_hd__clkbuf_2
Xoutput39 _5213_/Q vssd1 vssd1 vccd1 vccd1 data_out[23] sky130_fd_sc_hd__clkbuf_2
X_3559_ _3563_/A _3390_/Y _3391_/B _2878_/X vssd1 vssd1 vccd1 vccd1 _3559_/Y sky130_fd_sc_hd__a31oi_1
X_5229_ _5288_/CLK _5229_/D vssd1 vssd1 vccd1 vccd1 _5229_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_4_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _2930_/A _2930_/B vssd1 vssd1 vccd1 vccd1 _2930_/Y sky130_fd_sc_hd__nand2_1
XFILLER_50_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2861_ _5280_/Q vssd1 vssd1 vccd1 vccd1 _3721_/B sky130_fd_sc_hd__inv_2
X_4600_ _4779_/B _4775_/A vssd1 vssd1 vccd1 vccd1 _4600_/Y sky130_fd_sc_hd__nor2_2
XPHY_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2792_ _4968_/B _5317_/Q vssd1 vssd1 vccd1 vccd1 _2793_/C sky130_fd_sc_hd__and2_1
X_4531_ _4531_/A _4531_/B vssd1 vssd1 vccd1 vccd1 _4531_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4462_ _4462_/A _4462_/B _4462_/C vssd1 vssd1 vccd1 vccd1 _4463_/A sky130_fd_sc_hd__or3_2
X_3413_ _5139_/Q _3841_/B vssd1 vssd1 vccd1 vccd1 _3628_/A sky130_fd_sc_hd__nor2_1
X_4393_ _4375_/A _4704_/B _4449_/B vssd1 vssd1 vccd1 vccd1 _4395_/A sky130_fd_sc_hd__o21ai_1
X_3344_ _3785_/B _5161_/Q vssd1 vssd1 vccd1 vccd1 _3345_/B sky130_fd_sc_hd__nand2_1
X_3275_ _5238_/Q vssd1 vssd1 vccd1 vccd1 _3833_/B sky130_fd_sc_hd__inv_2
X_5014_ _5120_/CLK _5014_/D vssd1 vssd1 vccd1 vccd1 _5014_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4729_ _4735_/A _4735_/C _4735_/B vssd1 vssd1 vccd1 vccd1 _4736_/B sky130_fd_sc_hd__a21oi_1
XFILLER_1_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3060_ _5270_/Q vssd1 vssd1 vccd1 vccd1 _3747_/B sky130_fd_sc_hd__inv_2
XFILLER_35_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3962_ _3962_/A _4136_/B vssd1 vssd1 vccd1 vccd1 _4131_/B sky130_fd_sc_hd__and2_1
X_3893_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3893_/X sky130_fd_sc_hd__clkbuf_2
X_2913_ _2919_/A _2914_/C _2914_/B vssd1 vssd1 vccd1 vccd1 _2913_/Y sky130_fd_sc_hd__a21oi_1
X_2844_ _2844_/A vssd1 vssd1 vccd1 vccd1 _2846_/A sky130_fd_sc_hd__inv_2
XFILLER_12_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4514_ _4514_/A vssd1 vssd1 vccd1 vccd1 _4520_/A sky130_fd_sc_hd__inv_2
X_2775_ _2875_/A _2874_/B _2871_/C vssd1 vssd1 vccd1 vccd1 _2854_/B sky130_fd_sc_hd__and3_1
X_4445_ _4798_/A _4445_/B _4445_/C vssd1 vssd1 vccd1 vccd1 _4445_/X sky130_fd_sc_hd__or3_1
X_4376_ _4394_/A _4376_/B vssd1 vssd1 vccd1 vccd1 _4377_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3327_ _5229_/Q _3321_/X _3325_/Y _3326_/X _3316_/X vssd1 vssd1 vccd1 vccd1 _5229_/D
+ sky130_fd_sc_hd__o221a_1
X_3258_ _3145_/C _3274_/B _3063_/X vssd1 vssd1 vccd1 vccd1 _3266_/A sky130_fd_sc_hd__o21ba_1
XFILLER_37_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3189_ _3027_/Y _3199_/B _3190_/B _3190_/C vssd1 vssd1 vccd1 vccd1 _3189_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2560_ _2565_/A _4677_/A vssd1 vssd1 vccd1 vccd1 _2560_/Y sky130_fd_sc_hd__nand2_1
X_4230_ _4446_/A _4580_/A vssd1 vssd1 vccd1 vccd1 _4230_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4161_ _4356_/A _4115_/C _3533_/X vssd1 vssd1 vccd1 vccd1 _4161_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_67_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4092_ _4208_/D _4222_/A _4208_/B _4207_/A vssd1 vssd1 vccd1 vccd1 _4201_/C sky130_fd_sc_hd__a31oi_4
XFILLER_67_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3112_ _5168_/Q _3763_/B vssd1 vssd1 vccd1 vccd1 _3300_/B sky130_fd_sc_hd__or2_2
X_3043_ _5184_/Q _3721_/B vssd1 vssd1 vccd1 vccd1 _3047_/B sky130_fd_sc_hd__or2_2
XFILLER_36_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4994_ _5002_/CLK _4994_/D vssd1 vssd1 vccd1 vccd1 _4994_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3945_ _4214_/A vssd1 vssd1 vccd1 vccd1 _4116_/A sky130_fd_sc_hd__buf_2
XFILLER_23_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3876_ _5126_/Q _2841_/X _3870_/X _3875_/Y vssd1 vssd1 vccd1 vccd1 _5126_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2827_ _2827_/A _3563_/B _2827_/C vssd1 vssd1 vccd1 vccd1 _2827_/Y sky130_fd_sc_hd__nand3_1
X_2758_ _5308_/Q _4778_/B vssd1 vssd1 vccd1 vccd1 _2760_/A sky130_fd_sc_hd__or2_2
X_4428_ _4428_/A vssd1 vssd1 vccd1 vccd1 _4428_/Y sky130_fd_sc_hd__inv_2
X_2689_ _5288_/Q _4633_/A vssd1 vssd1 vccd1 vccd1 _3010_/A sky130_fd_sc_hd__nor2_4
XFILLER_58_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4359_ _4359_/A _4359_/B vssd1 vssd1 vccd1 vccd1 _4359_/Y sky130_fd_sc_hd__nor2_2
XFILLER_86_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3730_ _3739_/A _3730_/B vssd1 vssd1 vccd1 vccd1 _3730_/Y sky130_fd_sc_hd__nand2_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3661_ _3424_/Y _3673_/A _3442_/Y vssd1 vssd1 vccd1 vccd1 _3670_/A sky130_fd_sc_hd__o21ai_1
X_2612_ _5024_/Q vssd1 vssd1 vccd1 vccd1 _2698_/A sky130_fd_sc_hd__inv_2
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3592_ _5211_/Q _3365_/X _3589_/Y _3590_/X _3591_/X vssd1 vssd1 vccd1 vccd1 _5211_/D
+ sky130_fd_sc_hd__o221a_1
X_2543_ _5310_/Q _2528_/X _2522_/X _2542_/Y vssd1 vssd1 vccd1 vccd1 _5310_/D sky130_fd_sc_hd__o211a_1
X_5262_ _5267_/CLK _5262_/D vssd1 vssd1 vccd1 vccd1 _5262_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4213_ _4446_/A _5086_/Q vssd1 vssd1 vccd1 vccd1 _4213_/Y sky130_fd_sc_hd__nand2_1
X_5193_ _5195_/CLK _5193_/D vssd1 vssd1 vccd1 vccd1 _5193_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4144_ _4144_/A _4144_/B _4197_/B vssd1 vssd1 vccd1 vccd1 _5105_/D sky130_fd_sc_hd__and3_1
XFILLER_83_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4075_ _4091_/A vssd1 vssd1 vccd1 vccd1 _4180_/B sky130_fd_sc_hd__buf_2
X_3026_ _5188_/Q _3711_/B vssd1 vssd1 vccd1 vccd1 _3190_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4977_ _4938_/X _4938_/B _4979_/S vssd1 vssd1 vccd1 vccd1 _4977_/X sky130_fd_sc_hd__mux2_1
XFILLER_11_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3928_ _5008_/Q _3913_/B _4958_/B _5013_/Q vssd1 vssd1 vccd1 vccd1 _3928_/X sky130_fd_sc_hd__o22a_1
X_3859_ _5133_/Q _3849_/X _3857_/X _3858_/Y vssd1 vssd1 vccd1 vccd1 _5133_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4900_ _4902_/A hold40/X vssd1 vssd1 vccd1 vccd1 _5015_/D sky130_fd_sc_hd__and2_1
X_4831_ _4837_/B _4837_/A vssd1 vssd1 vccd1 vccd1 _4834_/A sky130_fd_sc_hd__or2_1
XFILLER_33_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_1_0_clk ANTENNA_10/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_2_1_0_clk/X sky130_fd_sc_hd__clkbuf_1
X_4762_ _4762_/A _4762_/B vssd1 vssd1 vccd1 vccd1 _4763_/B sky130_fd_sc_hd__nand2_1
XFILLER_33_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3713_ _3713_/A _3713_/B vssd1 vssd1 vccd1 vccd1 _3713_/Y sky130_fd_sc_hd__nand2_1
X_4693_ _4693_/A _4693_/B vssd1 vssd1 vccd1 vccd1 _4783_/A sky130_fd_sc_hd__nor2_1
X_3644_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3644_/X sky130_fd_sc_hd__clkbuf_2
X_3575_ _3575_/A _3575_/B vssd1 vssd1 vccd1 vccd1 _3614_/A sky130_fd_sc_hd__and2_1
X_5314_ _5317_/CLK _5314_/D vssd1 vssd1 vccd1 vccd1 _5314_/Q sky130_fd_sc_hd__dfxtp_1
X_2526_ _2888_/A vssd1 vssd1 vccd1 vccd1 _3767_/A sky130_fd_sc_hd__buf_1
X_5245_ _5252_/CLK _5245_/D vssd1 vssd1 vccd1 vccd1 _5245_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold17 oversample_in[5] vssd1 vssd1 vccd1 vccd1 input7/A sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 hold28/A vssd1 vssd1 vccd1 vccd1 hold28/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 hold39/A vssd1 vssd1 vccd1 vccd1 hold39/X sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ _5179_/CLK _5176_/D vssd1 vssd1 vccd1 vccd1 _5176_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4127_ _4370_/A _4127_/B vssd1 vssd1 vccd1 vccd1 _4128_/B sky130_fd_sc_hd__nor2_1
X_4058_ _5084_/Q vssd1 vssd1 vccd1 vccd1 _4580_/A sky130_fd_sc_hd__buf_2
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3009_ _3010_/A _3010_/B _3010_/C vssd1 vssd1 vccd1 vccd1 _3009_/X sky130_fd_sc_hd__o21a_1
XPHY_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3360_ _3367_/B _3360_/B vssd1 vssd1 vccd1 vccd1 _3360_/Y sky130_fd_sc_hd__nor2_1
X_5030_ _5301_/CLK _5030_/D vssd1 vssd1 vccd1 vccd1 _5030_/Q sky130_fd_sc_hd__dfxtp_1
X_3291_ _3291_/A _3291_/B vssd1 vssd1 vccd1 vccd1 _3291_/Y sky130_fd_sc_hd__nor2_1
XFILLER_38_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_45_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5197_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4814_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4872_/B sky130_fd_sc_hd__clkbuf_2
X_4745_ _4745_/A vssd1 vssd1 vccd1 vccd1 _4747_/A sky130_fd_sc_hd__inv_2
X_4676_ _5038_/Q _5070_/Q vssd1 vssd1 vccd1 vccd1 _4691_/C sky130_fd_sc_hd__nor2_1
X_3627_ _5204_/Q _3613_/X _3585_/X _3626_/X vssd1 vssd1 vccd1 vccd1 _5204_/D sky130_fd_sc_hd__o211a_1
X_3558_ _3563_/A _3391_/B _3390_/Y vssd1 vssd1 vccd1 vccd1 _3558_/X sky130_fd_sc_hd__a21o_1
Xoutput29 _5204_/Q vssd1 vssd1 vccd1 vccd1 data_out[14] sky130_fd_sc_hd__clkbuf_2
XFILLER_88_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2509_ _3843_/A vssd1 vssd1 vccd1 vccd1 _4807_/A sky130_fd_sc_hd__clkbuf_2
X_3489_ _3489_/A _3603_/B _3489_/C vssd1 vssd1 vccd1 vccd1 _3489_/X sky130_fd_sc_hd__or3_4
X_5228_ _5228_/CLK _5228_/D vssd1 vssd1 vccd1 vccd1 _5228_/Q sky130_fd_sc_hd__dfxtp_1
X_5159_ _5251_/CLK _5159_/D vssd1 vssd1 vccd1 vccd1 _5159_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_36_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5285_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_72_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 _5179_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2860_ _2634_/X _2856_/Y _2857_/X _2837_/X _2859_/Y vssd1 vssd1 vccd1 vccd1 _5281_/D
+ sky130_fd_sc_hd__o311a_1
XPHY_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2791_ _5317_/Q _4968_/B vssd1 vssd1 vccd1 vccd1 _2793_/B sky130_fd_sc_hd__nor2_2
XFILLER_7_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4530_ _4780_/B vssd1 vssd1 vccd1 vccd1 _4530_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_7_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4461_ _4462_/B _4462_/C _4462_/A vssd1 vssd1 vccd1 vccd1 _4461_/X sky130_fd_sc_hd__o21a_1
X_3412_ _3841_/B _5139_/Q vssd1 vssd1 vccd1 vccd1 _3470_/A sky130_fd_sc_hd__nand2_1
X_4392_ _4392_/A vssd1 vssd1 vccd1 vccd1 _4392_/Y sky130_fd_sc_hd__inv_2
X_3343_ _5226_/Q _3328_/X _3304_/X _3342_/Y vssd1 vssd1 vccd1 vccd1 _5226_/D sky130_fd_sc_hd__o211a_1
X_3274_ _3274_/A _3274_/B vssd1 vssd1 vccd1 vccd1 _3274_/Y sky130_fd_sc_hd__xnor2_1
X_5013_ _5120_/CLK _5013_/D vssd1 vssd1 vccd1 vccd1 _5013_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5301_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2989_ _2989_/A vssd1 vssd1 vccd1 vccd1 _2993_/A sky130_fd_sc_hd__inv_2
XFILLER_21_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4728_ _4728_/A _4728_/B vssd1 vssd1 vccd1 vccd1 _4735_/B sky130_fd_sc_hd__or2_1
X_4659_ _4832_/B _4832_/A _4837_/B vssd1 vssd1 vccd1 vccd1 _4659_/X sky130_fd_sc_hd__or3_1
XFILLER_1_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3961_ _4258_/A _4365_/A vssd1 vssd1 vccd1 vccd1 _4136_/B sky130_fd_sc_hd__nor2_1
XFILLER_90_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2912_ _2909_/X _2910_/Y _2911_/Y vssd1 vssd1 vccd1 vccd1 _2919_/A sky130_fd_sc_hd__a21o_1
X_3892_ _3887_/X _4971_/X _3870_/X _3891_/Y vssd1 vssd1 vccd1 vccd1 _5124_/D sky130_fd_sc_hd__o211a_1
XFILLER_31_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2843_ _2843_/A _2843_/B vssd1 vssd1 vccd1 vccd1 _2844_/A sky130_fd_sc_hd__nor2_1
XFILLER_31_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2774_ _4701_/A _5310_/Q vssd1 vssd1 vccd1 vccd1 _2871_/C sky130_fd_sc_hd__nand2_1
X_4513_ _4513_/A _4513_/B vssd1 vssd1 vccd1 vccd1 _4514_/A sky130_fd_sc_hd__or2_1
XFILLER_7_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4444_ _4444_/A _4444_/B _4444_/C vssd1 vssd1 vccd1 vccd1 _4445_/B sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_7_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5096_/CLK sky130_fd_sc_hd__clkbuf_16
X_4375_ _4375_/A _4704_/B vssd1 vssd1 vccd1 vccd1 _4376_/B sky130_fd_sc_hd__nor2_1
X_3326_ _3325_/B _3325_/A _3292_/X vssd1 vssd1 vccd1 vccd1 _3326_/X sky130_fd_sc_hd__a21o_1
X_3257_ _3257_/A _3257_/B vssd1 vssd1 vccd1 vccd1 _3274_/B sky130_fd_sc_hd__and2_1
XFILLER_54_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3188_ _3707_/B _5189_/Q vssd1 vssd1 vccd1 vccd1 _3190_/C sky130_fd_sc_hd__and2_1
XFILLER_54_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4160_ _4734_/A _4160_/B _4160_/C vssd1 vssd1 vccd1 vccd1 _5100_/D sky130_fd_sc_hd__nor3_1
XFILLER_4_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3111_ _5264_/Q vssd1 vssd1 vccd1 vccd1 _3763_/B sky130_fd_sc_hd__inv_2
X_4091_ _4091_/A vssd1 vssd1 vccd1 vccd1 _4106_/A sky130_fd_sc_hd__inv_2
X_3042_ _3042_/A _3047_/A vssd1 vssd1 vccd1 vccd1 _3172_/B sky130_fd_sc_hd__nor2_2
XFILLER_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4993_ _5002_/CLK hold9/X vssd1 vssd1 vccd1 vccd1 _4994_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3944_ _3907_/X _4979_/S _3911_/X _3943_/Y vssd1 vssd1 vccd1 vccd1 _5115_/D sky130_fd_sc_hd__o211a_1
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3875_ _4968_/A _3875_/B vssd1 vssd1 vccd1 vccd1 _3875_/Y sky130_fd_sc_hd__nand2_1
X_2826_ _2787_/Y _2826_/B _2826_/C vssd1 vssd1 vccd1 vccd1 _2827_/C sky130_fd_sc_hd__nand3b_1
X_2757_ _5309_/Q _4597_/A vssd1 vssd1 vccd1 vccd1 _2885_/A sky130_fd_sc_hd__nor2_2
X_2688_ _5289_/Q vssd1 vssd1 vccd1 vccd1 _3000_/B sky130_fd_sc_hd__inv_2
X_4427_ _4427_/A vssd1 vssd1 vccd1 vccd1 _4427_/Y sky130_fd_sc_hd__inv_2
XFILLER_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4358_ _4494_/A _4494_/B _4499_/B vssd1 vssd1 vccd1 vccd1 _4359_/B sky130_fd_sc_hd__or3_1
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4289_ _4289_/A _4628_/B vssd1 vssd1 vccd1 vccd1 _4291_/A sky130_fd_sc_hd__nand2_1
X_3309_ _3309_/A vssd1 vssd1 vccd1 vccd1 _3313_/A sky130_fd_sc_hd__inv_2
XFILLER_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3660_ _5198_/Q _3613_/X _3646_/X _3659_/X vssd1 vssd1 vccd1 vccd1 _5198_/D sky130_fd_sc_hd__o211a_1
X_2611_ _5292_/Q _2604_/X _2600_/X _2610_/Y vssd1 vssd1 vccd1 vccd1 _5292_/D sky130_fd_sc_hd__o211a_1
X_3591_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3591_/X sky130_fd_sc_hd__clkbuf_2
X_2542_ _2546_/A _4701_/A vssd1 vssd1 vccd1 vccd1 _2542_/Y sky130_fd_sc_hd__nand2_1
X_5261_ _5267_/CLK _5261_/D vssd1 vssd1 vccd1 vccd1 _5261_/Q sky130_fd_sc_hd__dfxtp_1
X_4212_ _4208_/X _4778_/A _4212_/C vssd1 vssd1 vccd1 vccd1 _4212_/Y sky130_fd_sc_hd__nand3b_1
X_5192_ _5195_/CLK _5192_/D vssd1 vssd1 vccd1 vccd1 _5192_/Q sky130_fd_sc_hd__dfxtp_1
X_4143_ _4807_/A vssd1 vssd1 vccd1 vccd1 _4197_/B sky130_fd_sc_hd__clkbuf_4
XFILLER_68_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4074_ _4417_/A _5088_/Q _5087_/Q vssd1 vssd1 vccd1 vccd1 _4091_/A sky130_fd_sc_hd__and3_1
XFILLER_83_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3025_ _5284_/Q vssd1 vssd1 vccd1 vccd1 _3711_/B sky130_fd_sc_hd__inv_2
XFILLER_83_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4976_ _4942_/X _4942_/B _4979_/S vssd1 vssd1 vccd1 vccd1 _4976_/X sky130_fd_sc_hd__mux2_1
X_3927_ _5006_/Q vssd1 vssd1 vccd1 vccd1 _3927_/Y sky130_fd_sc_hd__inv_2
X_3858_ _3860_/A _3858_/B vssd1 vssd1 vccd1 vccd1 _3858_/Y sky130_fd_sc_hd__nand2_1
X_3789_ _3794_/A _3789_/B vssd1 vssd1 vccd1 vccd1 _3789_/Y sky130_fd_sc_hd__nand2_1
X_2809_ _2933_/A _2933_/B _2743_/Y vssd1 vssd1 vccd1 vccd1 _2908_/B sky130_fd_sc_hd__a21oi_2
XFILLER_59_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4830_ _4830_/A _4830_/B vssd1 vssd1 vccd1 vccd1 _4837_/A sky130_fd_sc_hd__and2_1
XFILLER_33_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4761_ _4761_/A _4750_/X vssd1 vssd1 vccd1 vccd1 _4762_/A sky130_fd_sc_hd__or2b_1
X_3712_ _5188_/Q _3668_/X _3710_/X _3711_/Y vssd1 vssd1 vccd1 vccd1 _5188_/D sky130_fd_sc_hd__o211a_1
X_4692_ _4677_/A _4677_/B _4690_/Y _4688_/A _4691_/X vssd1 vssd1 vccd1 vccd1 _4771_/B
+ sky130_fd_sc_hd__o221a_1
X_3643_ _3641_/B _3641_/A _3642_/X vssd1 vssd1 vccd1 vccd1 _3643_/X sky130_fd_sc_hd__a21o_1
X_3574_ _5214_/Q _3328_/X _3304_/X _3573_/Y vssd1 vssd1 vccd1 vccd1 _5214_/D sky130_fd_sc_hd__o211a_1
X_5313_ _5317_/CLK _5313_/D vssd1 vssd1 vccd1 vccd1 _5313_/Q sky130_fd_sc_hd__dfxtp_1
X_2525_ _5314_/Q _2506_/X _2522_/X _2524_/Y vssd1 vssd1 vccd1 vccd1 _5314_/D sky130_fd_sc_hd__o211a_1
X_5244_ _5252_/CLK _5244_/D vssd1 vssd1 vccd1 vccd1 _5244_/Q sky130_fd_sc_hd__dfxtp_1
Xhold29 hold29/A vssd1 vssd1 vccd1 vccd1 hold29/X sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 hold18/A vssd1 vssd1 vccd1 vccd1 hold18/X sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _5179_/CLK _5175_/D vssd1 vssd1 vccd1 vccd1 _5175_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4126_ _4126_/A vssd1 vssd1 vccd1 vccd1 _4149_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_83_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4057_ _4057_/A _4057_/B vssd1 vssd1 vccd1 vccd1 _4057_/Y sky130_fd_sc_hd__nor2_2
XFILLER_24_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3008_ _3008_/A _3018_/B vssd1 vssd1 vccd1 vccd1 _3010_/C sky130_fd_sc_hd__nand2_1
XPHY_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4959_ _4962_/B _4960_/C vssd1 vssd1 vccd1 vccd1 _4959_/X sky130_fd_sc_hd__and2_1
XFILLER_24_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_87_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3290_ _3758_/B _5170_/Q _3289_/X vssd1 vssd1 vccd1 vccd1 _3291_/B sky130_fd_sc_hd__o21a_1
XFILLER_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_65_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4813_ _4813_/A _4813_/B vssd1 vssd1 vccd1 vccd1 _4813_/X sky130_fd_sc_hd__and2_1
X_4744_ _4744_/A _4744_/B vssd1 vssd1 vccd1 vccd1 _4745_/A sky130_fd_sc_hd__nor2_1
X_4675_ _4810_/A _4810_/B _4674_/Y vssd1 vssd1 vccd1 vccd1 _4790_/B sky130_fd_sc_hd__a21oi_2
X_3626_ _3622_/A _3625_/Y _3615_/X vssd1 vssd1 vccd1 vccd1 _3626_/X sky130_fd_sc_hd__a21o_1
X_3557_ _3562_/A _3381_/Y vssd1 vssd1 vccd1 vccd1 _3563_/A sky130_fd_sc_hd__or2b_1
X_2508_ _2821_/A vssd1 vssd1 vccd1 vccd1 _3843_/A sky130_fd_sc_hd__buf_2
X_3488_ _3608_/B _3608_/A _3614_/B vssd1 vssd1 vccd1 vccd1 _3489_/C sky130_fd_sc_hd__or3_1
X_5227_ _5274_/CLK _5227_/D vssd1 vssd1 vccd1 vccd1 _5227_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_69_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5158_ _5251_/CLK _5158_/D vssd1 vssd1 vccd1 vccd1 _5158_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5089_ _5118_/CLK _5089_/D vssd1 vssd1 vccd1 vccd1 _5089_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4109_ _4127_/B _4101_/B _4119_/C _2889_/X vssd1 vssd1 vccd1 vccd1 _4110_/B sky130_fd_sc_hd__o31ai_1
XFILLER_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_2_0_0_clk ANTENNA_10/DIODE vssd1 vssd1 vccd1 vccd1 clkbuf_2_0_0_clk/X sky130_fd_sc_hd__clkbuf_1
XFILLER_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2790_ _5050_/Q vssd1 vssd1 vccd1 vccd1 _4968_/B sky130_fd_sc_hd__inv_2
XFILLER_30_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4460_ _4460_/A _4460_/B vssd1 vssd1 vccd1 vccd1 _4462_/C sky130_fd_sc_hd__nor2_1
X_3411_ _5235_/Q vssd1 vssd1 vccd1 vccd1 _3841_/B sky130_fd_sc_hd__inv_2
XFILLER_7_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4391_ _4454_/A _4454_/B _4390_/Y vssd1 vssd1 vccd1 vccd1 _4428_/A sky130_fd_sc_hd__o21bai_2
X_3342_ _3333_/A _3341_/X _2951_/X vssd1 vssd1 vccd1 vccd1 _3342_/Y sky130_fd_sc_hd__o21ai_2
X_3273_ _5239_/Q _3269_/X _3271_/Y _3272_/X _3262_/X vssd1 vssd1 vccd1 vccd1 _5239_/D
+ sky130_fd_sc_hd__o221a_1
X_5012_ _5120_/CLK _5012_/D vssd1 vssd1 vccd1 vccd1 _5012_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2988_ _2901_/X _2985_/Y _2961_/X _2987_/Y vssd1 vssd1 vccd1 vccd1 _5260_/D sky130_fd_sc_hd__o211a_1
X_4727_ _5049_/Q _5081_/Q vssd1 vssd1 vccd1 vccd1 _4728_/A sky130_fd_sc_hd__nor2_1
X_4658_ _4658_/A _4834_/C vssd1 vssd1 vccd1 vccd1 _4837_/B sky130_fd_sc_hd__nand2_1
X_3609_ _3610_/A _3611_/A _3610_/B _2897_/X vssd1 vssd1 vccd1 vccd1 _3609_/X sky130_fd_sc_hd__a31o_1
X_4589_ _4589_/A vssd1 vssd1 vccd1 vccd1 _4906_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_67_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3960_ _5103_/Q vssd1 vssd1 vccd1 vccd1 _4365_/A sky130_fd_sc_hd__inv_2
XFILLER_90_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_opt_0_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 clkbuf_opt_0_clk/X sky130_fd_sc_hd__clkbuf_16
X_2911_ _2914_/C _2911_/B vssd1 vssd1 vccd1 vccd1 _2911_/Y sky130_fd_sc_hd__nand2_1
X_3891_ _4572_/A _4962_/A vssd1 vssd1 vccd1 vccd1 _3891_/Y sky130_fd_sc_hd__nand2_1
XFILLER_85_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2842_ _5047_/Q _2842_/B vssd1 vssd1 vccd1 vccd1 _2843_/B sky130_fd_sc_hd__nor2_1
X_2773_ _5310_/Q _4701_/A vssd1 vssd1 vccd1 vccd1 _2874_/B sky130_fd_sc_hd__or2_2
X_4512_ _4453_/X _5065_/Q _4473_/X _4511_/X vssd1 vssd1 vccd1 vccd1 _5065_/D sky130_fd_sc_hd__o211a_1
X_4443_ _4893_/A vssd1 vssd1 vccd1 vccd1 _4798_/A sky130_fd_sc_hd__clkbuf_2
X_4374_ _5076_/Q vssd1 vssd1 vccd1 vccd1 _4704_/B sky130_fd_sc_hd__inv_2
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3325_ _3325_/A _3325_/B vssd1 vssd1 vccd1 vccd1 _3325_/Y sky130_fd_sc_hd__nor2_1
X_3256_ _5242_/Q _3253_/X _3246_/X _3255_/X vssd1 vssd1 vccd1 vccd1 _5242_/D sky130_fd_sc_hd__o211a_1
XFILLER_37_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3187_ _5189_/Q _3707_/B vssd1 vssd1 vccd1 vccd1 _3190_/B sky130_fd_sc_hd__nor2_1
XFILLER_54_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_78_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3110_ _3310_/A _3310_/B _3109_/X vssd1 vssd1 vccd1 vccd1 _3298_/B sky130_fd_sc_hd__a21oi_2
XFILLER_67_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4090_ _4115_/B _4090_/B _4119_/C vssd1 vssd1 vccd1 vccd1 _4097_/B sky130_fd_sc_hd__nor3_2
X_3041_ _3719_/B _5185_/Q vssd1 vssd1 vccd1 vccd1 _3047_/A sky130_fd_sc_hd__and2_1
XFILLER_48_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4992_ _4992_/CLK _4992_/D vssd1 vssd1 vccd1 vccd1 _4992_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_51_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3943_ _4446_/A _4911_/B vssd1 vssd1 vccd1 vccd1 _3943_/Y sky130_fd_sc_hd__nand2_1
X_3874_ _5127_/Q _3862_/X _3870_/X _3873_/Y vssd1 vssd1 vccd1 vccd1 _5127_/D sky130_fd_sc_hd__o211a_1
X_2825_ _3011_/A vssd1 vssd1 vccd1 vccd1 _3563_/B sky130_fd_sc_hd__buf_2
X_2756_ _4597_/A _5309_/Q vssd1 vssd1 vccd1 vccd1 _2885_/B sky130_fd_sc_hd__and2_1
X_2687_ _5291_/Q _4863_/A _2993_/B vssd1 vssd1 vccd1 vccd1 _2687_/Y sky130_fd_sc_hd__o21ai_2
X_4426_ _4420_/X _4739_/B _4422_/X _4425_/Y _3695_/X vssd1 vssd1 vccd1 vccd1 _5080_/D
+ sky130_fd_sc_hd__o221a_1
X_4357_ _4496_/B _4357_/B vssd1 vssd1 vccd1 vccd1 _4499_/B sky130_fd_sc_hd__nand2_1
X_4288_ _5055_/Q vssd1 vssd1 vccd1 vccd1 _4628_/B sky130_fd_sc_hd__inv_2
X_3308_ _5232_/Q _3253_/X _3304_/X _3307_/X vssd1 vssd1 vccd1 vccd1 _5232_/D sky130_fd_sc_hd__o211a_1
X_3239_ _3164_/A _3238_/Y _3170_/Y vssd1 vssd1 vccd1 vccd1 _3247_/A sky130_fd_sc_hd__o21a_1
XFILLER_39_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2610_ _2622_/A _4643_/A vssd1 vssd1 vccd1 vccd1 _2610_/Y sky130_fd_sc_hd__nand2_1
X_3590_ _3578_/Y _3508_/Y _3494_/A _3604_/A vssd1 vssd1 vccd1 vccd1 _3590_/X sky130_fd_sc_hd__a31o_1
X_2541_ _4699_/A vssd1 vssd1 vccd1 vccd1 _4701_/A sky130_fd_sc_hd__buf_1
X_5260_ _5267_/CLK _5260_/D vssd1 vssd1 vccd1 vccd1 _5260_/Q sky130_fd_sc_hd__dfxtp_1
X_4211_ _4222_/A _4208_/D _4208_/A _4208_/B vssd1 vssd1 vccd1 vccd1 _4212_/C sky130_fd_sc_hd__a22o_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5191_ _5195_/CLK _5191_/D vssd1 vssd1 vccd1 vccd1 _5191_/Q sky130_fd_sc_hd__dfxtp_1
X_4142_ _4137_/A _4119_/C _4252_/A vssd1 vssd1 vccd1 vccd1 _4144_/A sky130_fd_sc_hd__o21ai_1
X_4073_ _5015_/Q vssd1 vssd1 vccd1 vccd1 _4417_/A sky130_fd_sc_hd__buf_2
XFILLER_83_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3024_ _5254_/Q _2977_/X _3022_/Y _3023_/Y _2971_/X vssd1 vssd1 vccd1 vccd1 _5254_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_48_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4975_ _4947_/X _4947_/B _4979_/S vssd1 vssd1 vccd1 vccd1 _4975_/X sky130_fd_sc_hd__mux2_1
X_3926_ _5013_/Q vssd1 vssd1 vccd1 vccd1 _4922_/B sky130_fd_sc_hd__inv_2
X_3857_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3857_/X sky130_fd_sc_hd__clkbuf_2
X_3788_ _5160_/Q _3783_/X _3778_/X _3787_/Y vssd1 vssd1 vccd1 vccd1 _5160_/D sky130_fd_sc_hd__o211a_1
X_2808_ _2808_/A vssd1 vssd1 vccd1 vccd1 _2933_/B sky130_fd_sc_hd__inv_2
X_2739_ _2739_/A _5033_/Q vssd1 vssd1 vccd1 vccd1 _2936_/B sky130_fd_sc_hd__nand2_1
XFILLER_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4409_ _4241_/Y _4407_/Y _4411_/C vssd1 vssd1 vccd1 vccd1 _4412_/A sky130_fd_sc_hd__o21bai_1
XFILLER_46_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4760_ _4758_/X _4759_/Y _4116_/A vssd1 vssd1 vccd1 vccd1 _5045_/D sky130_fd_sc_hd__a21oi_1
X_3711_ _3713_/A _3711_/B vssd1 vssd1 vccd1 vccd1 _3711_/Y sky130_fd_sc_hd__nand2_1
X_4691_ _4691_/A _4691_/B _4691_/C vssd1 vssd1 vccd1 vccd1 _4691_/X sky130_fd_sc_hd__or3_2
X_3642_ _3642_/A vssd1 vssd1 vccd1 vccd1 _3642_/X sky130_fd_sc_hd__buf_2
X_3573_ _3572_/X _3568_/B _2951_/X vssd1 vssd1 vccd1 vccd1 _3573_/Y sky130_fd_sc_hd__o21ai_1
X_5312_ _5317_/CLK _5312_/D vssd1 vssd1 vccd1 vccd1 _5312_/Q sky130_fd_sc_hd__dfxtp_1
X_2524_ _2524_/A _4592_/A vssd1 vssd1 vccd1 vccd1 _2524_/Y sky130_fd_sc_hd__nand2_1
X_5243_ _5274_/CLK _5243_/D vssd1 vssd1 vccd1 vccd1 _5243_/Q sky130_fd_sc_hd__dfxtp_1
Xhold19 input9/X vssd1 vssd1 vccd1 vccd1 hold19/X sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ _5179_/CLK _5174_/D vssd1 vssd1 vccd1 vccd1 _5174_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4125_ _4734_/A _4125_/B _4125_/C vssd1 vssd1 vccd1 vccd1 _5109_/D sky130_fd_sc_hd__nor3_1
XFILLER_83_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4056_ _4056_/A _4056_/B _4056_/C vssd1 vssd1 vccd1 vccd1 _4057_/B sky130_fd_sc_hd__nand3_2
X_3007_ _3007_/A vssd1 vssd1 vccd1 vccd1 _3010_/B sky130_fd_sc_hd__inv_2
XPHY_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4958_ _4958_/A _4958_/B vssd1 vssd1 vccd1 vccd1 _4960_/C sky130_fd_sc_hd__nand2_1
X_3909_ _3916_/A _4940_/A vssd1 vssd1 vccd1 vccd1 _3909_/Y sky130_fd_sc_hd__nand2_1
X_4889_ _4898_/A _4892_/A _4898_/B vssd1 vssd1 vccd1 vccd1 _4891_/A sky130_fd_sc_hd__or3_1
XFILLER_10_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4812_ _4813_/B _4813_/A vssd1 vssd1 vccd1 vccd1 _4812_/Y sky130_fd_sc_hd__nor2_1
X_4743_ _4739_/A _4574_/X _4740_/X _4742_/Y _4584_/X vssd1 vssd1 vccd1 vccd1 _5048_/D
+ sky130_fd_sc_hd__o221a_1
X_4674_ _4813_/B _4817_/A vssd1 vssd1 vccd1 vccd1 _4674_/Y sky130_fd_sc_hd__nand2_1
X_3625_ _3625_/A _3625_/B vssd1 vssd1 vccd1 vccd1 _3625_/Y sky130_fd_sc_hd__nand2_1
X_3556_ _3519_/B _3567_/B _3386_/X vssd1 vssd1 vccd1 vccd1 _3562_/A sky130_fd_sc_hd__o21ba_1
XFILLER_88_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2507_ hold44/X vssd1 vssd1 vccd1 vccd1 _2821_/A sky130_fd_sc_hd__inv_2
X_3487_ _3610_/B _3487_/B vssd1 vssd1 vccd1 vccd1 _3614_/B sky130_fd_sc_hd__nand2_1
X_5226_ _5228_/CLK _5226_/D vssd1 vssd1 vccd1 vccd1 _5226_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5157_ _5251_/CLK _5157_/D vssd1 vssd1 vccd1 vccd1 _5157_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5088_ _5124_/CLK _5088_/D vssd1 vssd1 vccd1 vccd1 _5088_/Q sky130_fd_sc_hd__dfxtp_1
X_4108_ _4169_/B _5111_/Q _4095_/X _5112_/Q vssd1 vssd1 vccd1 vccd1 _4110_/A sky130_fd_sc_hd__a31oi_1
X_4039_ _4039_/A _4039_/B vssd1 vssd1 vccd1 vccd1 _4040_/B sky130_fd_sc_hd__and2_1
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3410_ _5138_/Q _3845_/B vssd1 vssd1 vccd1 vccd1 _3472_/A sky130_fd_sc_hd__nor2_1
X_4390_ _4390_/A _4390_/B vssd1 vssd1 vccd1 vccd1 _4390_/Y sky130_fd_sc_hd__nand2_1
X_3341_ _3341_/A _3341_/B _3345_/A vssd1 vssd1 vccd1 vccd1 _3341_/X sky130_fd_sc_hd__and3_1
XFILLER_85_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3272_ _3271_/B _3271_/A _2969_/X vssd1 vssd1 vccd1 vccd1 _3272_/X sky130_fd_sc_hd__a21o_1
XFILLER_87_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5011_ _5120_/CLK hold25/X vssd1 vssd1 vccd1 vccd1 _5011_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2987_ _3276_/A _3775_/B vssd1 vssd1 vccd1 vccd1 _2987_/Y sky130_fd_sc_hd__nand2_1
X_4726_ _4741_/A vssd1 vssd1 vccd1 vccd1 _4735_/C sky130_fd_sc_hd__inv_2
X_4657_ _4657_/A _4657_/B vssd1 vssd1 vccd1 vccd1 _4658_/A sky130_fd_sc_hd__nand2_1
X_3608_ _3608_/A _3608_/B vssd1 vssd1 vccd1 vccd1 _3611_/A sky130_fd_sc_hd__nor2_1
X_4588_ _4588_/A _4588_/B vssd1 vssd1 vccd1 vccd1 _4588_/Y sky130_fd_sc_hd__nor2_2
XFILLER_1_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3539_ _3539_/A _3539_/B vssd1 vssd1 vccd1 vccd1 _3540_/C sky130_fd_sc_hd__nor2_1
XFILLER_67_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5209_ _5228_/CLK _5209_/D vssd1 vssd1 vccd1 vccd1 _5209_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2910_ _2910_/A vssd1 vssd1 vccd1 vccd1 _2910_/Y sky130_fd_sc_hd__inv_2
X_3890_ _5124_/Q vssd1 vssd1 vccd1 vccd1 _4962_/A sky130_fd_sc_hd__inv_2
X_2841_ _3863_/A vssd1 vssd1 vccd1 vccd1 _2841_/X sky130_fd_sc_hd__buf_2
XFILLER_31_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2772_ _2772_/A _2772_/B vssd1 vssd1 vccd1 vccd1 _2875_/A sky130_fd_sc_hd__nor2_2
XPHY_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4511_ _4506_/A _4510_/Y _4204_/X vssd1 vssd1 vccd1 vccd1 _4511_/X sky130_fd_sc_hd__a21o_1
X_4442_ _4434_/X _4437_/X _4439_/X _2915_/X _4441_/Y vssd1 vssd1 vccd1 vccd1 _5078_/D
+ sky130_fd_sc_hd__o311a_1
X_4373_ _5108_/Q _5076_/Q vssd1 vssd1 vccd1 vccd1 _4394_/A sky130_fd_sc_hd__nor2_1
X_3324_ _3324_/A _3324_/B vssd1 vssd1 vccd1 vccd1 _3325_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3255_ _3254_/X _3238_/Y _2963_/X vssd1 vssd1 vccd1 vccd1 _3255_/X sky130_fd_sc_hd__a21o_1
XFILLER_66_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3186_ _5285_/Q vssd1 vssd1 vccd1 vccd1 _3707_/B sky130_fd_sc_hd__inv_2
XFILLER_81_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4709_ _4709_/A vssd1 vssd1 vccd1 vccd1 _4720_/B sky130_fd_sc_hd__inv_2
XFILLER_78_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_67_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3040_ _5185_/Q _3719_/B vssd1 vssd1 vccd1 vccd1 _3042_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4991_ _4992_/CLK hold5/X vssd1 vssd1 vccd1 vccd1 _4992_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3942_ _5121_/Q _3923_/Y _3925_/X _3933_/X _3941_/Y vssd1 vssd1 vccd1 vccd1 _4979_/S
+ sky130_fd_sc_hd__o2111a_4
X_3873_ _3873_/A _3873_/B vssd1 vssd1 vccd1 vccd1 _3873_/Y sky130_fd_sc_hd__nand2_1
X_2824_ _2795_/Y _2819_/Y _2823_/Y vssd1 vssd1 vccd1 vccd1 _5285_/D sky130_fd_sc_hd__a21oi_1
X_2755_ _2882_/B _2755_/B vssd1 vssd1 vccd1 vccd1 _2902_/C sky130_fd_sc_hd__nand2_1
X_2686_ _5290_/Q _4628_/A vssd1 vssd1 vccd1 vccd1 _2993_/B sky130_fd_sc_hd__or2_2
X_4425_ _4425_/A _4912_/B vssd1 vssd1 vccd1 vccd1 _4425_/Y sky130_fd_sc_hd__nand2_1
X_4356_ _4356_/A _4685_/B vssd1 vssd1 vccd1 vccd1 _4357_/B sky130_fd_sc_hd__nand2_1
XFILLER_58_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3307_ _3300_/A _3305_/Y _3306_/X vssd1 vssd1 vccd1 vccd1 _3307_/X sky130_fd_sc_hd__a21o_1
X_4287_ _4301_/B _4302_/A vssd1 vssd1 vccd1 vccd1 _4556_/A sky130_fd_sc_hd__nor2_4
X_3238_ _3254_/B _3254_/A vssd1 vssd1 vccd1 vccd1 _3238_/Y sky130_fd_sc_hd__nand2_2
XFILLER_39_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3169_ _3150_/A _3168_/Y _3150_/B vssd1 vssd1 vccd1 vccd1 _3170_/A sky130_fd_sc_hd__o21ba_1
XFILLER_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_89_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2540_ _5043_/Q vssd1 vssd1 vccd1 vccd1 _4699_/A sky130_fd_sc_hd__inv_2
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4210_ _4770_/A vssd1 vssd1 vccd1 vccd1 _4778_/A sky130_fd_sc_hd__buf_2
X_5190_ _5195_/CLK _5190_/D vssd1 vssd1 vccd1 vccd1 _5190_/Q sky130_fd_sc_hd__dfxtp_1
X_4141_ _5105_/Q vssd1 vssd1 vccd1 vccd1 _4252_/A sky130_fd_sc_hd__inv_2
X_4072_ _4208_/D _4222_/A _4208_/B _4207_/A vssd1 vssd1 vccd1 vccd1 _4180_/A sky130_fd_sc_hd__a31o_4
XFILLER_36_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3023_ _3705_/A _3023_/B vssd1 vssd1 vccd1 vccd1 _3023_/Y sky130_fd_sc_hd__nand2_1
XFILLER_24_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4974_ _4951_/X _4951_/B _4979_/S vssd1 vssd1 vccd1 vccd1 _4974_/X sky130_fd_sc_hd__mux2_1
X_3925_ _5117_/Q _3924_/Y _4930_/B _5006_/Q vssd1 vssd1 vccd1 vccd1 _3925_/X sky130_fd_sc_hd__o22a_1
X_3856_ _5134_/Q _3849_/X _3844_/X _3855_/Y vssd1 vssd1 vccd1 vccd1 _5134_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3787_ _3794_/A _3787_/B vssd1 vssd1 vccd1 vccd1 _3787_/Y sky130_fd_sc_hd__nand2_1
X_2807_ _2797_/Y _2806_/Y _2733_/Y vssd1 vssd1 vccd1 vccd1 _2933_/A sky130_fd_sc_hd__o21bai_2
X_2738_ _5300_/Q vssd1 vssd1 vccd1 vccd1 _2739_/A sky130_fd_sc_hd__inv_2
X_4408_ _5114_/Q _5082_/Q vssd1 vssd1 vccd1 vccd1 _4411_/C sky130_fd_sc_hd__xnor2_1
X_2669_ _5303_/Q _4682_/A vssd1 vssd1 vccd1 vccd1 _2747_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4339_ _4504_/B _4504_/A _4510_/B vssd1 vssd1 vccd1 vccd1 _4339_/X sky130_fd_sc_hd__or3_4
XFILLER_59_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3710_ _3762_/A vssd1 vssd1 vccd1 vccd1 _3710_/X sky130_fd_sc_hd__buf_2
X_4690_ _4801_/B _4684_/A _4801_/A vssd1 vssd1 vccd1 vccd1 _4690_/Y sky130_fd_sc_hd__o21bai_1
X_3641_ _3641_/A _3641_/B vssd1 vssd1 vccd1 vccd1 _3641_/Y sky130_fd_sc_hd__nor2_1
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3572_ _3572_/A _3572_/B _3572_/C vssd1 vssd1 vccd1 vccd1 _3572_/X sky130_fd_sc_hd__and3_1
X_2523_ _5047_/Q vssd1 vssd1 vccd1 vccd1 _4592_/A sky130_fd_sc_hd__inv_2
X_5311_ _5311_/CLK _5311_/D vssd1 vssd1 vccd1 vccd1 _5311_/Q sky130_fd_sc_hd__dfxtp_1
X_5242_ _5251_/CLK _5242_/D vssd1 vssd1 vccd1 vccd1 _5242_/Q sky130_fd_sc_hd__dfxtp_1
X_5173_ _5179_/CLK _5173_/D vssd1 vssd1 vccd1 vccd1 _5173_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4124_ _4111_/X _4112_/X _4094_/X _4118_/A _5109_/Q vssd1 vssd1 vccd1 vccd1 _4125_/B
+ sky130_fd_sc_hd__a41oi_1
Xinput1 enable_in vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_1
XFILLER_56_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4055_ _4055_/A _4055_/B vssd1 vssd1 vccd1 vccd1 _4056_/A sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_48_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5112_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_83_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3006_ _4633_/A _5288_/Q vssd1 vssd1 vccd1 vccd1 _3007_/A sky130_fd_sc_hd__nand2_1
XPHY_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4957_ _4961_/B vssd1 vssd1 vccd1 vccd1 _4962_/B sky130_fd_sc_hd__inv_2
X_3908_ _5119_/Q vssd1 vssd1 vccd1 vccd1 _4940_/A sky130_fd_sc_hd__inv_2
X_4888_ _5016_/Q vssd1 vssd1 vccd1 vccd1 _4898_/B sky130_fd_sc_hd__inv_2
X_3839_ _3847_/A _3839_/B vssd1 vssd1 vccd1 vccd1 _3839_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_39_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5277_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4811_ _4673_/A _4817_/B _4611_/Y vssd1 vssd1 vccd1 vccd1 _4813_/A sky130_fd_sc_hd__o21a_1
X_4742_ _4742_/A _4742_/B vssd1 vssd1 vccd1 vccd1 _4742_/Y sky130_fd_sc_hd__nand2_1
XFILLER_33_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4673_ _4673_/A _4673_/B vssd1 vssd1 vccd1 vccd1 _4817_/A sky130_fd_sc_hd__nor2_1
X_3624_ _5205_/Q _3596_/X _3621_/X _3623_/Y _3591_/X vssd1 vssd1 vccd1 vccd1 _5205_/D
+ sky130_fd_sc_hd__o221a_1
X_3555_ _3572_/A _3572_/C vssd1 vssd1 vccd1 vccd1 _3567_/B sky130_fd_sc_hd__and2_1
X_3486_ _3833_/B _5142_/Q vssd1 vssd1 vccd1 vccd1 _3487_/B sky130_fd_sc_hd__nand2_1
X_2506_ _3011_/A vssd1 vssd1 vccd1 vccd1 _2506_/X sky130_fd_sc_hd__buf_2
XFILLER_88_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5225_ _5280_/CLK _5225_/D vssd1 vssd1 vccd1 vccd1 _5225_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5156_ _5250_/CLK _5156_/D vssd1 vssd1 vccd1 vccd1 _5156_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5087_ _5118_/CLK _5087_/D vssd1 vssd1 vccd1 vccd1 _5087_/Q sky130_fd_sc_hd__dfxtp_1
X_4107_ _4126_/A vssd1 vssd1 vccd1 vccd1 _4169_/B sky130_fd_sc_hd__clkbuf_2
X_4038_ _4038_/A vssd1 vssd1 vccd1 vccd1 _4040_/A sky130_fd_sc_hd__inv_2
XFILLER_71_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3340_ _5227_/Q _3321_/X _3336_/X _3339_/Y _3316_/X vssd1 vssd1 vccd1 vccd1 _5227_/D
+ sky130_fd_sc_hd__o221a_1
X_5010_ _5118_/CLK hold18/X vssd1 vssd1 vccd1 vccd1 _5010_/Q sky130_fd_sc_hd__dfxtp_1
X_3271_ _3271_/A _3271_/B vssd1 vssd1 vccd1 vccd1 _3271_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_66_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2986_ _5260_/Q vssd1 vssd1 vccd1 vccd1 _3775_/B sky130_fd_sc_hd__inv_2
X_4725_ _4725_/A _4725_/B vssd1 vssd1 vccd1 vccd1 _4741_/A sky130_fd_sc_hd__nor2_2
X_4656_ _4653_/A _4650_/B _4653_/B vssd1 vssd1 vccd1 vccd1 _4830_/B sky130_fd_sc_hd__o21ba_1
X_4587_ _4912_/B _4587_/B vssd1 vssd1 vccd1 vccd1 _4587_/Y sky130_fd_sc_hd__nand2_1
X_3607_ _3614_/B _3614_/A vssd1 vssd1 vccd1 vccd1 _3610_/A sky130_fd_sc_hd__or2_1
X_3538_ _3521_/Y _3524_/Y _3544_/B vssd1 vssd1 vccd1 vccd1 _3540_/B sky130_fd_sc_hd__a21o_1
X_3469_ _3465_/B _3640_/B _3465_/A vssd1 vssd1 vccd1 vccd1 _3629_/B sky130_fd_sc_hd__o21ba_1
X_5208_ _5228_/CLK _5208_/D vssd1 vssd1 vccd1 vccd1 _5208_/Q sky130_fd_sc_hd__dfxtp_1
X_5139_ _5204_/CLK _5139_/D vssd1 vssd1 vccd1 vccd1 _5139_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2840_ _2634_/X _2835_/Y _2836_/X _2837_/X _2839_/Y vssd1 vssd1 vccd1 vccd1 _5283_/D
+ sky130_fd_sc_hd__o311a_1
XPHY_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2771_ _2760_/A _2885_/B _2767_/Y _2770_/Y vssd1 vssd1 vccd1 vccd1 _2853_/B sky130_fd_sc_hd__o211a_1
XPHY_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4510_ _4510_/A _4510_/B vssd1 vssd1 vccd1 vccd1 _4510_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4441_ _4528_/A _4713_/B vssd1 vssd1 vccd1 vccd1 _4441_/Y sky130_fd_sc_hd__nand2_1
X_4372_ _4372_/A _4449_/B vssd1 vssd1 vccd1 vccd1 _4378_/A sky130_fd_sc_hd__nand2_1
X_3323_ _3775_/B _5164_/Q _3330_/A vssd1 vssd1 vccd1 vccd1 _3324_/A sky130_fd_sc_hd__a21o_1
X_3254_ _3254_/A _3254_/B vssd1 vssd1 vccd1 vccd1 _3254_/X sky130_fd_sc_hd__or2_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3185_ _3197_/B _3197_/A _3204_/A _3184_/Y vssd1 vssd1 vccd1 vccd1 _3199_/B sky130_fd_sc_hd__o22ai_4
XFILLER_81_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2969_ _3361_/A vssd1 vssd1 vccd1 vccd1 _2969_/X sky130_fd_sc_hd__buf_2
X_4708_ _4710_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4709_/A sky130_fd_sc_hd__nor2_1
X_4639_ _5021_/Q _5053_/Q vssd1 vssd1 vccd1 vccd1 _4878_/B sky130_fd_sc_hd__nand2_2
XFILLER_89_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4990_ _4990_/CLK _4990_/D vssd1 vssd1 vccd1 vccd1 _4990_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_90_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3941_ _3898_/B _5012_/Q _3934_/Y _3936_/X _3940_/X vssd1 vssd1 vccd1 vccd1 _3941_/Y
+ sky130_fd_sc_hd__a2111oi_2
XFILLER_90_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3872_ _5128_/Q _3862_/X _3870_/X _3871_/Y vssd1 vssd1 vccd1 vccd1 _5128_/D sky130_fd_sc_hd__o211a_1
X_2823_ _5285_/Q _3199_/C _4238_/B vssd1 vssd1 vccd1 vccd1 _2823_/Y sky130_fd_sc_hd__o21ai_1
X_2754_ _4788_/A _5306_/Q vssd1 vssd1 vccd1 vccd1 _2755_/B sky130_fd_sc_hd__nand2_1
XFILLER_8_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2685_ _2954_/B vssd1 vssd1 vccd1 vccd1 _2685_/Y sky130_fd_sc_hd__inv_2
X_4424_ _4770_/A vssd1 vssd1 vccd1 vccd1 _4912_/B sky130_fd_sc_hd__clkbuf_4
X_4355_ _4355_/A vssd1 vssd1 vccd1 vccd1 _4496_/B sky130_fd_sc_hd__inv_2
X_3306_ _3615_/A vssd1 vssd1 vccd1 vccd1 _3306_/X sky130_fd_sc_hd__buf_2
X_4286_ _4286_/A _4626_/B vssd1 vssd1 vccd1 vccd1 _4302_/A sky130_fd_sc_hd__nor2_2
X_3237_ _3237_/A vssd1 vssd1 vccd1 vccd1 _3254_/A sky130_fd_sc_hd__inv_2
XFILLER_27_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3168_ _5178_/Q _3737_/B vssd1 vssd1 vccd1 vccd1 _3168_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3099_ _3324_/B _3099_/B vssd1 vssd1 vccd1 vccd1 _3330_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4140_ _4250_/A _4144_/B _4139_/Y vssd1 vssd1 vccd1 vccd1 _5106_/D sky130_fd_sc_hd__a21oi_1
X_4071_ _4070_/A _4070_/C _4558_/A vssd1 vssd1 vccd1 vccd1 _4207_/A sky130_fd_sc_hd__a21oi_4
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3022_ _5286_/Q _3022_/B vssd1 vssd1 vccd1 vccd1 _3022_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4973_ _4955_/X _4954_/X _4979_/S vssd1 vssd1 vccd1 vccd1 _4973_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3924_ _5007_/Q vssd1 vssd1 vccd1 vccd1 _3924_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3855_ _3860_/A _3855_/B vssd1 vssd1 vccd1 vccd1 _3855_/Y sky130_fd_sc_hd__nand2_1
X_2806_ _2954_/A _2954_/B _2724_/Y vssd1 vssd1 vccd1 vccd1 _2806_/Y sky130_fd_sc_hd__a21oi_1
X_3786_ _5161_/Q _3783_/X _3778_/X _3785_/Y vssd1 vssd1 vccd1 vccd1 _5161_/D sky130_fd_sc_hd__o211a_1
X_2737_ _2735_/Y _2737_/B vssd1 vssd1 vccd1 vccd1 _2937_/A sky130_fd_sc_hd__and2b_1
X_2668_ _2914_/B _2914_/C _2911_/B vssd1 vssd1 vccd1 vccd1 _2674_/A sky130_fd_sc_hd__and3_1
X_4407_ _4416_/A _4403_/Y _4416_/B vssd1 vssd1 vccd1 vccd1 _4407_/Y sky130_fd_sc_hd__a21oi_1
X_2599_ _5295_/Q _2586_/X _2582_/X _2598_/Y vssd1 vssd1 vccd1 vccd1 _5295_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4338_ _4506_/B _4338_/B vssd1 vssd1 vccd1 vccd1 _4510_/B sky130_fd_sc_hd__nand2_1
XFILLER_59_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4269_ _5065_/Q vssd1 vssd1 vccd1 vccd1 _4610_/B sky130_fd_sc_hd__inv_2
XFILLER_86_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3640_ _3640_/A _3640_/B vssd1 vssd1 vccd1 vccd1 _3641_/B sky130_fd_sc_hd__nand2_1
X_3571_ _5215_/Q _3365_/X _3569_/Y _3570_/X _3363_/X vssd1 vssd1 vccd1 vccd1 _5215_/D
+ sky130_fd_sc_hd__o221a_1
X_2522_ _4550_/A vssd1 vssd1 vccd1 vccd1 _2522_/X sky130_fd_sc_hd__clkbuf_2
X_5310_ _5311_/CLK _5310_/D vssd1 vssd1 vccd1 vccd1 _5310_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5241_ _5274_/CLK _5241_/D vssd1 vssd1 vccd1 vccd1 _5241_/Q sky130_fd_sc_hd__dfxtp_1
X_5172_ _5179_/CLK _5172_/D vssd1 vssd1 vccd1 vccd1 _5172_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4123_ _4589_/A vssd1 vssd1 vccd1 vccd1 _4734_/A sky130_fd_sc_hd__buf_2
Xinput2 oversample_in[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__clkbuf_1
X_4054_ _4054_/A vssd1 vssd1 vccd1 vccd1 _4057_/A sky130_fd_sc_hd__inv_2
X_3005_ _5257_/Q _2977_/X _3003_/Y _3004_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _5257_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4956_ _4958_/B _4958_/A vssd1 vssd1 vccd1 vccd1 _4961_/B sky130_fd_sc_hd__nor2_1
X_3907_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3907_/X sky130_fd_sc_hd__clkbuf_2
X_4887_ _5017_/Q vssd1 vssd1 vccd1 vccd1 _4892_/A sky130_fd_sc_hd__inv_2
XFILLER_20_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3838_ _5141_/Q _3835_/X _3830_/X _3837_/Y vssd1 vssd1 vccd1 vccd1 _5141_/D sky130_fd_sc_hd__o211a_1
XFILLER_3_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3769_ _3769_/A vssd1 vssd1 vccd1 vccd1 _3823_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_3_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4810_ _4810_/A _4810_/B vssd1 vssd1 vccd1 vccd1 _4817_/B sky130_fd_sc_hd__and2_1
XFILLER_21_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4741_ _4741_/A _4741_/B _4744_/B _4741_/D vssd1 vssd1 vccd1 vccd1 _4742_/A sky130_fd_sc_hd__or4_4
X_4672_ _5033_/Q _5065_/Q vssd1 vssd1 vccd1 vccd1 _4673_/A sky130_fd_sc_hd__nor2_1
X_3623_ _3623_/A _3623_/B vssd1 vssd1 vccd1 vccd1 _3623_/Y sky130_fd_sc_hd__nor2_1
X_3554_ _5218_/Q _3365_/X _3552_/Y _3553_/X _3363_/X vssd1 vssd1 vccd1 vccd1 _5218_/D
+ sky130_fd_sc_hd__o221a_1
X_3485_ _3485_/A vssd1 vssd1 vccd1 vccd1 _3610_/B sky130_fd_sc_hd__inv_2
X_2505_ _2888_/A vssd1 vssd1 vccd1 vccd1 _3011_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_88_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5224_ _5280_/CLK _5224_/D vssd1 vssd1 vccd1 vccd1 _5224_/Q sky130_fd_sc_hd__dfxtp_2
X_5155_ _5250_/CLK _5155_/D vssd1 vssd1 vccd1 vccd1 _5155_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5086_ _5125_/CLK _5086_/D vssd1 vssd1 vccd1 vccd1 _5086_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4106_ _4106_/A _4106_/B _4201_/C vssd1 vssd1 vccd1 vccd1 _4126_/A sky130_fd_sc_hd__nor3_4
X_4037_ _4037_/A _4037_/B _4037_/C vssd1 vssd1 vccd1 vccd1 _4045_/C sky130_fd_sc_hd__nand3_4
XFILLER_56_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4939_ _5119_/Q _4939_/B vssd1 vssd1 vccd1 vccd1 _4941_/A sky130_fd_sc_hd__nor2_1
XFILLER_24_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3270_ _3142_/B _3274_/B _3142_/A vssd1 vssd1 vccd1 vccd1 _3271_/B sky130_fd_sc_hd__o21ba_1
XFILLER_87_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2985_ _2984_/Y _2799_/A _2979_/B vssd1 vssd1 vccd1 vccd1 _2985_/Y sky130_fd_sc_hd__a21oi_2
X_4724_ _4739_/A _4739_/B _4744_/B _4741_/D vssd1 vssd1 vccd1 vccd1 _4735_/A sky130_fd_sc_hd__o22ai_1
XFILLER_21_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4655_ _4840_/A _4840_/B _4654_/Y vssd1 vssd1 vccd1 vccd1 _4830_/A sky130_fd_sc_hd__o21ai_1
X_4586_ _5051_/Q vssd1 vssd1 vccd1 vccd1 _4588_/B sky130_fd_sc_hd__inv_2
X_3606_ _3604_/X _3605_/Y _3202_/X vssd1 vssd1 vccd1 vccd1 _5208_/D sky130_fd_sc_hd__a21oi_1
X_3537_ _5251_/Q _3537_/B vssd1 vssd1 vccd1 vccd1 _3544_/B sky130_fd_sc_hd__nor2_1
XFILLER_67_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3468_ _3638_/A _3638_/B _3467_/X vssd1 vssd1 vccd1 vccd1 _3629_/A sky130_fd_sc_hd__o21bai_1
X_3399_ _3828_/B _5144_/Q vssd1 vssd1 vccd1 vccd1 _3400_/B sky130_fd_sc_hd__nand2_1
X_5207_ _5228_/CLK _5207_/D vssd1 vssd1 vccd1 vccd1 _5207_/Q sky130_fd_sc_hd__dfxtp_1
X_5138_ _5204_/CLK _5138_/D vssd1 vssd1 vccd1 vccd1 _5138_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5069_ _5098_/CLK _5069_/D vssd1 vssd1 vccd1 vccd1 _5069_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_25_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2770_ _2770_/A vssd1 vssd1 vccd1 vccd1 _2770_/Y sky130_fd_sc_hd__inv_2
XPHY_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4440_ _4440_/A vssd1 vssd1 vccd1 vccd1 _4528_/A sky130_fd_sc_hd__buf_2
X_4371_ _5107_/Q _5075_/Q vssd1 vssd1 vccd1 vccd1 _4449_/B sky130_fd_sc_hd__nand2_1
X_3322_ _3079_/Y _3333_/A _3096_/Y vssd1 vssd1 vccd1 vccd1 _3330_/A sky130_fd_sc_hd__o21ai_1
XFILLER_85_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3253_ _3613_/A vssd1 vssd1 vccd1 vccd1 _3253_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_85_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3184_ _3713_/B _5187_/Q _3180_/Y _3183_/Y vssd1 vssd1 vccd1 vccd1 _3184_/Y sky130_fd_sc_hd__a22oi_4
XFILLER_66_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2968_ _2968_/A _2968_/B vssd1 vssd1 vccd1 vccd1 _2968_/Y sky130_fd_sc_hd__nor2_1
X_4707_ _4761_/A _4763_/A vssd1 vssd1 vccd1 vccd1 _4717_/A sky130_fd_sc_hd__nor2_2
X_4638_ _5022_/Q _5054_/Q vssd1 vssd1 vccd1 vccd1 _4871_/B sky130_fd_sc_hd__nand2_1
X_2899_ _3262_/A vssd1 vssd1 vccd1 vccd1 _2899_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_89_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4569_ _4569_/A vssd1 vssd1 vccd1 vccd1 _4571_/A sky130_fd_sc_hd__inv_2
XFILLER_1_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_75_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3940_ _5124_/Q _3937_/Y _5119_/Q _3938_/Y _3939_/X vssd1 vssd1 vccd1 vccd1 _3940_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_90_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3871_ _3873_/A _3871_/B vssd1 vssd1 vccd1 vccd1 _3871_/Y sky130_fd_sc_hd__nand2_1
XFILLER_16_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2822_ _4132_/A vssd1 vssd1 vccd1 vccd1 _4238_/B sky130_fd_sc_hd__buf_4
XFILLER_31_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2753_ _2753_/A vssd1 vssd1 vccd1 vccd1 _2882_/B sky130_fd_sc_hd__inv_2
X_2684_ _2714_/B _2712_/A _2683_/Y vssd1 vssd1 vccd1 vccd1 _2954_/B sky130_fd_sc_hd__o21a_1
XFILLER_8_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4423_ _4423_/A _4423_/B _4429_/B _4423_/D vssd1 vssd1 vccd1 vccd1 _4425_/A sky130_fd_sc_hd__or4_4
X_4354_ _4354_/A _4685_/B vssd1 vssd1 vccd1 vccd1 _4355_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3305_ _3305_/A _3305_/B vssd1 vssd1 vccd1 vccd1 _3305_/Y sky130_fd_sc_hd__nand2_1
X_4285_ _5056_/Q vssd1 vssd1 vccd1 vccd1 _4626_/B sky130_fd_sc_hd__inv_2
X_3236_ _3236_/A _3236_/B vssd1 vssd1 vccd1 vccd1 _3254_/B sky130_fd_sc_hd__or2_1
XFILLER_39_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3167_ _3167_/A _3241_/A vssd1 vssd1 vccd1 vccd1 _3167_/Y sky130_fd_sc_hd__nor2_1
X_3098_ _3775_/B _5164_/Q vssd1 vssd1 vccd1 vccd1 _3099_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4070_ _4070_/A _4558_/A _4070_/C vssd1 vssd1 vccd1 vccd1 _4208_/B sky130_fd_sc_hd__nand3_4
X_3021_ _3015_/Y _3020_/Y _2869_/X vssd1 vssd1 vccd1 vccd1 _5255_/D sky130_fd_sc_hd__o21a_1
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4972_ _4960_/X _4959_/X _4979_/S vssd1 vssd1 vccd1 vccd1 _4972_/X sky130_fd_sc_hd__mux2_1
XFILLER_63_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3923_ _5011_/Q vssd1 vssd1 vccd1 vccd1 _3923_/Y sky130_fd_sc_hd__inv_2
X_3854_ _5135_/Q _3849_/X _3844_/X _3853_/Y vssd1 vssd1 vccd1 vccd1 _5135_/D sky130_fd_sc_hd__o211a_1
X_2805_ _2966_/A _2966_/B _2805_/C vssd1 vssd1 vccd1 vccd1 _2954_/A sky130_fd_sc_hd__nand3_2
X_3785_ _3794_/A _3785_/B vssd1 vssd1 vccd1 vccd1 _3785_/Y sky130_fd_sc_hd__nand2_1
X_2736_ _4815_/A _5301_/Q vssd1 vssd1 vccd1 vccd1 _2737_/B sky130_fd_sc_hd__nand2_1
X_2667_ _4691_/A _5304_/Q vssd1 vssd1 vccd1 vccd1 _2911_/B sky130_fd_sc_hd__nand2_1
X_4406_ _4406_/A _4406_/B vssd1 vssd1 vccd1 vccd1 _4416_/B sky130_fd_sc_hd__nor2_1
X_2598_ _2602_/A _4652_/A vssd1 vssd1 vccd1 vccd1 _2598_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_86_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4337_ _4337_/A _4610_/B vssd1 vssd1 vccd1 vccd1 _4338_/B sky130_fd_sc_hd__nand2_1
XFILLER_75_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4268_ _5098_/Q _5066_/Q vssd1 vssd1 vccd1 vccd1 _4504_/A sky130_fd_sc_hd__nor2_2
XFILLER_74_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3219_ _3223_/B _3223_/C _3223_/A vssd1 vssd1 vccd1 vccd1 _3224_/C sky130_fd_sc_hd__o21ai_2
XFILLER_46_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4199_ _4199_/A vssd1 vssd1 vccd1 vccd1 _4542_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_27_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3570_ _3569_/B _3569_/A _3361_/X vssd1 vssd1 vccd1 vccd1 _3570_/X sky130_fd_sc_hd__a21o_1
X_2521_ _3315_/A vssd1 vssd1 vccd1 vccd1 _4550_/A sky130_fd_sc_hd__buf_1
XFILLER_5_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5240_ _5280_/CLK _5240_/D vssd1 vssd1 vccd1 vccd1 _5240_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5171_ _5171_/CLK _5171_/D vssd1 vssd1 vccd1 vccd1 _5171_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4122_ _5110_/Q _4125_/C _4121_/Y vssd1 vssd1 vccd1 vccd1 _5110_/D sky130_fd_sc_hd__o21a_1
XFILLER_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4053_ _4070_/A _5085_/Q _4053_/C vssd1 vssd1 vccd1 vccd1 _4222_/B sky130_fd_sc_hd__nand3_4
XFILLER_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 oversample_in[1] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_1
X_3004_ _3003_/B _3003_/A _2969_/X vssd1 vssd1 vccd1 vccd1 _3004_/X sky130_fd_sc_hd__a21o_1
XFILLER_24_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4955_ _4966_/B _4958_/A _4955_/C vssd1 vssd1 vccd1 vccd1 _4955_/X sky130_fd_sc_hd__and3_1
X_3906_ _3887_/X _4975_/X _3893_/X _3905_/Y vssd1 vssd1 vccd1 vccd1 _5120_/D sky130_fd_sc_hd__o211a_1
X_4886_ _4980_/X vssd1 vssd1 vccd1 vccd1 _4898_/A sky130_fd_sc_hd__inv_2
XFILLER_32_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3837_ _3847_/A _3837_/B vssd1 vssd1 vccd1 vccd1 _3837_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3768_ _3822_/A vssd1 vssd1 vccd1 vccd1 _3768_/X sky130_fd_sc_hd__clkbuf_2
X_2719_ _2957_/B _2719_/B vssd1 vssd1 vccd1 vccd1 _2720_/A sky130_fd_sc_hd__nand2_1
X_3699_ _3873_/B _5127_/Q vssd1 vssd1 vccd1 vccd1 _3700_/A sky130_fd_sc_hd__nand2_1
XFILLER_15_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4740_ _4741_/A _4741_/B _4744_/B _4741_/D vssd1 vssd1 vccd1 vccd1 _4740_/X sky130_fd_sc_hd__o22a_1
X_4671_ _4671_/A _4671_/B vssd1 vssd1 vccd1 vccd1 _4813_/B sky130_fd_sc_hd__nor2_1
X_3622_ _3622_/A _3622_/B vssd1 vssd1 vccd1 vccd1 _3623_/B sky130_fd_sc_hd__and2_1
X_3553_ _3552_/B _3552_/A _3361_/X vssd1 vssd1 vccd1 vccd1 _3553_/X sky130_fd_sc_hd__a21o_1
XFILLER_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3484_ _3620_/B _3622_/B _3620_/A vssd1 vssd1 vccd1 vccd1 _3575_/B sky130_fd_sc_hd__o21ba_1
X_2504_ _2632_/A vssd1 vssd1 vccd1 vccd1 _2888_/A sky130_fd_sc_hd__buf_1
X_5223_ _5251_/CLK _5223_/D vssd1 vssd1 vccd1 vccd1 _5223_/Q sky130_fd_sc_hd__dfxtp_2
X_5154_ _5219_/CLK _5154_/D vssd1 vssd1 vccd1 vccd1 _5154_/Q sky130_fd_sc_hd__dfxtp_1
X_4105_ _4105_/A vssd1 vssd1 vccd1 vccd1 _4106_/B sky130_fd_sc_hd__inv_2
X_5085_ _5085_/CLK _5085_/D vssd1 vssd1 vccd1 vccd1 _5085_/Q sky130_fd_sc_hd__dfxtp_2
X_4036_ _4036_/A _4036_/B vssd1 vssd1 vccd1 vccd1 _4037_/B sky130_fd_sc_hd__nand2_1
XFILLER_2_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4938_ _4951_/A _4938_/B vssd1 vssd1 vccd1 vccd1 _4938_/X sky130_fd_sc_hd__and2_1
XFILLER_52_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4869_ _4869_/A vssd1 vssd1 vccd1 vccd1 _4871_/A sky130_fd_sc_hd__inv_2
XFILLER_20_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2984_ _2687_/Y _2989_/A _2798_/A vssd1 vssd1 vccd1 vccd1 _2984_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4723_ _4746_/A _4746_/B _4744_/A vssd1 vssd1 vccd1 vccd1 _4741_/D sky130_fd_sc_hd__a21oi_2
X_4654_ _4845_/A _4842_/A vssd1 vssd1 vccd1 vccd1 _4654_/Y sky130_fd_sc_hd__nor2_1
X_4585_ _4574_/X _4634_/B _4582_/Y _4583_/X _4584_/X vssd1 vssd1 vccd1 vccd1 _5052_/D
+ sky130_fd_sc_hd__o221a_1
X_3605_ _3605_/A _5208_/Q vssd1 vssd1 vccd1 vccd1 _3605_/Y sky130_fd_sc_hd__nand2_1
X_3536_ _5155_/Q vssd1 vssd1 vccd1 vccd1 _3537_/B sky130_fd_sc_hd__inv_2
X_3467_ _3647_/B _3641_/A vssd1 vssd1 vccd1 vccd1 _3467_/X sky130_fd_sc_hd__or2_1
X_5206_ _5228_/CLK _5206_/D vssd1 vssd1 vccd1 vccd1 _5206_/Q sky130_fd_sc_hd__dfxtp_1
X_3398_ _5144_/Q _3828_/B vssd1 vssd1 vccd1 vccd1 _3406_/B sky130_fd_sc_hd__or2_2
X_5137_ _5204_/CLK _5137_/D vssd1 vssd1 vccd1 vccd1 _5137_/Q sky130_fd_sc_hd__dfxtp_1
X_5068_ _5098_/CLK _5068_/D vssd1 vssd1 vccd1 vccd1 _5068_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4019_ _4023_/B _4023_/A _4028_/A _4018_/X vssd1 vssd1 vccd1 vccd1 _4063_/A sky130_fd_sc_hd__o22ai_4
XFILLER_25_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4370_ _4370_/A _4701_/B vssd1 vssd1 vccd1 vccd1 _4372_/A sky130_fd_sc_hd__nand2_1
X_3321_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3321_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_3_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3252_ _5243_/Q _3210_/X _3250_/Y _3251_/X _3208_/X vssd1 vssd1 vccd1 vccd1 _5243_/D
+ sky130_fd_sc_hd__o221a_1
X_3183_ _3212_/A vssd1 vssd1 vccd1 vccd1 _3183_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2967_ _2973_/A _2973_/B _2712_/A vssd1 vssd1 vccd1 vccd1 _2968_/B sky130_fd_sc_hd__o21a_1
X_4706_ _4706_/A vssd1 vssd1 vccd1 vccd1 _4763_/A sky130_fd_sc_hd__inv_2
X_2898_ _2903_/B _2764_/X _2882_/B _2897_/X vssd1 vssd1 vccd1 vccd1 _2898_/X sky130_fd_sc_hd__a31o_1
X_4637_ _4875_/A _4878_/C _4877_/B vssd1 vssd1 vccd1 vccd1 _4868_/A sky130_fd_sc_hd__nand3b_2
X_4568_ _4568_/A _4576_/B vssd1 vssd1 vccd1 vccd1 _4569_/A sky130_fd_sc_hd__nand2_1
XFILLER_1_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3519_ _3562_/B _3519_/B _3390_/Y vssd1 vssd1 vccd1 vccd1 _3519_/X sky130_fd_sc_hd__or3b_4
X_4499_ _4499_/A _4499_/B vssd1 vssd1 vccd1 vccd1 _4499_/Y sky130_fd_sc_hd__nand2_1
XFILLER_89_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_20_clk clkbuf_opt_0_clk/X vssd1 vssd1 vccd1 vccd1 _4990_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_21_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3870_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3870_/X sky130_fd_sc_hd__buf_2
X_2821_ _2821_/A vssd1 vssd1 vccd1 vccd1 _4132_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_11_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5120_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2752_ _5306_/Q _4788_/A vssd1 vssd1 vccd1 vccd1 _2753_/A sky130_fd_sc_hd__nor2_2
X_2683_ _2714_/A vssd1 vssd1 vccd1 vccd1 _2683_/Y sky130_fd_sc_hd__inv_2
X_4422_ _4423_/A _4423_/B _4429_/B _4423_/D vssd1 vssd1 vccd1 vccd1 _4422_/X sky130_fd_sc_hd__o22a_1
X_4353_ _5067_/Q vssd1 vssd1 vccd1 vccd1 _4685_/B sky130_fd_sc_hd__inv_2
X_4284_ _5088_/Q _5056_/Q vssd1 vssd1 vccd1 vccd1 _4301_/B sky130_fd_sc_hd__nor2_2
X_3304_ _3646_/A vssd1 vssd1 vccd1 vccd1 _3304_/X sky130_fd_sc_hd__clkbuf_2
X_3235_ _2901_/X _3232_/Y _2961_/X _3234_/Y vssd1 vssd1 vccd1 vccd1 _5246_/D sky130_fd_sc_hd__o211a_1
XFILLER_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166_ _3236_/A _3236_/B _3165_/Y vssd1 vssd1 vccd1 vccd1 _3231_/A sky130_fd_sc_hd__o21bai_2
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3097_ _5164_/Q _3775_/B vssd1 vssd1 vccd1 vccd1 _3324_/B sky130_fd_sc_hd__or2_1
XFILLER_39_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3999_ _4031_/B _4031_/A vssd1 vssd1 vccd1 vccd1 _4000_/B sky130_fd_sc_hd__nor2_2
XFILLER_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_70_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_0_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5108_/CLK sky130_fd_sc_hd__clkbuf_16
X_3020_ _3023_/B _3018_/X _3019_/Y vssd1 vssd1 vccd1 vccd1 _3020_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_63_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4971_ _4964_/X _4964_/A _4979_/S vssd1 vssd1 vccd1 vccd1 _4971_/X sky130_fd_sc_hd__mux2_1
XFILLER_36_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3922_ _3907_/X _4979_/X _3911_/X _3921_/Y vssd1 vssd1 vccd1 vccd1 _5116_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3853_ _3860_/A _3853_/B vssd1 vssd1 vccd1 vccd1 _3853_/Y sky130_fd_sc_hd__nand2_1
X_2804_ _2804_/A vssd1 vssd1 vccd1 vccd1 _2805_/C sky130_fd_sc_hd__inv_2
X_3784_ _3823_/A vssd1 vssd1 vccd1 vccd1 _3794_/A sky130_fd_sc_hd__clkbuf_2
X_2735_ _5301_/Q _4815_/A vssd1 vssd1 vccd1 vccd1 _2735_/Y sky130_fd_sc_hd__nor2_1
X_2666_ _2675_/A _2666_/B vssd1 vssd1 vccd1 vccd1 _2914_/B sky130_fd_sc_hd__nor2_1
X_4405_ _5081_/Q _4405_/B vssd1 vssd1 vccd1 vccd1 _4406_/B sky130_fd_sc_hd__nor2_1
X_2597_ _5028_/Q vssd1 vssd1 vccd1 vccd1 _4652_/A sky130_fd_sc_hd__inv_2
XFILLER_5_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4336_ _4332_/A _4328_/B _4332_/B vssd1 vssd1 vccd1 vccd1 _4502_/B sky130_fd_sc_hd__o21ba_1
X_4267_ _4267_/A vssd1 vssd1 vccd1 vccd1 _4454_/A sky130_fd_sc_hd__inv_2
XFILLER_86_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4198_ _5088_/Q vssd1 vssd1 vccd1 vccd1 _4286_/A sky130_fd_sc_hd__inv_2
X_3218_ _3218_/A _3227_/B vssd1 vssd1 vccd1 vccd1 _3223_/C sky130_fd_sc_hd__nor2_1
XFILLER_67_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3149_ _3734_/B _5179_/Q vssd1 vssd1 vccd1 vccd1 _3150_/B sky130_fd_sc_hd__and2_1
XFILLER_82_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2520_ _2821_/A vssd1 vssd1 vccd1 vccd1 _3315_/A sky130_fd_sc_hd__buf_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_5170_ _5171_/CLK _5170_/D vssd1 vssd1 vccd1 vccd1 _5170_/Q sky130_fd_sc_hd__dfxtp_1
X_4121_ _4169_/B _4095_/X _4910_/A vssd1 vssd1 vccd1 vccd1 _4121_/Y sky130_fd_sc_hd__a21oi_1
X_4052_ _4052_/A _4059_/A _4052_/C vssd1 vssd1 vccd1 vccd1 _4053_/C sky130_fd_sc_hd__nand3_4
XFILLER_83_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput4 input4/A vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_1
X_3003_ _3003_/A _3003_/B vssd1 vssd1 vccd1 vccd1 _3003_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4954_ _4955_/C _4958_/A vssd1 vssd1 vccd1 vccd1 _4954_/X sky130_fd_sc_hd__and2_1
X_3905_ _3916_/A _3934_/B vssd1 vssd1 vccd1 vccd1 _3905_/Y sky130_fd_sc_hd__nand2_1
X_4885_ _4434_/X _4880_/A _5019_/Q _4588_/Y _2837_/X vssd1 vssd1 vccd1 vccd1 _5019_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3836_ _3863_/A vssd1 vssd1 vccd1 vccd1 _3847_/A sky130_fd_sc_hd__buf_1
X_3767_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3822_/A sky130_fd_sc_hd__clkbuf_2
X_2718_ _4657_/A _5296_/Q vssd1 vssd1 vccd1 vccd1 _2719_/B sky130_fd_sc_hd__nand2_1
X_3698_ _3875_/B _5126_/Q vssd1 vssd1 vccd1 vccd1 _3705_/B sky130_fd_sc_hd__nand2_1
XFILLER_10_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2649_ _2653_/B _2857_/C vssd1 vssd1 vccd1 vccd1 _2661_/B sky130_fd_sc_hd__nor2_1
XFILLER_59_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4319_ _4316_/A _4536_/B _4316_/B vssd1 vssd1 vccd1 vccd1 _4523_/B sky130_fd_sc_hd__o21ba_1
X_5299_ _5301_/CLK _5299_/D vssd1 vssd1 vccd1 vccd1 _5299_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4670_ _4667_/A _4823_/B _4667_/B vssd1 vssd1 vccd1 vccd1 _4810_/B sky130_fd_sc_hd__o21ba_1
X_3621_ _3622_/A _3623_/A _3622_/B _2897_/X vssd1 vssd1 vccd1 vccd1 _3621_/X sky130_fd_sc_hd__a31o_1
X_3552_ _3552_/A _3552_/B vssd1 vssd1 vccd1 vccd1 _3552_/Y sky130_fd_sc_hd__nor2_1
X_2503_ _4199_/A _4911_/B vssd1 vssd1 vccd1 vccd1 _2632_/A sky130_fd_sc_hd__nor2_2
X_3483_ _3618_/A _3618_/B _3482_/X vssd1 vssd1 vccd1 vccd1 _3575_/A sky130_fd_sc_hd__o21bai_1
X_5222_ _5251_/CLK _5222_/D vssd1 vssd1 vccd1 vccd1 _5222_/Q sky130_fd_sc_hd__dfxtp_2
X_5153_ _5219_/CLK _5153_/D vssd1 vssd1 vccd1 vccd1 _5153_/Q sky130_fd_sc_hd__dfxtp_1
X_4104_ _5113_/Q _4101_/Y _4103_/Y vssd1 vssd1 vccd1 vccd1 _5113_/D sky130_fd_sc_hd__o21a_1
XFILLER_29_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5084_ _5085_/CLK _5084_/D vssd1 vssd1 vccd1 vccd1 _5084_/Q sky130_fd_sc_hd__dfxtp_1
X_4035_ _4030_/Y _4045_/B _4032_/Y vssd1 vssd1 vccd1 vccd1 _4037_/A sky130_fd_sc_hd__a21o_1
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4937_ _5118_/Q _4931_/B _4940_/B vssd1 vssd1 vccd1 vccd1 _4938_/B sky130_fd_sc_hd__o21a_1
X_4868_ _4868_/A _4878_/B vssd1 vssd1 vccd1 vccd1 _4869_/A sky130_fd_sc_hd__nand2_1
X_3819_ _5148_/Q _3809_/X _3817_/X _3818_/Y vssd1 vssd1 vccd1 vccd1 _5148_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4799_ _4799_/A _5037_/Q vssd1 vssd1 vccd1 vccd1 _4799_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2983_ _5261_/Q _2977_/X _2981_/Y _2982_/X _2971_/X vssd1 vssd1 vccd1 vccd1 _5261_/D
+ sky130_fd_sc_hd__o221a_1
X_4722_ _5047_/Q _5079_/Q vssd1 vssd1 vccd1 vccd1 _4744_/A sky130_fd_sc_hd__nor2_1
X_4653_ _4653_/A _4653_/B vssd1 vssd1 vccd1 vccd1 _4842_/A sky130_fd_sc_hd__or2_1
X_3604_ _3604_/A _3604_/B _3604_/C vssd1 vssd1 vccd1 vccd1 _3604_/X sky130_fd_sc_hd__or3_1
X_4584_ _4785_/A vssd1 vssd1 vccd1 vccd1 _4584_/X sky130_fd_sc_hd__buf_2
X_3535_ _3530_/Y _3532_/Y _3534_/Y vssd1 vssd1 vccd1 vccd1 _5221_/D sky130_fd_sc_hd__a21oi_1
X_3466_ _3466_/A vssd1 vssd1 vccd1 vccd1 _3641_/A sky130_fd_sc_hd__inv_2
X_5205_ _5285_/CLK _5205_/D vssd1 vssd1 vccd1 vccd1 _5205_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3397_ _3599_/A vssd1 vssd1 vccd1 vccd1 _3489_/A sky130_fd_sc_hd__inv_2
XFILLER_57_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5136_ _5204_/CLK _5136_/D vssd1 vssd1 vccd1 vccd1 _5136_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5067_ _5098_/CLK _5067_/D vssd1 vssd1 vccd1 vccd1 _5067_/Q sky130_fd_sc_hd__dfxtp_1
X_4018_ _4005_/X _4015_/Y _4022_/B _4022_/A vssd1 vssd1 vccd1 vccd1 _4018_/X sky130_fd_sc_hd__o211a_2
XFILLER_25_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3320_ _5230_/Q _3253_/X _3304_/X _3319_/X vssd1 vssd1 vccd1 vccd1 _5230_/D sky130_fd_sc_hd__o211a_1
X_3251_ _3238_/Y _3151_/A _3154_/A _3206_/X vssd1 vssd1 vccd1 vccd1 _3251_/X sky130_fd_sc_hd__a31o_1
XFILLER_78_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3182_ _5186_/Q _3717_/B vssd1 vssd1 vccd1 vccd1 _3212_/A sky130_fd_sc_hd__nor2_2
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2966_ _2966_/A _2966_/B vssd1 vssd1 vccd1 vccd1 _2973_/B sky130_fd_sc_hd__nand2_1
X_2897_ _3642_/A vssd1 vssd1 vccd1 vccd1 _2897_/X sky130_fd_sc_hd__buf_2
X_4705_ _4705_/A _4705_/B vssd1 vssd1 vccd1 vccd1 _4706_/A sky130_fd_sc_hd__nor2_1
X_4636_ _4881_/B _4880_/A vssd1 vssd1 vccd1 vccd1 _4877_/B sky130_fd_sc_hd__nand2_1
X_4567_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4567_/X sky130_fd_sc_hd__buf_2
XFILLER_89_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3518_ _3566_/B _3566_/A _3572_/B vssd1 vssd1 vccd1 vccd1 _3519_/B sky130_fd_sc_hd__or3_1
X_4498_ _4492_/X _5068_/Q _4495_/X _4497_/Y _4432_/X vssd1 vssd1 vccd1 vccd1 _5068_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_89_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3449_ _3858_/B _5133_/Q vssd1 vssd1 vccd1 vccd1 _3450_/B sky130_fd_sc_hd__and2_1
X_5119_ _5120_/CLK _5119_/D vssd1 vssd1 vccd1 vccd1 _5119_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2820_ _3011_/A vssd1 vssd1 vccd1 vccd1 _3199_/C sky130_fd_sc_hd__buf_2
XPHY_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2751_ _2744_/Y _2746_/Y _2750_/X vssd1 vssd1 vccd1 vccd1 _2751_/Y sky130_fd_sc_hd__a21oi_2
X_2682_ _5295_/Q _4652_/A vssd1 vssd1 vccd1 vccd1 _2714_/A sky130_fd_sc_hd__nor2_2
XFILLER_8_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4421_ _5112_/Q _4739_/B vssd1 vssd1 vccd1 vccd1 _4423_/B sky130_fd_sc_hd__nor2_1
X_4352_ _4352_/A _4682_/B vssd1 vssd1 vccd1 vccd1 _4494_/B sky130_fd_sc_hd__nor2_1
X_4283_ _4306_/A _4549_/C _4306_/B vssd1 vssd1 vccd1 vccd1 _4534_/A sky130_fd_sc_hd__o21bai_1
X_3303_ _5233_/Q _3269_/X _3301_/Y _3302_/X _3262_/X vssd1 vssd1 vccd1 vccd1 _5233_/D
+ sky130_fd_sc_hd__o221a_1
X_3234_ _3276_/A _3813_/B vssd1 vssd1 vccd1 vccd1 _3234_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3165_ _3165_/A vssd1 vssd1 vccd1 vccd1 _3165_/Y sky130_fd_sc_hd__inv_2
XFILLER_66_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3096_ _3335_/A vssd1 vssd1 vccd1 vccd1 _3096_/Y sky130_fd_sc_hd__inv_2
XFILLER_54_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3998_ _4032_/A _4000_/A _4031_/A _4031_/B vssd1 vssd1 vccd1 vccd1 _4011_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_22_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2949_ _2949_/A _2949_/B vssd1 vssd1 vccd1 vccd1 _2949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_13_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4619_ _4832_/A _4834_/C _4618_/Y vssd1 vssd1 vccd1 vccd1 _4620_/A sky130_fd_sc_hd__o21a_1
XFILLER_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4970_ _4966_/X _4966_/A _4979_/S vssd1 vssd1 vccd1 vccd1 _4970_/X sky130_fd_sc_hd__mux2_1
XFILLER_51_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3921_ _4446_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _3921_/Y sky130_fd_sc_hd__nand2_1
X_3852_ _5136_/Q _3849_/X _3844_/X _3851_/Y vssd1 vssd1 vccd1 vccd1 _5136_/D sky130_fd_sc_hd__o211a_1
X_2803_ _2978_/A _2803_/B vssd1 vssd1 vccd1 vccd1 _2966_/A sky130_fd_sc_hd__nand2_1
X_3783_ _3822_/A vssd1 vssd1 vccd1 vccd1 _3783_/X sky130_fd_sc_hd__clkbuf_2
X_2734_ _2943_/A _2943_/B _2733_/Y vssd1 vssd1 vccd1 vccd1 _2734_/Y sky130_fd_sc_hd__a21oi_1
X_2665_ _2666_/B _2914_/C vssd1 vssd1 vccd1 vccd1 _2675_/B sky130_fd_sc_hd__nor2_1
X_2596_ _5296_/Q _2586_/X _2582_/X _2595_/Y vssd1 vssd1 vccd1 vccd1 _5296_/D sky130_fd_sc_hd__o211a_1
X_4404_ _5113_/Q _4591_/B vssd1 vssd1 vccd1 vccd1 _4406_/A sky130_fd_sc_hd__nor2_1
X_4335_ _4513_/A _4513_/B _4334_/Y vssd1 vssd1 vccd1 vccd1 _4502_/A sky130_fd_sc_hd__o21ai_2
X_4266_ _4254_/A _4253_/A _4251_/Y _4265_/Y vssd1 vssd1 vccd1 vccd1 _4267_/A sky130_fd_sc_hd__o211a_1
XFILLER_86_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4197_ _4197_/A _4197_/B _4197_/C vssd1 vssd1 vccd1 vccd1 _5089_/D sky130_fd_sc_hd__and3_1
X_3217_ _3231_/A _3231_/C vssd1 vssd1 vccd1 vccd1 _3227_/B sky130_fd_sc_hd__and2_1
XFILLER_39_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3148_ _5179_/Q _3734_/B vssd1 vssd1 vccd1 vccd1 _3150_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3079_ _3779_/B _5163_/Q _3337_/B vssd1 vssd1 vccd1 vccd1 _3079_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4120_ _4589_/A vssd1 vssd1 vccd1 vccd1 _4910_/A sky130_fd_sc_hd__buf_1
X_4051_ _4070_/C _4051_/B vssd1 vssd1 vccd1 vccd1 _4052_/C sky130_fd_sc_hd__nand2_1
XFILLER_68_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput5 input5/A vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_1
X_3002_ _3010_/A _3002_/B vssd1 vssd1 vccd1 vccd1 _3003_/B sky130_fd_sc_hd__or2_1
XFILLER_64_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4953_ _4953_/A _5122_/Q vssd1 vssd1 vccd1 vccd1 _4958_/A sky130_fd_sc_hd__nand2_1
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3904_ _5120_/Q vssd1 vssd1 vccd1 vccd1 _3934_/B sky130_fd_sc_hd__inv_2
X_4884_ _4631_/A _4475_/X _4882_/Y _4883_/X _2837_/X vssd1 vssd1 vccd1 vccd1 _5020_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3835_ _3862_/A vssd1 vssd1 vccd1 vccd1 _3835_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3766_ _5167_/Q _3754_/X _3762_/X _3765_/Y vssd1 vssd1 vccd1 vccd1 _5167_/D sky130_fd_sc_hd__o211a_1
X_2717_ _5296_/Q _4657_/A vssd1 vssd1 vccd1 vccd1 _2957_/B sky130_fd_sc_hd__or2_2
X_3697_ _5222_/Q vssd1 vssd1 vccd1 vccd1 _3875_/B sky130_fd_sc_hd__inv_2
X_2648_ _5312_/Q _4710_/A vssd1 vssd1 vccd1 vccd1 _2857_/C sky130_fd_sc_hd__or2_2
XFILLER_59_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2579_ _5033_/Q vssd1 vssd1 vccd1 vccd1 _4818_/A sky130_fd_sc_hd__inv_2
XFILLER_59_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4318_ _4534_/A _4534_/B _4317_/Y vssd1 vssd1 vccd1 vccd1 _4523_/A sky130_fd_sc_hd__o21ai_1
X_5298_ _5301_/CLK _5298_/D vssd1 vssd1 vccd1 vccd1 _5298_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4249_ _5074_/Q vssd1 vssd1 vccd1 vccd1 _4597_/B sky130_fd_sc_hd__inv_2
XFILLER_67_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_76_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3620_ _3620_/A _3620_/B vssd1 vssd1 vccd1 vccd1 _3623_/A sky130_fd_sc_hd__nor2_1
X_3551_ _3551_/A _3551_/B vssd1 vssd1 vccd1 vccd1 _3552_/B sky130_fd_sc_hd__nor2_1
X_2502_ _5115_/Q vssd1 vssd1 vccd1 vccd1 _4911_/B sky130_fd_sc_hd__inv_2
X_3482_ _3620_/A _3620_/B _3625_/B vssd1 vssd1 vccd1 vccd1 _3482_/X sky130_fd_sc_hd__or3_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5221_ _5221_/CLK _5221_/D vssd1 vssd1 vccd1 vccd1 _5221_/Q sky130_fd_sc_hd__dfxtp_1
X_5152_ _5219_/CLK _5152_/D vssd1 vssd1 vccd1 vccd1 _5152_/Q sky130_fd_sc_hd__dfxtp_1
X_4103_ _4194_/A _4094_/X _4095_/X _3967_/A _4169_/A vssd1 vssd1 vccd1 vccd1 _4103_/Y
+ sky130_fd_sc_hd__a41oi_1
X_5083_ _5085_/CLK _5083_/D vssd1 vssd1 vccd1 vccd1 _5083_/Q sky130_fd_sc_hd__dfxtp_1
X_4034_ _4036_/A _4004_/Y _4033_/Y _4036_/B vssd1 vssd1 vccd1 vccd1 _4041_/A sky130_fd_sc_hd__o211ai_4
XFILLER_2_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4936_ _4939_/B vssd1 vssd1 vccd1 vccd1 _4940_/B sky130_fd_sc_hd__inv_2
XANTENNA_10 ANTENNA_10/DIODE vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4867_ _5023_/Q _4217_/X _4197_/B _4866_/X vssd1 vssd1 vccd1 vccd1 _5023_/D sky130_fd_sc_hd__o211a_1
X_3818_ _3820_/A _3818_/B vssd1 vssd1 vccd1 vccd1 _3818_/Y sky130_fd_sc_hd__nand2_1
X_4798_ _4798_/A _4798_/B _4792_/Y vssd1 vssd1 vccd1 vccd1 _4798_/X sky130_fd_sc_hd__or3b_1
XFILLER_21_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3749_ _3762_/A vssd1 vssd1 vccd1 vccd1 _3749_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_75_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2982_ _2981_/B _2981_/A _2969_/X vssd1 vssd1 vccd1 vccd1 _2982_/X sky130_fd_sc_hd__a21o_1
XFILLER_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4721_ _4717_/B _4719_/X _4714_/B _4720_/Y vssd1 vssd1 vccd1 vccd1 _4746_/B sky130_fd_sc_hd__a211oi_4
X_4652_ _4652_/A _4652_/B vssd1 vssd1 vccd1 vccd1 _4653_/B sky130_fd_sc_hd__nor2_1
X_3603_ _3603_/A _3603_/B vssd1 vssd1 vccd1 vccd1 _3604_/C sky130_fd_sc_hd__and2_1
X_4583_ _4581_/X _5083_/Q _5051_/Q _4440_/A vssd1 vssd1 vccd1 vccd1 _4583_/X sky130_fd_sc_hd__a31o_1
X_3534_ _5221_/Q _3199_/C _3533_/X vssd1 vssd1 vccd1 vccd1 _3534_/Y sky130_fd_sc_hd__o21ai_1
X_3465_ _3465_/A _3465_/B vssd1 vssd1 vccd1 vccd1 _3466_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5204_ _5204_/CLK _5204_/D vssd1 vssd1 vccd1 vccd1 _5204_/Q sky130_fd_sc_hd__dfxtp_1
X_3396_ _3407_/A _3406_/A vssd1 vssd1 vccd1 vccd1 _3599_/A sky130_fd_sc_hd__nor2_2
XFILLER_57_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5135_ _5196_/CLK _5135_/D vssd1 vssd1 vccd1 vccd1 _5135_/Q sky130_fd_sc_hd__dfxtp_1
X_5066_ _5096_/CLK _5066_/D vssd1 vssd1 vccd1 vccd1 _5066_/Q sky130_fd_sc_hd__dfxtp_2
X_4017_ _4017_/A _4017_/B vssd1 vssd1 vccd1 vccd1 _4022_/B sky130_fd_sc_hd__nor2_4
XFILLER_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4919_ _3898_/B _5011_/Q _3920_/A _5005_/Q _4918_/X vssd1 vssd1 vccd1 vccd1 _4920_/C
+ sky130_fd_sc_hd__o221a_1
XFILLER_20_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_87_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3250_ _3238_/Y _3154_/A _3151_/A vssd1 vssd1 vccd1 vccd1 _3250_/Y sky130_fd_sc_hd__a21oi_1
X_3181_ _5282_/Q vssd1 vssd1 vccd1 vccd1 _3717_/B sky130_fd_sc_hd__inv_2
XFILLER_39_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4704_ _4704_/A _4704_/B vssd1 vssd1 vccd1 vccd1 _4705_/B sky130_fd_sc_hd__nor2_1
X_2965_ _5264_/Q _2939_/X _2961_/X _2964_/X vssd1 vssd1 vccd1 vccd1 _5264_/D sky130_fd_sc_hd__o211a_1
XFILLER_30_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2896_ _2903_/B _2882_/B _2764_/X vssd1 vssd1 vccd1 vccd1 _2896_/Y sky130_fd_sc_hd__a21oi_1
X_4635_ _5019_/Q _5051_/Q vssd1 vssd1 vccd1 vccd1 _4880_/A sky130_fd_sc_hd__nand2_1
X_4566_ _4530_/X _5055_/Q _4540_/X _4565_/Y vssd1 vssd1 vccd1 vccd1 _5055_/D sky130_fd_sc_hd__o211a_1
X_3517_ _3517_/A _3517_/B vssd1 vssd1 vccd1 vccd1 _3572_/B sky130_fd_sc_hd__nand2_1
X_4497_ _4497_/A _4497_/B vssd1 vssd1 vccd1 vccd1 _4497_/Y sky130_fd_sc_hd__nor2_1
X_3448_ _5133_/Q _3858_/B vssd1 vssd1 vccd1 vccd1 _3450_/A sky130_fd_sc_hd__nor2_1
XFILLER_76_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3379_ _3807_/B _5152_/Q vssd1 vssd1 vccd1 vccd1 _3380_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5118_ _5118_/CLK _5118_/D vssd1 vssd1 vccd1 vccd1 _5118_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5049_ _5196_/CLK _5049_/D vssd1 vssd1 vccd1 vccd1 _5049_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_40_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2750_ _2927_/A _2930_/B _2674_/A vssd1 vssd1 vccd1 vccd1 _2750_/X sky130_fd_sc_hd__or3b_1
X_2681_ _5294_/Q _4846_/A vssd1 vssd1 vccd1 vccd1 _2712_/A sky130_fd_sc_hd__or2_2
XFILLER_8_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4420_ _4780_/B vssd1 vssd1 vccd1 vccd1 _4420_/X sky130_fd_sc_hd__clkbuf_2
X_4351_ _5068_/Q vssd1 vssd1 vccd1 vccd1 _4682_/B sky130_fd_sc_hd__inv_2
X_4282_ _4282_/A _4623_/B vssd1 vssd1 vccd1 vccd1 _4306_/B sky130_fd_sc_hd__nor2_1
X_3302_ _3301_/B _3301_/A _3292_/X vssd1 vssd1 vccd1 vccd1 _3302_/X sky130_fd_sc_hd__a21o_1
XFILLER_86_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3233_ _5246_/Q vssd1 vssd1 vccd1 vccd1 _3813_/B sky130_fd_sc_hd__inv_2
XFILLER_79_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3164_ _3164_/A _3237_/A _3164_/C vssd1 vssd1 vccd1 vccd1 _3165_/A sky130_fd_sc_hd__nor3_2
XFILLER_27_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3095_ _5259_/Q _3095_/B vssd1 vssd1 vccd1 vccd1 _3335_/A sky130_fd_sc_hd__nor2_1
XFILLER_22_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3997_ _4994_/Q _3997_/B vssd1 vssd1 vccd1 vccd1 _4031_/B sky130_fd_sc_hd__nor2_4
XFILLER_10_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2948_ _5267_/Q _2924_/X _2946_/Y _2947_/X _2899_/X vssd1 vssd1 vccd1 vccd1 _5267_/D
+ sky130_fd_sc_hd__o221a_1
X_4618_ _4832_/B vssd1 vssd1 vccd1 vccd1 _4618_/Y sky130_fd_sc_hd__inv_2
X_2879_ _2877_/X _2874_/A _2878_/X vssd1 vssd1 vccd1 vccd1 _2879_/X sky130_fd_sc_hd__a21o_1
X_4549_ _4549_/A _4549_/B _4549_/C vssd1 vssd1 vccd1 vccd1 _4549_/X sky130_fd_sc_hd__and3_1
XFILLER_49_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3920_ _3920_/A vssd1 vssd1 vccd1 vccd1 _4930_/B sky130_fd_sc_hd__buf_1
XFILLER_51_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3851_ _3860_/A _3851_/B vssd1 vssd1 vccd1 vccd1 _3851_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2802_ _2802_/A _2979_/A vssd1 vssd1 vccd1 vccd1 _2803_/B sky130_fd_sc_hd__nor2_1
X_3782_ _5162_/Q _3768_/X _3778_/X _3781_/Y vssd1 vssd1 vccd1 vccd1 _5162_/D sky130_fd_sc_hd__o211a_1
X_2733_ _2946_/A _2949_/A vssd1 vssd1 vccd1 vccd1 _2733_/Y sky130_fd_sc_hd__nand2_1
X_2664_ _5304_/Q _4691_/A vssd1 vssd1 vccd1 vccd1 _2914_/C sky130_fd_sc_hd__or2_2
X_2595_ _2602_/A _4657_/A vssd1 vssd1 vccd1 vccd1 _2595_/Y sky130_fd_sc_hd__nand2_1
X_4403_ _4423_/A vssd1 vssd1 vccd1 vccd1 _4403_/Y sky130_fd_sc_hd__inv_2
X_4334_ _4520_/B _4516_/A vssd1 vssd1 vccd1 vccd1 _4334_/Y sky130_fd_sc_hd__nor2_1
X_4265_ _4367_/A _4265_/B vssd1 vssd1 vccd1 vccd1 _4265_/Y sky130_fd_sc_hd__nand2_1
X_4196_ _4106_/A _4201_/C _4304_/A vssd1 vssd1 vccd1 vccd1 _4197_/C sky130_fd_sc_hd__o21ai_1
X_3216_ _5250_/Q _3210_/X _3214_/X _3215_/Y _3208_/X vssd1 vssd1 vccd1 vccd1 _5250_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_27_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3147_ _5275_/Q vssd1 vssd1 vccd1 vccd1 _3734_/B sky130_fd_sc_hd__inv_2
XFILLER_82_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3078_ _5162_/Q _3781_/B vssd1 vssd1 vccd1 vccd1 _3337_/B sky130_fd_sc_hd__or2_2
XFILLER_82_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4050_ _4056_/B _4045_/C _4045_/B vssd1 vssd1 vccd1 vccd1 _4070_/C sky130_fd_sc_hd__a21o_2
XFILLER_1_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 input6/A vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_1
XFILLER_76_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3001_ _3001_/A _2997_/C vssd1 vssd1 vccd1 vccd1 _3003_/A sky130_fd_sc_hd__or2b_1
XFILLER_36_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4952_ _5122_/Q _4953_/A vssd1 vssd1 vccd1 vccd1 _4955_/C sky130_fd_sc_hd__or2_1
XFILLER_64_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3903_ _3887_/X _4974_/X _3893_/X _3902_/Y vssd1 vssd1 vccd1 vccd1 _5121_/D sky130_fd_sc_hd__o211a_1
X_4883_ _4882_/B _4882_/A _3907_/A vssd1 vssd1 vccd1 vccd1 _4883_/X sky130_fd_sc_hd__a21o_1
XFILLER_51_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3834_ _5142_/Q _3822_/X _3830_/X _3833_/Y vssd1 vssd1 vccd1 vccd1 _5142_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3765_ _3765_/A _3765_/B vssd1 vssd1 vccd1 vccd1 _3765_/Y sky130_fd_sc_hd__nand2_1
X_2716_ _2708_/Y _2710_/Y _2804_/A vssd1 vssd1 vccd1 vccd1 _2716_/Y sky130_fd_sc_hd__a21oi_1
X_3696_ _5192_/Q _3650_/X _3692_/X _3694_/X _3695_/X vssd1 vssd1 vccd1 vccd1 _5192_/D
+ sky130_fd_sc_hd__o221a_1
X_2647_ _4755_/A _5313_/Q vssd1 vssd1 vccd1 vccd1 _2653_/B sky130_fd_sc_hd__and2_1
XFILLER_10_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2578_ _5301_/Q _2567_/X _2563_/X _2577_/Y vssd1 vssd1 vccd1 vccd1 _5301_/D sky130_fd_sc_hd__o211a_1
X_4317_ _4541_/B _4537_/A vssd1 vssd1 vccd1 vccd1 _4317_/Y sky130_fd_sc_hd__nor2_1
X_5297_ _5301_/CLK _5297_/D vssd1 vssd1 vccd1 vccd1 _5297_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_19_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4248_ _4462_/B vssd1 vssd1 vccd1 vccd1 _4253_/A sky130_fd_sc_hd__inv_2
XFILLER_74_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4179_ _5091_/Q _5090_/Q _5089_/Q vssd1 vssd1 vccd1 vccd1 _4180_/C sky130_fd_sc_hd__and3_1
XFILLER_27_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3550_ _3550_/A _3550_/B vssd1 vssd1 vccd1 vccd1 _3552_/A sky130_fd_sc_hd__nor2_1
X_2501_ _5015_/Q vssd1 vssd1 vccd1 vccd1 _4199_/A sky130_fd_sc_hd__inv_2
X_3481_ _3622_/B _3481_/B vssd1 vssd1 vccd1 vccd1 _3625_/B sky130_fd_sc_hd__nand2_1
X_5220_ _5250_/CLK _5220_/D vssd1 vssd1 vccd1 vccd1 _5220_/Q sky130_fd_sc_hd__dfxtp_1
X_5151_ _5221_/CLK _5151_/D vssd1 vssd1 vccd1 vccd1 _5151_/Q sky130_fd_sc_hd__dfxtp_1
X_5082_ _5108_/CLK _5082_/D vssd1 vssd1 vccd1 vccd1 _5082_/Q sky130_fd_sc_hd__dfxtp_1
X_4102_ _4202_/B vssd1 vssd1 vccd1 vccd1 _4194_/A sky130_fd_sc_hd__buf_2
X_4033_ _4030_/Y _4045_/B _4032_/Y vssd1 vssd1 vccd1 vccd1 _4033_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_56_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4935_ _5118_/Q _5117_/Q _5116_/Q vssd1 vssd1 vccd1 vccd1 _4939_/B sky130_fd_sc_hd__and3_1
X_4866_ _4865_/X _4862_/A _4588_/A vssd1 vssd1 vccd1 vccd1 _4866_/X sky130_fd_sc_hd__a21o_1
X_4797_ _4797_/A _4797_/B vssd1 vssd1 vccd1 vccd1 _4798_/B sky130_fd_sc_hd__nor2_1
X_3817_ _3830_/A vssd1 vssd1 vccd1 vccd1 _3817_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3748_ _5174_/Q _3741_/X _3736_/X _3747_/Y vssd1 vssd1 vccd1 vccd1 _5174_/D sky130_fd_sc_hd__o211a_1
X_3679_ _3679_/A _3679_/B vssd1 vssd1 vccd1 vccd1 _3679_/Y sky130_fd_sc_hd__nor2_1
XFILLER_87_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2981_ _2981_/A _2981_/B vssd1 vssd1 vccd1 vccd1 _2981_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_41_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5317_/CLK sky130_fd_sc_hd__clkbuf_16
X_4720_ _4720_/A _4720_/B vssd1 vssd1 vccd1 vccd1 _4720_/Y sky130_fd_sc_hd__nor2_2
X_4651_ _5028_/Q _5060_/Q vssd1 vssd1 vccd1 vccd1 _4653_/A sky130_fd_sc_hd__nor2_1
Xinput20 phase_in[7] vssd1 vssd1 vccd1 vccd1 hold45/A sky130_fd_sc_hd__clkbuf_1
X_3602_ _3603_/B _3603_/A vssd1 vssd1 vccd1 vccd1 _3604_/B sky130_fd_sc_hd__nor2_1
X_4582_ _4587_/B _5051_/Q _4581_/X vssd1 vssd1 vccd1 vccd1 _4582_/Y sky130_fd_sc_hd__a21oi_1
X_3533_ _4132_/A vssd1 vssd1 vccd1 vccd1 _3533_/X sky130_fd_sc_hd__clkbuf_4
X_3464_ _3847_/B _5137_/Q vssd1 vssd1 vccd1 vccd1 _3465_/B sky130_fd_sc_hd__and2_1
X_5203_ _5204_/CLK _5203_/D vssd1 vssd1 vccd1 vccd1 _5203_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5134_ _5199_/CLK _5134_/D vssd1 vssd1 vccd1 vccd1 _5134_/Q sky130_fd_sc_hd__dfxtp_1
X_3395_ _3826_/B _5145_/Q vssd1 vssd1 vccd1 vccd1 _3406_/A sky130_fd_sc_hd__and2_1
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5065_ _5096_/CLK _5065_/D vssd1 vssd1 vccd1 vccd1 _5065_/Q sky130_fd_sc_hd__dfxtp_1
X_4016_ _4016_/A vssd1 vssd1 vccd1 vccd1 _4017_/B sky130_fd_sc_hd__inv_2
XFILLER_25_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4918_ _5125_/Q _3937_/Y _5123_/Q _3935_/Y vssd1 vssd1 vccd1 vccd1 _4918_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5221_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_32_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4849_ _4849_/A _4849_/B vssd1 vssd1 vccd1 vccd1 _4855_/A sky130_fd_sc_hd__and2_1
XFILLER_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_23_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 _5267_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3180_ _5282_/Q _3211_/B _3048_/X _3179_/Y vssd1 vssd1 vccd1 vccd1 _3180_/Y sky130_fd_sc_hd__o22ai_4
XFILLER_66_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2964_ _2962_/X _2957_/A _2963_/X vssd1 vssd1 vccd1 vccd1 _2964_/X sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_14_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5002_/CLK sky130_fd_sc_hd__clkbuf_16
X_4703_ _5044_/Q _5076_/Q vssd1 vssd1 vccd1 vccd1 _4705_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2895_ _5276_/Q _2625_/X _2892_/X _2894_/X vssd1 vssd1 vccd1 vccd1 _5276_/D sky130_fd_sc_hd__o211a_1
X_4634_ _5020_/Q _4634_/B vssd1 vssd1 vccd1 vccd1 _4881_/B sky130_fd_sc_hd__nand2_1
XFILLER_30_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4565_ _4564_/Y _4559_/X _4778_/A vssd1 vssd1 vccd1 vccd1 _4565_/Y sky130_fd_sc_hd__o21ai_1
X_3516_ _3813_/B _5150_/Q vssd1 vssd1 vccd1 vccd1 _3517_/B sky130_fd_sc_hd__nand2_1
X_4496_ _4496_/A _4496_/B vssd1 vssd1 vccd1 vccd1 _4497_/B sky130_fd_sc_hd__and2_1
X_3447_ _5229_/Q vssd1 vssd1 vccd1 vccd1 _3858_/B sky130_fd_sc_hd__inv_2
XFILLER_69_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3378_ _5152_/Q _3807_/B vssd1 vssd1 vccd1 vccd1 _3391_/B sky130_fd_sc_hd__or2_2
XFILLER_69_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5117_ _5118_/CLK _5117_/D vssd1 vssd1 vccd1 vccd1 _5117_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5048_ _5317_/CLK _5048_/D vssd1 vssd1 vccd1 vccd1 _5048_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2680_ _4652_/A _5295_/Q vssd1 vssd1 vccd1 vccd1 _2714_/B sky130_fd_sc_hd__and2_1
XFILLER_8_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4350_ _5100_/Q _5068_/Q vssd1 vssd1 vccd1 vccd1 _4494_/A sky130_fd_sc_hd__nor2_1
X_3301_ _3301_/A _3301_/B vssd1 vssd1 vccd1 vccd1 _3301_/Y sky130_fd_sc_hd__nor2_1
X_4281_ _5058_/Q vssd1 vssd1 vccd1 vccd1 _4623_/B sky130_fd_sc_hd__inv_2
XFILLER_86_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_3_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5076_/CLK sky130_fd_sc_hd__clkbuf_16
X_3232_ _3232_/A _3232_/B vssd1 vssd1 vccd1 vccd1 _3232_/Y sky130_fd_sc_hd__nor2_1
XFILLER_79_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3163_ _3241_/B _3241_/A _3247_/B vssd1 vssd1 vccd1 vccd1 _3164_/C sky130_fd_sc_hd__or3_1
XFILLER_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3094_ _5163_/Q vssd1 vssd1 vccd1 vccd1 _3095_/B sky130_fd_sc_hd__inv_2
XFILLER_39_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3996_ _3997_/B _4994_/Q vssd1 vssd1 vccd1 vccd1 _4031_/A sky130_fd_sc_hd__and2_1
XFILLER_22_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2947_ _2946_/B _2946_/A _2848_/X vssd1 vssd1 vccd1 vccd1 _2947_/X sky130_fd_sc_hd__a21o_1
XFILLER_13_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4617_ _4835_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4832_/B sky130_fd_sc_hd__nor2_2
X_2878_ _3361_/A vssd1 vssd1 vccd1 vccd1 _2878_/X sky130_fd_sc_hd__buf_2
X_4548_ _4549_/A _4549_/C _4549_/B vssd1 vssd1 vccd1 vccd1 _4548_/Y sky130_fd_sc_hd__a21oi_1
X_4479_ _4479_/A _4479_/B vssd1 vssd1 vccd1 vccd1 _4499_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3850_ _3863_/A vssd1 vssd1 vccd1 vccd1 _3860_/A sky130_fd_sc_hd__buf_1
XFILLER_32_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2801_ _2801_/A vssd1 vssd1 vccd1 vccd1 _2979_/A sky130_fd_sc_hd__inv_2
X_3781_ _3781_/A _3781_/B vssd1 vssd1 vccd1 vccd1 _3781_/Y sky130_fd_sc_hd__nand2_1
X_2732_ _2950_/A vssd1 vssd1 vccd1 vccd1 _2949_/A sky130_fd_sc_hd__inv_2
X_2663_ _4677_/A _5305_/Q vssd1 vssd1 vccd1 vccd1 _2666_/B sky130_fd_sc_hd__and2_1
X_2594_ _5029_/Q vssd1 vssd1 vccd1 vccd1 _4657_/A sky130_fd_sc_hd__inv_2
X_4402_ _4402_/A _4725_/B vssd1 vssd1 vccd1 vccd1 _4423_/A sky130_fd_sc_hd__nor2_4
X_4333_ _4333_/A vssd1 vssd1 vccd1 vccd1 _4516_/A sky130_fd_sc_hd__inv_2
X_4264_ _4259_/Y _4457_/A _4364_/A vssd1 vssd1 vccd1 vccd1 _4265_/B sky130_fd_sc_hd__a21oi_1
X_3215_ _3048_/X _3213_/Y _3179_/Y _2888_/X vssd1 vssd1 vccd1 vccd1 _3215_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_39_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4195_ _4194_/A _4190_/B _4197_/A _4282_/A _4734_/A vssd1 vssd1 vccd1 vccd1 _5090_/D
+ sky130_fd_sc_hd__a221oi_2
X_3146_ _3257_/A _3257_/B _3145_/X vssd1 vssd1 vccd1 vccd1 _3236_/B sky130_fd_sc_hd__a21oi_2
XFILLER_54_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3077_ _5258_/Q vssd1 vssd1 vccd1 vccd1 _3781_/B sky130_fd_sc_hd__inv_2
XFILLER_82_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3979_ _4990_/Q _4990_/D vssd1 vssd1 vccd1 vccd1 _3980_/B sky130_fd_sc_hd__and2_1
XFILLER_10_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 input7/A vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_1
X_3000_ _3000_/A _3000_/B vssd1 vssd1 vccd1 vccd1 _3001_/A sky130_fd_sc_hd__nor2_1
XFILLER_76_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4951_ _4951_/A _4951_/B vssd1 vssd1 vccd1 vccd1 _4951_/X sky130_fd_sc_hd__and2_1
X_3902_ _3916_/A _4948_/A vssd1 vssd1 vccd1 vccd1 _3902_/Y sky130_fd_sc_hd__nand2_1
X_4882_ _4882_/A _4882_/B vssd1 vssd1 vccd1 vccd1 _4882_/Y sky130_fd_sc_hd__nor2_1
X_3833_ _3833_/A _3833_/B vssd1 vssd1 vccd1 vccd1 _3833_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3764_ _5168_/Q _3754_/X _3762_/X _3763_/Y vssd1 vssd1 vccd1 vccd1 _5168_/D sky130_fd_sc_hd__o211a_1
X_2715_ _2715_/A _2968_/A vssd1 vssd1 vccd1 vccd1 _2804_/A sky130_fd_sc_hd__nand2_1
X_3695_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3695_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_10_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2646_ _5313_/Q _4755_/A vssd1 vssd1 vccd1 vccd1 _2661_/A sky130_fd_sc_hd__nor2_1
X_2577_ _2584_/A _4815_/A vssd1 vssd1 vccd1 vccd1 _2577_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4316_ _4316_/A _4316_/B vssd1 vssd1 vccd1 vccd1 _4537_/A sky130_fd_sc_hd__or2_1
X_5296_ _5301_/CLK _5296_/D vssd1 vssd1 vccd1 vccd1 _5296_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4247_ _4252_/A _4594_/B vssd1 vssd1 vccd1 vccd1 _4462_/B sky130_fd_sc_hd__nor2_2
XFILLER_55_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4178_ _5095_/Q _4174_/A _4177_/X vssd1 vssd1 vccd1 vccd1 _5095_/D sky130_fd_sc_hd__o21a_1
XFILLER_82_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3129_ _5269_/Q vssd1 vssd1 vccd1 vccd1 _3750_/B sky130_fd_sc_hd__inv_2
XFILLER_35_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_76_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3480_ _3839_/B _5140_/Q vssd1 vssd1 vccd1 vccd1 _3481_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5150_ _5221_/CLK _5150_/D vssd1 vssd1 vccd1 vccd1 _5150_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_69_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5081_ _5197_/CLK _5081_/D vssd1 vssd1 vccd1 vccd1 _5081_/Q sky130_fd_sc_hd__dfxtp_1
X_4101_ _4127_/B _4101_/B _4119_/C vssd1 vssd1 vccd1 vccd1 _4101_/Y sky130_fd_sc_hd__nor3_2
X_4032_ _4032_/A vssd1 vssd1 vccd1 vccd1 _4032_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_1_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 clkbuf_2_3_0_clk/A sky130_fd_sc_hd__clkbuf_1
XFILLER_2_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4934_ _4951_/A _4934_/B vssd1 vssd1 vccd1 vccd1 _4934_/X sky130_fd_sc_hd__and2_1
XFILLER_24_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4865_ _4865_/A _4865_/B vssd1 vssd1 vccd1 vccd1 _4865_/X sky130_fd_sc_hd__or2_1
XFILLER_32_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3816_ _5149_/Q _3809_/X _3804_/X _3815_/Y vssd1 vssd1 vccd1 vccd1 _5149_/D sky130_fd_sc_hd__o211a_1
X_4796_ _5038_/Q _4770_/X _4794_/Y _4795_/X _4785_/X vssd1 vssd1 vccd1 vccd1 _5038_/D
+ sky130_fd_sc_hd__o221a_1
X_3747_ _3752_/A _3747_/B vssd1 vssd1 vccd1 vccd1 _3747_/Y sky130_fd_sc_hd__nand2_1
X_3678_ _3678_/A vssd1 vssd1 vccd1 vccd1 _3679_/B sky130_fd_sc_hd__inv_2
X_2629_ _3713_/A _4633_/A vssd1 vssd1 vccd1 vccd1 _2629_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5279_ _5280_/CLK _5279_/D vssd1 vssd1 vccd1 vccd1 _5279_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2980_ _2980_/A vssd1 vssd1 vccd1 vccd1 _2981_/B sky130_fd_sc_hd__inv_2
XFILLER_14_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4650_ _4650_/A _4650_/B vssd1 vssd1 vccd1 vccd1 _4845_/A sky130_fd_sc_hd__nand2_1
Xinput21 phase_in[8] vssd1 vssd1 vccd1 vccd1 hold43/A sky130_fd_sc_hd__clkbuf_1
Xinput10 hold30/X vssd1 vssd1 vccd1 vccd1 hold29/A sky130_fd_sc_hd__clkbuf_1
X_3601_ _5209_/Q _3596_/X _3599_/Y _3600_/X _3591_/X vssd1 vssd1 vccd1 vccd1 _5209_/D
+ sky130_fd_sc_hd__o221a_1
X_4581_ _4581_/A _4581_/B vssd1 vssd1 vccd1 vccd1 _4581_/X sky130_fd_sc_hd__or2_1
X_3532_ _3541_/B _3531_/Y _3605_/A vssd1 vssd1 vccd1 vccd1 _3532_/Y sky130_fd_sc_hd__a21oi_1
X_3463_ _5137_/Q _3847_/B vssd1 vssd1 vccd1 vccd1 _3465_/A sky130_fd_sc_hd__nor2_1
XFILLER_6_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5202_ _5204_/CLK _5202_/D vssd1 vssd1 vccd1 vccd1 _5202_/Q sky130_fd_sc_hd__dfxtp_1
X_5133_ _5196_/CLK _5133_/D vssd1 vssd1 vccd1 vccd1 _5133_/Q sky130_fd_sc_hd__dfxtp_1
X_3394_ _5145_/Q _3826_/B vssd1 vssd1 vccd1 vccd1 _3407_/A sky130_fd_sc_hd__nor2_2
XFILLER_69_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5064_ _5096_/CLK _5064_/D vssd1 vssd1 vccd1 vccd1 _5064_/Q sky130_fd_sc_hd__dfxtp_1
X_4015_ _4037_/C _4015_/B vssd1 vssd1 vccd1 vccd1 _4015_/Y sky130_fd_sc_hd__nand2_1
XFILLER_65_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4917_ _5120_/Q _3938_/Y _5119_/Q _3931_/Y _4916_/X vssd1 vssd1 vccd1 vccd1 _4920_/B
+ sky130_fd_sc_hd__o221a_1
X_4848_ _4848_/A vssd1 vssd1 vccd1 vccd1 _4855_/B sky130_fd_sc_hd__inv_2
XFILLER_20_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4779_ _4779_/A _4779_/B vssd1 vssd1 vccd1 vccd1 _4780_/C sky130_fd_sc_hd__nand2_1
XFILLER_4_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2963_ _3615_/A vssd1 vssd1 vccd1 vccd1 _2963_/X sky130_fd_sc_hd__buf_2
X_4702_ _4762_/B _4702_/B vssd1 vssd1 vccd1 vccd1 _4761_/A sky130_fd_sc_hd__nand2_1
X_2894_ _2884_/X _2893_/Y _2878_/X vssd1 vssd1 vccd1 vccd1 _2894_/X sky130_fd_sc_hd__a21o_1
X_4633_ _4633_/A _4633_/B vssd1 vssd1 vccd1 vccd1 _4878_/C sky130_fd_sc_hd__nand2_1
X_4564_ _4559_/A _4571_/C _4559_/C vssd1 vssd1 vccd1 vccd1 _4564_/Y sky130_fd_sc_hd__a21oi_1
X_3515_ _3568_/A vssd1 vssd1 vccd1 vccd1 _3517_/A sky130_fd_sc_hd__inv_2
X_4495_ _4496_/A _4497_/A _4496_/B _3879_/A vssd1 vssd1 vccd1 vccd1 _4495_/X sky130_fd_sc_hd__a31o_1
X_3446_ _3663_/B _3446_/B vssd1 vssd1 vccd1 vccd1 _3670_/B sky130_fd_sc_hd__nand2_1
XFILLER_69_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3377_ _5248_/Q vssd1 vssd1 vccd1 vccd1 _3807_/B sky130_fd_sc_hd__inv_2
XFILLER_84_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5116_ _5118_/CLK _5116_/D vssd1 vssd1 vccd1 vccd1 _5116_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5047_ _5317_/CLK _5047_/D vssd1 vssd1 vccd1 vccd1 _5047_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_72_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3300_ _3300_/A _3300_/B vssd1 vssd1 vccd1 vccd1 _3301_/B sky130_fd_sc_hd__nand2_1
X_4280_ _5089_/Q _5057_/Q vssd1 vssd1 vccd1 vccd1 _4549_/C sky130_fd_sc_hd__nand2_1
XFILLER_3_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3231_ _3231_/A _3231_/B _3231_/C vssd1 vssd1 vccd1 vccd1 _3232_/A sky130_fd_sc_hd__and3_1
X_3162_ _3243_/B _3162_/B vssd1 vssd1 vccd1 vccd1 _3247_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3093_ _3341_/A _3345_/A _3341_/B vssd1 vssd1 vccd1 vccd1 _3333_/A sky130_fd_sc_hd__a21oi_4
XFILLER_62_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3995_ _4994_/D vssd1 vssd1 vccd1 vccd1 _3997_/B sky130_fd_sc_hd__inv_2
XFILLER_22_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2946_ _2946_/A _2946_/B vssd1 vssd1 vccd1 vccd1 _2946_/Y sky130_fd_sc_hd__nor2_1
X_2877_ _2874_/B _2871_/C _2871_/A vssd1 vssd1 vccd1 vccd1 _2877_/X sky130_fd_sc_hd__a21o_1
X_4616_ _5029_/Q _5061_/Q vssd1 vssd1 vccd1 vccd1 _4834_/C sky130_fd_sc_hd__nand2_1
X_4547_ _4553_/B _4553_/A vssd1 vssd1 vccd1 vccd1 _4549_/A sky130_fd_sc_hd__or2_1
X_4478_ _4478_/A vssd1 vssd1 vccd1 vccd1 _4483_/A sky130_fd_sc_hd__inv_2
XFILLER_89_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3429_ _5126_/Q vssd1 vssd1 vccd1 vccd1 _3429_/Y sky130_fd_sc_hd__inv_2
XFILLER_57_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_79_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_76_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2800_ _2687_/Y _2989_/A _2799_/X vssd1 vssd1 vccd1 vccd1 _2978_/A sky130_fd_sc_hd__o21bai_1
X_3780_ _5163_/Q _3768_/X _3778_/X _3779_/Y vssd1 vssd1 vccd1 vccd1 _5163_/D sky130_fd_sc_hd__o211a_1
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2731_ _2731_/A _2731_/B vssd1 vssd1 vccd1 vccd1 _2950_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4401_ _5080_/Q vssd1 vssd1 vccd1 vccd1 _4725_/B sky130_fd_sc_hd__inv_2
X_2662_ _5305_/Q _4677_/A vssd1 vssd1 vccd1 vccd1 _2675_/A sky130_fd_sc_hd__nor2_1
X_2593_ _5297_/Q _2586_/X _2582_/X _2592_/Y vssd1 vssd1 vccd1 vccd1 _5297_/D sky130_fd_sc_hd__o211a_1
X_4332_ _4332_/A _4332_/B vssd1 vssd1 vccd1 vccd1 _4333_/A sky130_fd_sc_hd__nor2_1
X_4263_ _5104_/Q _5072_/Q vssd1 vssd1 vccd1 vccd1 _4364_/A sky130_fd_sc_hd__nor2_1
X_3214_ _3048_/X _3179_/Y _3213_/Y vssd1 vssd1 vccd1 vccd1 _3214_/X sky130_fd_sc_hd__o21a_1
XFILLER_79_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4194_ _4194_/A _5089_/Q vssd1 vssd1 vccd1 vccd1 _4197_/A sky130_fd_sc_hd__nand2_1
X_3145_ _3266_/B _3145_/B _3145_/C vssd1 vssd1 vccd1 vccd1 _3145_/X sky130_fd_sc_hd__or3_1
XFILLER_39_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3076_ _3076_/A _3108_/A vssd1 vssd1 vccd1 vccd1 _3298_/A sky130_fd_sc_hd__nand2_1
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3978_ _4990_/Q _4990_/D vssd1 vssd1 vccd1 vccd1 _3980_/A sky130_fd_sc_hd__nor2_1
XFILLER_10_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2929_ _5271_/Q _2924_/X _2927_/Y _2928_/X _2899_/X vssd1 vssd1 vccd1 vccd1 _5271_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_50_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 input8/A vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_1
XFILLER_39_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4950_ _4953_/A _4950_/B vssd1 vssd1 vccd1 vccd1 _4951_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3901_ _5121_/Q vssd1 vssd1 vccd1 vccd1 _4948_/A sky130_fd_sc_hd__inv_2
X_4881_ _4881_/A _4881_/B vssd1 vssd1 vccd1 vccd1 _4882_/B sky130_fd_sc_hd__nand2_1
X_3832_ _5143_/Q _3822_/X _3830_/X _3831_/Y vssd1 vssd1 vccd1 vccd1 _5143_/D sky130_fd_sc_hd__o211a_1
X_3763_ _3765_/A _3763_/B vssd1 vssd1 vccd1 vccd1 _3763_/Y sky130_fd_sc_hd__nand2_1
X_2714_ _2714_/A _2714_/B vssd1 vssd1 vccd1 vccd1 _2968_/A sky130_fd_sc_hd__nor2_2
X_3694_ _3691_/A _3691_/B _3693_/X vssd1 vssd1 vccd1 vccd1 _3694_/X sky130_fd_sc_hd__o21ba_1
X_2645_ _5314_/Q vssd1 vssd1 vccd1 vccd1 _2842_/B sky130_fd_sc_hd__inv_2
X_2576_ _5034_/Q vssd1 vssd1 vccd1 vccd1 _4815_/A sky130_fd_sc_hd__inv_2
X_4315_ _4315_/A _4652_/B vssd1 vssd1 vccd1 vccd1 _4316_/B sky130_fd_sc_hd__nor2_1
XFILLER_87_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5295_ _5301_/CLK _5295_/D vssd1 vssd1 vccd1 vccd1 _5295_/Q sky130_fd_sc_hd__dfxtp_1
X_4246_ _5073_/Q vssd1 vssd1 vccd1 vccd1 _4594_/B sky130_fd_sc_hd__inv_2
X_4177_ _4326_/A _4183_/A _2889_/X vssd1 vssd1 vccd1 vccd1 _4177_/X sky130_fd_sc_hd__o21a_1
XFILLER_82_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3128_ _5268_/Q _5172_/Q vssd1 vssd1 vccd1 vccd1 _3284_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3059_ _5175_/Q _3745_/B vssd1 vssd1 vccd1 vccd1 _3143_/A sky130_fd_sc_hd__nor2_1
XPHY_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_73_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5080_ _5197_/CLK _5080_/D vssd1 vssd1 vccd1 vccd1 _5080_/Q sky130_fd_sc_hd__dfxtp_1
X_4100_ _4402_/A _4244_/A _4100_/C vssd1 vssd1 vccd1 vccd1 _4101_/B sky130_fd_sc_hd__or3_1
X_4031_ _4031_/A _4031_/B _4031_/C _4031_/D vssd1 vssd1 vccd1 vccd1 _4045_/B sky130_fd_sc_hd__or4_4
XFILLER_2_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4933_ _4966_/B vssd1 vssd1 vccd1 vccd1 _4951_/A sky130_fd_sc_hd__buf_1
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4864_ _4528_/A _4861_/Y _4862_/X _2510_/X _4863_/Y vssd1 vssd1 vccd1 vccd1 _5024_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3815_ _3820_/A _3815_/B vssd1 vssd1 vccd1 vccd1 _3815_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4795_ _4794_/B _4794_/A _4764_/X vssd1 vssd1 vccd1 vccd1 _4795_/X sky130_fd_sc_hd__a21o_1
X_3746_ _5175_/Q _3741_/X _3736_/X _3745_/Y vssd1 vssd1 vccd1 vccd1 _5175_/D sky130_fd_sc_hd__o211a_1
X_3677_ _3677_/A _3677_/B vssd1 vssd1 vccd1 vccd1 _3678_/A sky130_fd_sc_hd__nand2_1
X_2628_ _5021_/Q vssd1 vssd1 vccd1 vccd1 _4633_/A sky130_fd_sc_hd__inv_2
X_2559_ _5038_/Q vssd1 vssd1 vccd1 vccd1 _4677_/A sky130_fd_sc_hd__inv_2
X_5278_ _5280_/CLK _5278_/D vssd1 vssd1 vccd1 vccd1 _5278_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4229_ _4221_/B _4226_/Y _4228_/Y vssd1 vssd1 vccd1 vccd1 _4229_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_46_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_70_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput22 hold22/X vssd1 vssd1 vccd1 vccd1 hold21/A sky130_fd_sc_hd__buf_1
Xinput11 hold35/X vssd1 vssd1 vccd1 vccd1 hold34/A sky130_fd_sc_hd__clkbuf_1
X_4580_ _4580_/A _4634_/B vssd1 vssd1 vccd1 vccd1 _4581_/A sky130_fd_sc_hd__nor2_1
X_3600_ _3599_/B _3599_/A _3361_/X vssd1 vssd1 vccd1 vccd1 _3600_/X sky130_fd_sc_hd__a21o_1
X_3531_ _3531_/A _3531_/B _3531_/C vssd1 vssd1 vccd1 vccd1 _3531_/Y sky130_fd_sc_hd__nor3_1
X_3462_ _5233_/Q vssd1 vssd1 vccd1 vccd1 _3847_/B sky130_fd_sc_hd__inv_2
X_3393_ _5241_/Q vssd1 vssd1 vccd1 vccd1 _3826_/B sky130_fd_sc_hd__inv_2
X_5201_ _5204_/CLK _5201_/D vssd1 vssd1 vccd1 vccd1 _5201_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5132_ _5196_/CLK _5132_/D vssd1 vssd1 vccd1 vccd1 _5132_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5063_ _5096_/CLK _5063_/D vssd1 vssd1 vccd1 vccd1 _5063_/Q sky130_fd_sc_hd__dfxtp_1
X_4014_ _3973_/Y _4016_/A _4022_/A _4022_/C vssd1 vssd1 vccd1 vccd1 _4028_/A sky130_fd_sc_hd__a22oi_4
XFILLER_80_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4916_ _5009_/Q _3934_/B _3933_/B _5014_/Q vssd1 vssd1 vccd1 vccd1 _4916_/X sky130_fd_sc_hd__o22a_1
XFILLER_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4847_ _3879_/X _4845_/Y _4807_/X _4846_/Y vssd1 vssd1 vccd1 vccd1 _5027_/D sky130_fd_sc_hd__o211a_1
X_4778_ _4778_/A _4778_/B vssd1 vssd1 vccd1 vccd1 _4778_/Y sky130_fd_sc_hd__nor2_1
X_3729_ _3755_/A vssd1 vssd1 vccd1 vccd1 _3739_/A sky130_fd_sc_hd__buf_1
XFILLER_0_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_1_0_0_clk clkbuf_0_clk/X vssd1 vssd1 vccd1 vccd1 ANTENNA_10/DIODE sky130_fd_sc_hd__clkbuf_1
XFILLER_3_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_66_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2962_ _2962_/A _2962_/B vssd1 vssd1 vccd1 vccd1 _2962_/X sky130_fd_sc_hd__or2_1
XFILLER_22_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4701_ _4701_/A _4701_/B vssd1 vssd1 vccd1 vccd1 _4702_/B sky130_fd_sc_hd__nand2_1
X_4632_ _5053_/Q vssd1 vssd1 vccd1 vccd1 _4633_/B sky130_fd_sc_hd__inv_2
X_2893_ _2893_/A _2893_/B vssd1 vssd1 vccd1 vccd1 _2893_/Y sky130_fd_sc_hd__nand2_1
X_4563_ _4492_/X _5056_/Q _4561_/Y _4562_/X _4508_/X vssd1 vssd1 vccd1 vccd1 _5056_/D
+ sky130_fd_sc_hd__o221a_1
X_3514_ _3503_/B _3511_/Y _3513_/X _3509_/B vssd1 vssd1 vccd1 vccd1 _3572_/C sky130_fd_sc_hd__o22a_2
X_4494_ _4494_/A _4494_/B vssd1 vssd1 vccd1 vccd1 _4497_/A sky130_fd_sc_hd__nor2_1
X_3445_ _3860_/B _5132_/Q vssd1 vssd1 vccd1 vccd1 _3446_/B sky130_fd_sc_hd__nand2_1
X_3376_ _5154_/Q vssd1 vssd1 vccd1 vccd1 _3549_/B sky130_fd_sc_hd__inv_2
X_5115_ _5118_/CLK _5115_/D vssd1 vssd1 vccd1 vccd1 _5115_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5046_ _5076_/CLK _5046_/D vssd1 vssd1 vccd1 vccd1 _5046_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_68_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_84_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3230_ _5247_/Q _3210_/X _3228_/X _3229_/Y _3208_/X vssd1 vssd1 vccd1 vccd1 _5247_/D
+ sky130_fd_sc_hd__o221a_1
X_3161_ _3732_/B _5180_/Q vssd1 vssd1 vccd1 vccd1 _3162_/B sky130_fd_sc_hd__nand2_1
XFILLER_39_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3092_ _3337_/B _3092_/B vssd1 vssd1 vccd1 vccd1 _3341_/B sky130_fd_sc_hd__nand2_2
XFILLER_81_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3994_ _3994_/A _4031_/C vssd1 vssd1 vccd1 vccd1 _4000_/A sky130_fd_sc_hd__nand2_2
XFILLER_22_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _2950_/A _2950_/B _2731_/A vssd1 vssd1 vccd1 vccd1 _2946_/B sky130_fd_sc_hd__o21a_1
X_2876_ _5279_/Q _2841_/X _2873_/X _2875_/Y _4902_/A vssd1 vssd1 vccd1 vccd1 _5279_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4615_ _5030_/Q _5062_/Q vssd1 vssd1 vccd1 vccd1 _4832_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4546_ _4546_/A _4546_/B vssd1 vssd1 vccd1 vccd1 _4553_/A sky130_fd_sc_hd__and2_1
X_4477_ _4453_/X _5071_/Q _4473_/X _4476_/Y vssd1 vssd1 vccd1 vccd1 _5071_/D sky130_fd_sc_hd__o211a_1
X_3428_ _5223_/Q vssd1 vssd1 vccd1 vccd1 _3873_/B sky130_fd_sc_hd__inv_2
X_3359_ _3359_/A _3359_/B vssd1 vssd1 vccd1 vccd1 _3360_/B sky130_fd_sc_hd__nand2_1
X_5029_ _5301_/CLK _5029_/D vssd1 vssd1 vccd1 vccd1 _5029_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2730_ _4661_/A _5298_/Q vssd1 vssd1 vccd1 vccd1 _2731_/B sky130_fd_sc_hd__nand2_1
X_2661_ _2661_/A _2661_/B _2660_/Y vssd1 vssd1 vccd1 vccd1 _2814_/A sky130_fd_sc_hd__or3b_4
X_4400_ _5112_/Q _4739_/B _4429_/B _4423_/D vssd1 vssd1 vccd1 vccd1 _4416_/A sky130_fd_sc_hd__o22ai_4
X_2592_ _2602_/A _4835_/A vssd1 vssd1 vccd1 vccd1 _2592_/Y sky130_fd_sc_hd__nand2_1
X_4331_ _4331_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4332_/B sky130_fd_sc_hd__nor2_1
X_4262_ _4468_/A vssd1 vssd1 vccd1 vccd1 _4457_/A sky130_fd_sc_hd__inv_2
X_3213_ _3213_/A vssd1 vssd1 vccd1 vccd1 _3213_/Y sky130_fd_sc_hd__inv_2
X_4193_ _4190_/Y _4310_/A _4192_/X vssd1 vssd1 vccd1 vccd1 _5091_/D sky130_fd_sc_hd__a21oi_1
XFILLER_39_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3144_ _3274_/A _3271_/A vssd1 vssd1 vccd1 vccd1 _3145_/C sky130_fd_sc_hd__nand2_1
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3075_ _5167_/Q _3765_/B vssd1 vssd1 vccd1 vccd1 _3108_/A sky130_fd_sc_hd__or2_1
XFILLER_27_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3977_ _4986_/Q _4986_/D vssd1 vssd1 vccd1 vccd1 _3981_/B sky130_fd_sc_hd__and2b_1
X_2928_ _2927_/B _2927_/A _2848_/X vssd1 vssd1 vccd1 vccd1 _2928_/X sky130_fd_sc_hd__a21o_1
X_2859_ _2995_/A _3719_/B vssd1 vssd1 vccd1 vccd1 _2859_/Y sky130_fd_sc_hd__nand2_1
X_4529_ _4434_/X _4526_/Y _4527_/X _2915_/X _4528_/Y vssd1 vssd1 vccd1 vccd1 _5062_/D
+ sky130_fd_sc_hd__o311a_1
XFILLER_77_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput9 input9/A vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_1
XFILLER_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3900_ _4440_/A vssd1 vssd1 vccd1 vccd1 _3916_/A sky130_fd_sc_hd__clkbuf_2
X_4880_ _4880_/A vssd1 vssd1 vccd1 vccd1 _4882_/A sky130_fd_sc_hd__inv_2
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3831_ _3833_/A _3831_/B vssd1 vssd1 vccd1 vccd1 _3831_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3762_ _3762_/A vssd1 vssd1 vccd1 vccd1 _3762_/X sky130_fd_sc_hd__clkbuf_2
X_2713_ _2973_/A vssd1 vssd1 vccd1 vccd1 _2715_/A sky130_fd_sc_hd__inv_2
X_3693_ _3693_/A _3700_/B vssd1 vssd1 vccd1 vccd1 _3693_/X sky130_fd_sc_hd__and2_1
X_2644_ _5315_/Q _4725_/A vssd1 vssd1 vccd1 vccd1 _2834_/A sky130_fd_sc_hd__nor2_2
X_2575_ _5302_/Q _2567_/X _2563_/X _2574_/Y vssd1 vssd1 vccd1 vccd1 _5302_/D sky130_fd_sc_hd__o211a_1
X_4314_ _5060_/Q vssd1 vssd1 vccd1 vccd1 _4652_/B sky130_fd_sc_hd__inv_2
XFILLER_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5294_ _5301_/CLK _5294_/D vssd1 vssd1 vccd1 vccd1 _5294_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4245_ _5106_/Q _5074_/Q vssd1 vssd1 vccd1 vccd1 _4254_/A sky130_fd_sc_hd__nor2_1
X_4176_ _4174_/Y _4331_/A _4175_/Y vssd1 vssd1 vccd1 vccd1 _5096_/D sky130_fd_sc_hd__a21oi_1
XFILLER_67_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3127_ _3288_/A _3288_/B _3126_/X vssd1 vssd1 vccd1 vccd1 _3278_/B sky130_fd_sc_hd__a21oi_1
XFILLER_55_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3058_ _5271_/Q vssd1 vssd1 vccd1 vccd1 _3745_/B sky130_fd_sc_hd__inv_2
XPHY_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_73_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_69_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4030_ _4030_/A _4031_/D vssd1 vssd1 vccd1 vccd1 _4030_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4932_ _4932_/A vssd1 vssd1 vccd1 vccd1 _4966_/B sky130_fd_sc_hd__inv_2
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_44_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5196_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_45_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4863_ _4863_/A _4872_/B vssd1 vssd1 vccd1 vccd1 _4863_/Y sky130_fd_sc_hd__nand2_1
X_4794_ _4794_/A _4794_/B vssd1 vssd1 vccd1 vccd1 _4794_/Y sky130_fd_sc_hd__nor2_1
X_3814_ _5150_/Q _3809_/X _3804_/X _3813_/Y vssd1 vssd1 vccd1 vccd1 _5150_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3745_ _3752_/A _3745_/B vssd1 vssd1 vccd1 vccd1 _3745_/Y sky130_fd_sc_hd__nand2_1
X_3676_ _3677_/A _3677_/B _3679_/A _2897_/X vssd1 vssd1 vccd1 vccd1 _3676_/X sky130_fd_sc_hd__a31o_1
X_2627_ _3755_/A vssd1 vssd1 vccd1 vccd1 _3713_/A sky130_fd_sc_hd__clkbuf_2
X_2558_ _5306_/Q _2548_/X _2544_/X _2557_/Y vssd1 vssd1 vccd1 vccd1 _5306_/D sky130_fd_sc_hd__o211a_1
X_5277_ _5277_/CLK _5277_/D vssd1 vssd1 vccd1 vccd1 _5277_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4228_ _4226_/Y _4221_/B _4588_/A vssd1 vssd1 vccd1 vccd1 _4228_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4159_ _5099_/Q _4111_/X _4112_/X _4094_/X _5100_/Q vssd1 vssd1 vccd1 vccd1 _4160_/B
+ sky130_fd_sc_hd__a41oi_1
XFILLER_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_35_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5228_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_26_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 _5268_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_14_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput12 hold12/X vssd1 vssd1 vccd1 vccd1 hold11/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput23 rst vssd1 vssd1 vccd1 vccd1 hold44/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3530_ _3371_/Y _3541_/B _3531_/B _3531_/C vssd1 vssd1 vccd1 vccd1 _3530_/Y sky130_fd_sc_hd__o2bb2ai_1
XFILLER_6_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3461_ _3640_/B _3461_/B vssd1 vssd1 vccd1 vccd1 _3647_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3392_ _3381_/Y _3386_/X _3390_/Y _3390_/A _3391_/Y vssd1 vssd1 vccd1 vccd1 _3551_/A
+ sky130_fd_sc_hd__a311o_2
X_5200_ _5204_/CLK _5200_/D vssd1 vssd1 vccd1 vccd1 _5200_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5131_ _5197_/CLK _5131_/D vssd1 vssd1 vccd1 vccd1 _5131_/Q sky130_fd_sc_hd__dfxtp_1
X_5062_ _5062_/CLK _5062_/D vssd1 vssd1 vccd1 vccd1 _5062_/Q sky130_fd_sc_hd__dfxtp_1
X_4013_ _4037_/C _4036_/B _4015_/B vssd1 vssd1 vccd1 vccd1 _4022_/C sky130_fd_sc_hd__nand3_4
XFILLER_84_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_17_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5027_/CLK sky130_fd_sc_hd__clkbuf_16
X_4915_ _4958_/B _5012_/Q _4940_/A _5008_/Q _4914_/X vssd1 vssd1 vccd1 vccd1 _4920_/A
+ sky130_fd_sc_hd__o221a_1
X_4846_ _4846_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4846_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4777_ _5042_/Q _4770_/X _4775_/Y _4776_/X _4584_/X vssd1 vssd1 vccd1 vccd1 _5042_/D
+ sky130_fd_sc_hd__o221a_1
X_3728_ _3754_/A vssd1 vssd1 vccd1 vccd1 _3728_/X sky130_fd_sc_hd__buf_1
X_3659_ _3653_/X _3658_/Y _3615_/X vssd1 vssd1 vccd1 vccd1 _3659_/X sky130_fd_sc_hd__a21o_1
XFILLER_57_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2961_ _3646_/A vssd1 vssd1 vccd1 vccd1 _2961_/X sky130_fd_sc_hd__clkbuf_2
X_4700_ _4700_/A vssd1 vssd1 vccd1 vccd1 _4762_/B sky130_fd_sc_hd__inv_2
X_4631_ _4631_/A _4634_/B vssd1 vssd1 vccd1 vccd1 _4875_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2892_ _2892_/A vssd1 vssd1 vccd1 vccd1 _2892_/X sky130_fd_sc_hd__buf_2
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4562_ _4561_/B _4561_/A _4484_/X vssd1 vssd1 vccd1 vccd1 _4562_/X sky130_fd_sc_hd__a21o_1
X_3513_ _3512_/Y _3494_/A _3508_/B vssd1 vssd1 vccd1 vccd1 _3513_/X sky130_fd_sc_hd__a21o_1
X_4493_ _4499_/B _4499_/A vssd1 vssd1 vccd1 vccd1 _4496_/A sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_6_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5062_/CLK sky130_fd_sc_hd__clkbuf_16
X_3444_ _5132_/Q _3860_/B vssd1 vssd1 vccd1 vccd1 _3663_/B sky130_fd_sc_hd__or2_1
XFILLER_69_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3375_ _5155_/Q _3800_/B vssd1 vssd1 vccd1 vccd1 _3544_/A sky130_fd_sc_hd__nor2_2
XFILLER_69_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5114_ _5114_/CLK _5114_/D vssd1 vssd1 vccd1 vccd1 _5114_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5045_ _5317_/CLK _5045_/D vssd1 vssd1 vccd1 vccd1 _5045_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_72_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_65_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4829_ _5031_/Q _4217_/X _4807_/X _4828_/X vssd1 vssd1 vccd1 vccd1 _5031_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_84_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3160_ _3167_/A vssd1 vssd1 vccd1 vccd1 _3243_/B sky130_fd_sc_hd__inv_2
Xhold1 hold1/A vssd1 vssd1 vccd1 vccd1 hold1/X sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _3781_/B _5162_/Q vssd1 vssd1 vccd1 vccd1 _3092_/B sky130_fd_sc_hd__nand2_1
XFILLER_81_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3993_ _3993_/A _4031_/D vssd1 vssd1 vccd1 vccd1 _3994_/A sky130_fd_sc_hd__nand2_1
XFILLER_13_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2944_ _2949_/B vssd1 vssd1 vccd1 vccd1 _2950_/B sky130_fd_sc_hd__inv_2
X_2875_ _2875_/A _2875_/B vssd1 vssd1 vccd1 vccd1 _2875_/Y sky130_fd_sc_hd__nor2_1
X_4614_ _4671_/A _4611_/Y _4671_/B vssd1 vssd1 vccd1 vccd1 _4790_/A sky130_fd_sc_hd__o21bai_1
X_4545_ _4545_/A vssd1 vssd1 vccd1 vccd1 _4553_/B sky130_fd_sc_hd__inv_2
X_4476_ _4468_/B _4474_/X _4475_/X vssd1 vssd1 vccd1 vccd1 _4476_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_89_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3427_ _5128_/Q _3871_/B vssd1 vssd1 vccd1 vccd1 _3691_/A sky130_fd_sc_hd__nor2_4
XFILLER_85_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3358_ _3789_/B _5159_/Q vssd1 vssd1 vccd1 vccd1 _3359_/A sky130_fd_sc_hd__nand2_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3289_ _3295_/B _3295_/A vssd1 vssd1 vccd1 vccd1 _3289_/X sky130_fd_sc_hd__or2_1
X_5028_ _5062_/CLK _5028_/D vssd1 vssd1 vccd1 vccd1 _5028_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2660_ _2776_/A _2865_/B vssd1 vssd1 vccd1 vccd1 _2660_/Y sky130_fd_sc_hd__nand2_1
X_2591_ _5030_/Q vssd1 vssd1 vccd1 vccd1 _4835_/A sky130_fd_sc_hd__inv_2
XFILLER_5_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4330_ _5064_/Q vssd1 vssd1 vccd1 vccd1 _4666_/B sky130_fd_sc_hd__inv_2
XFILLER_4_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4261_ _4365_/A _4602_/B vssd1 vssd1 vccd1 vccd1 _4468_/A sky130_fd_sc_hd__nor2_1
XFILLER_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3212_ _3212_/A _3212_/B vssd1 vssd1 vccd1 vccd1 _3213_/A sky130_fd_sc_hd__nor2_1
X_4192_ _4111_/X _4112_/X _4180_/C _4214_/A vssd1 vssd1 vccd1 vccd1 _4192_/X sky130_fd_sc_hd__a31o_1
XFILLER_39_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3143_ _3143_/A _3143_/B vssd1 vssd1 vccd1 vccd1 _3271_/A sky130_fd_sc_hd__nor2_2
X_3074_ _3771_/B _5166_/Q _3108_/B vssd1 vssd1 vccd1 vccd1 _3076_/A sky130_fd_sc_hd__or3b_2
XFILLER_35_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3976_ _4986_/D _4986_/Q vssd1 vssd1 vccd1 vccd1 _3981_/A sky130_fd_sc_hd__and2b_1
X_2927_ _2927_/A _2927_/B vssd1 vssd1 vccd1 vccd1 _2927_/Y sky130_fd_sc_hd__nor2_1
X_2858_ _5281_/Q vssd1 vssd1 vccd1 vccd1 _3719_/B sky130_fd_sc_hd__inv_2
X_2789_ _5316_/Q _4591_/A vssd1 vssd1 vccd1 vccd1 _2793_/A sky130_fd_sc_hd__nor2_1
X_4528_ _4528_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4528_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4459_ _4468_/B _4470_/B _4265_/B vssd1 vssd1 vccd1 vccd1 _4460_/B sky130_fd_sc_hd__a21oi_1
XFILLER_73_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3830_ _3830_/A vssd1 vssd1 vccd1 vccd1 _3830_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_20_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3761_ _5169_/Q _3754_/X _3749_/X _3760_/Y vssd1 vssd1 vccd1 vccd1 _5169_/D sky130_fd_sc_hd__o211a_1
X_2712_ _2712_/A _2712_/B vssd1 vssd1 vccd1 vccd1 _2973_/A sky130_fd_sc_hd__nand2_2
XFILLER_72_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3692_ _3691_/Y _3700_/B _3693_/A _2897_/X vssd1 vssd1 vccd1 vccd1 _3692_/X sky130_fd_sc_hd__a31o_1
X_2643_ _5286_/Q _2625_/X _2619_/X _2642_/Y vssd1 vssd1 vccd1 vccd1 _5286_/D sky130_fd_sc_hd__o211a_1
X_2574_ _2584_/A _4808_/A vssd1 vssd1 vccd1 vccd1 _2574_/Y sky130_fd_sc_hd__nand2_1
X_4313_ _5092_/Q _5060_/Q vssd1 vssd1 vccd1 vccd1 _4316_/A sky130_fd_sc_hd__nor2_1
X_5293_ _5301_/CLK _5293_/D vssd1 vssd1 vccd1 vccd1 _5293_/Q sky130_fd_sc_hd__dfxtp_1
X_4244_ _4244_/A _4592_/B vssd1 vssd1 vccd1 vccd1 _4429_/B sky130_fd_sc_hd__nor2_4
X_4175_ _4168_/B _4183_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4175_/Y sky130_fd_sc_hd__o21ai_1
X_3126_ _3287_/A _3287_/B _3295_/B vssd1 vssd1 vccd1 vccd1 _3126_/X sky130_fd_sc_hd__or3_1
XFILLER_55_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3057_ _3266_/B _3145_/B vssd1 vssd1 vccd1 vccd1 _3057_/Y sky130_fd_sc_hd__nor2_1
XPHY_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3959_ _5104_/Q vssd1 vssd1 vccd1 vccd1 _4258_/A sky130_fd_sc_hd__inv_2
XFILLER_18_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4931_ _4931_/A _4931_/B vssd1 vssd1 vccd1 vccd1 _4934_/B sky130_fd_sc_hd__nor2_1
X_4862_ _4862_/A _4862_/B _4862_/C vssd1 vssd1 vccd1 vccd1 _4862_/X sky130_fd_sc_hd__and3_1
X_3813_ _3820_/A _3813_/B vssd1 vssd1 vccd1 vccd1 _3813_/Y sky130_fd_sc_hd__nand2_1
X_4793_ _4691_/A _4691_/B _4792_/Y vssd1 vssd1 vccd1 vccd1 _4794_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3744_ _5176_/Q _3741_/X _3736_/X _3743_/Y vssd1 vssd1 vccd1 vccd1 _5176_/D sky130_fd_sc_hd__o211a_1
X_3675_ _3675_/A _3675_/B vssd1 vssd1 vccd1 vccd1 _3679_/A sky130_fd_sc_hd__nor2_1
X_2626_ _3769_/A vssd1 vssd1 vccd1 vccd1 _3755_/A sky130_fd_sc_hd__buf_2
X_2557_ _2565_/A _4788_/A vssd1 vssd1 vccd1 vccd1 _2557_/Y sky130_fd_sc_hd__nand2_1
X_5276_ _5280_/CLK _5276_/D vssd1 vssd1 vccd1 vccd1 _5276_/Q sky130_fd_sc_hd__dfxtp_1
X_4227_ _4764_/A vssd1 vssd1 vccd1 vccd1 _4588_/A sky130_fd_sc_hd__clkbuf_4
X_4158_ _5101_/Q _4160_/C _4157_/Y vssd1 vssd1 vccd1 vccd1 _5101_/D sky130_fd_sc_hd__o21a_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4089_ _4156_/C vssd1 vssd1 vccd1 vccd1 _4119_/C sky130_fd_sc_hd__buf_2
X_3109_ _3318_/B _3309_/A vssd1 vssd1 vccd1 vccd1 _3109_/X sky130_fd_sc_hd__or2_1
XFILLER_43_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput13 phase_in[10] vssd1 vssd1 vccd1 vccd1 hold42/A sky130_fd_sc_hd__buf_1
X_3460_ _3851_/B _5136_/Q vssd1 vssd1 vccd1 vccd1 _3461_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3391_ _3391_/A _3391_/B vssd1 vssd1 vccd1 vccd1 _3391_/Y sky130_fd_sc_hd__nor2_1
X_5130_ _5196_/CLK _5130_/D vssd1 vssd1 vccd1 vccd1 _5130_/Q sky130_fd_sc_hd__dfxtp_1
X_5061_ _5062_/CLK _5061_/D vssd1 vssd1 vccd1 vccd1 _5061_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4012_ _4029_/A _4029_/B vssd1 vssd1 vccd1 vccd1 _4015_/B sky130_fd_sc_hd__nor2_2
XFILLER_84_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4914_ _5122_/Q _3923_/Y _5117_/Q _3927_/Y vssd1 vssd1 vccd1 vccd1 _4914_/X sky130_fd_sc_hd__o22a_1
XFILLER_52_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4845_ _4845_/A _4845_/B vssd1 vssd1 vccd1 vccd1 _4845_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4776_ _4775_/B _4775_/A _4764_/X vssd1 vssd1 vccd1 vccd1 _4776_/X sky130_fd_sc_hd__a21o_1
XFILLER_20_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3727_ _5182_/Q _3715_/X _3723_/X _3726_/Y vssd1 vssd1 vccd1 vccd1 _5182_/D sky130_fd_sc_hd__o211a_1
X_3658_ _3658_/A _3658_/B vssd1 vssd1 vccd1 vccd1 _3658_/Y sky130_fd_sc_hd__nand2_1
X_2609_ _5025_/Q vssd1 vssd1 vccd1 vccd1 _4643_/A sky130_fd_sc_hd__inv_2
X_3589_ _3578_/Y _3494_/A _3508_/Y vssd1 vssd1 vccd1 vccd1 _3589_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5259_ _5288_/CLK _5259_/D vssd1 vssd1 vccd1 vccd1 _5259_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2960_ _3843_/A vssd1 vssd1 vccd1 vccd1 _3646_/A sky130_fd_sc_hd__clkbuf_2
X_2891_ _2886_/Y _2887_/X _2890_/X vssd1 vssd1 vccd1 vccd1 _5277_/D sky130_fd_sc_hd__o21a_1
XPHY_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4630_ _4630_/A _4862_/C vssd1 vssd1 vccd1 vccd1 _4865_/A sky130_fd_sc_hd__and2_1
XFILLER_30_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4561_ _4561_/A _4561_/B vssd1 vssd1 vccd1 vccd1 _4561_/Y sky130_fd_sc_hd__nor2_1
X_3512_ _3512_/A vssd1 vssd1 vccd1 vccd1 _3512_/Y sky130_fd_sc_hd__inv_2
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4492_ _4780_/B vssd1 vssd1 vccd1 vccd1 _4492_/X sky130_fd_sc_hd__clkbuf_2
X_3443_ _5228_/Q vssd1 vssd1 vccd1 vccd1 _3860_/B sky130_fd_sc_hd__inv_2
XFILLER_69_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5113_ _5114_/CLK _5113_/D vssd1 vssd1 vccd1 vccd1 _5113_/Q sky130_fd_sc_hd__dfxtp_1
X_3374_ _5251_/Q vssd1 vssd1 vccd1 vccd1 _3800_/B sky130_fd_sc_hd__inv_2
XFILLER_57_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5044_ _5317_/CLK _5044_/D vssd1 vssd1 vccd1 vccd1 _5044_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_27_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4828_ _4827_/X _4823_/A _4542_/X vssd1 vssd1 vccd1 vccd1 _4828_/X sky130_fd_sc_hd__a21o_1
X_4759_ _4799_/A _5045_/Q vssd1 vssd1 vccd1 vccd1 _4759_/Y sky130_fd_sc_hd__nand2_1
XFILLER_88_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_88_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold2 phase_in[1] vssd1 vssd1 vccd1 vccd1 hold2/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3090_ _3090_/A vssd1 vssd1 vccd1 vccd1 _3345_/A sky130_fd_sc_hd__inv_2
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3992_ _4031_/C _3993_/A _4031_/D vssd1 vssd1 vccd1 vccd1 _4032_/A sky130_fd_sc_hd__nand3b_4
X_2943_ _2943_/A _2943_/B vssd1 vssd1 vccd1 vccd1 _2949_/B sky130_fd_sc_hd__nand2_1
X_2874_ _2874_/A _2874_/B vssd1 vssd1 vccd1 vccd1 _2875_/B sky130_fd_sc_hd__and2_1
X_4613_ _4815_/A _4613_/B vssd1 vssd1 vccd1 vccd1 _4671_/B sky130_fd_sc_hd__nor2_1
X_4544_ _4530_/X _5059_/Q _4540_/X _4543_/X vssd1 vssd1 vccd1 vccd1 _5059_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4475_ _4770_/A vssd1 vssd1 vccd1 vccd1 _4475_/X sky130_fd_sc_hd__buf_2
X_3426_ _5224_/Q vssd1 vssd1 vccd1 vccd1 _3871_/B sky130_fd_sc_hd__inv_2
X_3357_ _3792_/B _5158_/Q vssd1 vssd1 vccd1 vccd1 _3367_/B sky130_fd_sc_hd__nand2_1
XFILLER_85_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5027_ _5027_/CLK _5027_/D vssd1 vssd1 vccd1 vccd1 _5027_/Q sky130_fd_sc_hd__dfxtp_1
X_3288_ _3288_/A _3288_/B vssd1 vssd1 vccd1 vccd1 _3295_/A sky130_fd_sc_hd__and2_1
XFILLER_38_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_70_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2590_ _5298_/Q _2586_/X _2582_/X _2589_/Y vssd1 vssd1 vccd1 vccd1 _5298_/D sky130_fd_sc_hd__o211a_1
XFILLER_5_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4260_ _5071_/Q vssd1 vssd1 vccd1 vccd1 _4602_/B sky130_fd_sc_hd__inv_2
X_4191_ _5091_/Q vssd1 vssd1 vccd1 vccd1 _4310_/A sky130_fd_sc_hd__inv_2
X_3211_ _5282_/Q _3211_/B vssd1 vssd1 vccd1 vccd1 _3212_/B sky130_fd_sc_hd__nor2_1
XFILLER_79_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3142_ _3142_/A _3142_/B vssd1 vssd1 vccd1 vccd1 _3274_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073_ _3765_/B _5167_/Q vssd1 vssd1 vccd1 vccd1 _3108_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3975_ _4982_/Q _4982_/D vssd1 vssd1 vccd1 vccd1 _4039_/B sky130_fd_sc_hd__xor2_4
XFILLER_50_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2926_ _2926_/A _2926_/B vssd1 vssd1 vccd1 vccd1 _2927_/B sky130_fd_sc_hd__nand2_1
X_2857_ _2867_/C _2857_/B _2857_/C vssd1 vssd1 vccd1 vccd1 _2857_/X sky130_fd_sc_hd__and3_1
X_2788_ _2834_/A _2784_/Y _2787_/Y vssd1 vssd1 vccd1 vccd1 _2827_/A sky130_fd_sc_hd__o21ai_1
X_4527_ _4527_/A _4527_/B _4527_/C vssd1 vssd1 vccd1 vccd1 _4527_/X sky130_fd_sc_hd__and3_1
X_4458_ _4474_/A _4474_/B _4474_/C vssd1 vssd1 vccd1 vccd1 _4468_/B sky130_fd_sc_hd__a21oi_2
XFILLER_49_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3409_ _5234_/Q vssd1 vssd1 vccd1 vccd1 _3845_/B sky130_fd_sc_hd__inv_2
X_4389_ _4444_/B _4396_/C vssd1 vssd1 vccd1 vccd1 _4390_/B sky130_fd_sc_hd__nor2_1
XFILLER_85_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3760_ _3765_/A _3760_/B vssd1 vssd1 vccd1 vccd1 _3760_/Y sky130_fd_sc_hd__nand2_1
XFILLER_32_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2711_ _4846_/A _5294_/Q vssd1 vssd1 vccd1 vccd1 _2712_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3691_ _3691_/A _3691_/B vssd1 vssd1 vccd1 vccd1 _3691_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2642_ _3713_/A _3022_/B vssd1 vssd1 vccd1 vccd1 _2642_/Y sky130_fd_sc_hd__nand2_1
X_2573_ _4683_/A vssd1 vssd1 vccd1 vccd1 _4808_/A sky130_fd_sc_hd__buf_1
X_5292_ _5292_/CLK _5292_/D vssd1 vssd1 vccd1 vccd1 _5292_/Q sky130_fd_sc_hd__dfxtp_1
X_4312_ _4312_/A _4536_/B vssd1 vssd1 vccd1 vccd1 _4541_/B sky130_fd_sc_hd__nand2_1
X_4243_ _5079_/Q vssd1 vssd1 vccd1 vccd1 _4592_/B sky130_fd_sc_hd__inv_2
X_4174_ _4174_/A _5095_/Q vssd1 vssd1 vccd1 vccd1 _4174_/Y sky130_fd_sc_hd__nand2_1
XFILLER_82_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3125_ _3125_/A _3125_/B vssd1 vssd1 vccd1 vccd1 _3295_/B sky130_fd_sc_hd__or2_1
XFILLER_82_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3056_ _3056_/A vssd1 vssd1 vccd1 vccd1 _3145_/B sky130_fd_sc_hd__inv_2
XFILLER_82_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3958_ _4149_/B _5106_/Q _5105_/Q vssd1 vssd1 vccd1 vccd1 _3962_/A sky130_fd_sc_hd__and3_1
X_3889_ _4440_/A vssd1 vssd1 vccd1 vccd1 _4572_/A sky130_fd_sc_hd__clkbuf_2
X_2909_ _2927_/A _2930_/B _2930_/A vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__or3_1
XFILLER_76_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4930_ _4930_/A _4930_/B vssd1 vssd1 vccd1 vccd1 _4931_/B sky130_fd_sc_hd__nor2_1
XFILLER_64_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4861_ _4862_/A _4862_/C _4862_/B vssd1 vssd1 vccd1 vccd1 _4861_/Y sky130_fd_sc_hd__a21oi_1
X_3812_ _5151_/Q _3809_/X _3804_/X _3811_/Y vssd1 vssd1 vccd1 vccd1 _5151_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4792_ _4797_/B _4797_/A vssd1 vssd1 vccd1 vccd1 _4792_/Y sky130_fd_sc_hd__nand2_1
X_3743_ _3752_/A _3743_/B vssd1 vssd1 vccd1 vccd1 _3743_/Y sky130_fd_sc_hd__nand2_1
X_3674_ _5131_/Q _3864_/B vssd1 vssd1 vccd1 vccd1 _3675_/B sky130_fd_sc_hd__nor2_1
X_2625_ _3613_/A vssd1 vssd1 vccd1 vccd1 _2625_/X sky130_fd_sc_hd__clkbuf_2
X_2556_ _5039_/Q vssd1 vssd1 vccd1 vccd1 _4788_/A sky130_fd_sc_hd__inv_2
X_5275_ _5277_/CLK _5275_/D vssd1 vssd1 vccd1 vccd1 _5275_/Q sky130_fd_sc_hd__dfxtp_1
X_4226_ _4226_/A _4226_/B vssd1 vssd1 vccd1 vccd1 _4226_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4157_ _4169_/B _4152_/X _4169_/A vssd1 vssd1 vccd1 vccd1 _4157_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_28_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108_ _3108_/A _3108_/B vssd1 vssd1 vccd1 vccd1 _3309_/A sky130_fd_sc_hd__nand2_1
XFILLER_28_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4088_ _4180_/A _4180_/B _4105_/A vssd1 vssd1 vccd1 vccd1 _4156_/C sky130_fd_sc_hd__nand3_4
X_3039_ _3034_/Y _3174_/A _3175_/B vssd1 vssd1 vccd1 vccd1 _3223_/B sky130_fd_sc_hd__a21oi_4
XFILLER_36_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput14 hold2/X vssd1 vssd1 vccd1 vccd1 hold1/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3390_ _3390_/A _3391_/A vssd1 vssd1 vccd1 vccd1 _3390_/Y sky130_fd_sc_hd__nor2_2
X_5060_ _5118_/CLK _5060_/D vssd1 vssd1 vccd1 vccd1 _5060_/Q sky130_fd_sc_hd__dfxtp_1
X_4011_ _4011_/A _4030_/A _4011_/C vssd1 vssd1 vccd1 vccd1 _4036_/B sky130_fd_sc_hd__nand3_4
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4913_ _4913_/A _4913_/B vssd1 vssd1 vccd1 vccd1 _5003_/D sky130_fd_sc_hd__nor2_1
XFILLER_33_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4844_ _5028_/Q _4475_/X _4842_/Y _4843_/X _4785_/X vssd1 vssd1 vccd1 vccd1 _5028_/D
+ sky130_fd_sc_hd__o221a_1
X_4775_ _4775_/A _4775_/B vssd1 vssd1 vccd1 vccd1 _4775_/Y sky130_fd_sc_hd__nor2_1
X_3726_ _3726_/A _3726_/B vssd1 vssd1 vccd1 vccd1 _3726_/Y sky130_fd_sc_hd__nand2_1
X_3657_ _5199_/Q _3650_/X _3655_/Y _3656_/X _3644_/X vssd1 vssd1 vccd1 vccd1 _5199_/D
+ sky130_fd_sc_hd__o221a_1
X_2608_ _5293_/Q _2604_/X _2600_/X _2607_/Y vssd1 vssd1 vccd1 vccd1 _5293_/D sky130_fd_sc_hd__o211a_1
X_3588_ _5212_/Q _3328_/X _3585_/X _3587_/X vssd1 vssd1 vccd1 vccd1 _5212_/D sky130_fd_sc_hd__o211a_1
X_2539_ _5311_/Q _2528_/X _2522_/X _2538_/Y vssd1 vssd1 vccd1 vccd1 _5311_/D sky130_fd_sc_hd__o211a_1
XFILLER_0_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5258_ _5267_/CLK _5258_/D vssd1 vssd1 vccd1 vccd1 _5258_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5189_ _5285_/CLK _5189_/D vssd1 vssd1 vccd1 vccd1 _5189_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4209_ _4417_/A vssd1 vssd1 vccd1 vccd1 _4770_/A sky130_fd_sc_hd__buf_1
XFILLER_56_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2890_ _5277_/Q _2888_/X _2889_/X vssd1 vssd1 vccd1 vccd1 _2890_/X sky130_fd_sc_hd__o21a_1
XPHY_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4560_ _5087_/Q _5055_/Q _4559_/X vssd1 vssd1 vccd1 vccd1 _4561_/B sky130_fd_sc_hd__a21o_1
XFILLER_8_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3511_ _3511_/A _3511_/B vssd1 vssd1 vccd1 vccd1 _3511_/Y sky130_fd_sc_hd__nor2_1
X_4491_ _4488_/X _4490_/Y _4214_/X vssd1 vssd1 vccd1 vccd1 _5069_/D sky130_fd_sc_hd__a21oi_1
X_3442_ _3675_/A vssd1 vssd1 vccd1 vccd1 _3442_/Y sky130_fd_sc_hd__inv_2
X_3373_ _5252_/Q _5156_/Q vssd1 vssd1 vccd1 vccd1 _3539_/A sky130_fd_sc_hd__nor2_2
X_5112_ _5112_/CLK _5112_/D vssd1 vssd1 vccd1 vccd1 _5112_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5043_ _5311_/CLK _5043_/D vssd1 vssd1 vccd1 vccd1 _5043_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4827_ _4827_/A _4827_/B vssd1 vssd1 vccd1 vccd1 _4827_/X sky130_fd_sc_hd__or2_1
X_4758_ _4798_/A _4758_/B _4758_/C vssd1 vssd1 vccd1 vccd1 _4758_/X sky130_fd_sc_hd__or3_1
XFILLER_4_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3709_ _3843_/A vssd1 vssd1 vccd1 vccd1 _3762_/A sky130_fd_sc_hd__clkbuf_2
X_4689_ _4790_/A _4790_/B _4688_/X vssd1 vssd1 vccd1 vccd1 _4771_/A sky130_fd_sc_hd__o21bai_1
XFILLER_0_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold3 hold3/A vssd1 vssd1 vccd1 vccd1 hold3/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3991_ _3990_/A _3990_/B _3990_/C vssd1 vssd1 vccd1 vccd1 _4031_/D sky130_fd_sc_hd__o21ai_4
XFILLER_74_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2942_ _5268_/Q _2939_/X _2892_/X _2941_/X vssd1 vssd1 vccd1 vccd1 _5268_/D sky130_fd_sc_hd__o211a_1
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2873_ _2874_/A _2875_/A _2874_/B _2901_/A vssd1 vssd1 vccd1 vccd1 _2873_/X sky130_fd_sc_hd__a31o_1
X_4612_ _5066_/Q vssd1 vssd1 vccd1 vccd1 _4613_/B sky130_fd_sc_hd__inv_2
X_4543_ _4536_/A _4541_/Y _4542_/X vssd1 vssd1 vccd1 vccd1 _4543_/X sky130_fd_sc_hd__a21o_1
XFILLER_89_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4474_ _4474_/A _4474_/B _4474_/C vssd1 vssd1 vccd1 vccd1 _4474_/X sky130_fd_sc_hd__and3_1
X_3425_ _5129_/Q vssd1 vssd1 vccd1 vccd1 _3425_/Y sky130_fd_sc_hd__inv_2
X_3356_ _5254_/Q vssd1 vssd1 vccd1 vccd1 _3792_/B sky130_fd_sc_hd__inv_2
XFILLER_57_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3287_ _3287_/A _3287_/B vssd1 vssd1 vccd1 vccd1 _3291_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5026_ _5085_/CLK _5026_/D vssd1 vssd1 vccd1 vccd1 _5026_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3210_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3210_/X sky130_fd_sc_hd__clkbuf_2
X_4190_ _4194_/A _4190_/B vssd1 vssd1 vccd1 vccd1 _4190_/Y sky130_fd_sc_hd__nand2_1
XFILLER_79_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3141_ _3141_/A vssd1 vssd1 vccd1 vccd1 _3142_/B sky130_fd_sc_hd__inv_2
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3072_ _5263_/Q vssd1 vssd1 vccd1 vccd1 _3765_/B sky130_fd_sc_hd__inv_2
XFILLER_90_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3974_ _3974_/A _4992_/D vssd1 vssd1 vccd1 vccd1 _4016_/A sky130_fd_sc_hd__nand2_2
X_2925_ _2930_/B _2930_/A vssd1 vssd1 vccd1 vccd1 _2926_/A sky130_fd_sc_hd__or2_1
XFILLER_50_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2856_ _2867_/C _2857_/C _2857_/B vssd1 vssd1 vccd1 vccd1 _2856_/Y sky130_fd_sc_hd__a21oi_1
X_2787_ _2787_/A _2787_/B vssd1 vssd1 vccd1 vccd1 _2787_/Y sky130_fd_sc_hd__nand2_1
X_4526_ _4527_/A _4527_/C _4527_/B vssd1 vssd1 vccd1 vccd1 _4526_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_2_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4457_ _4457_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4474_/C sky130_fd_sc_hd__nand2_1
XFILLER_49_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3408_ _3489_/A _3603_/B _3608_/B _3405_/Y _3407_/Y vssd1 vssd1 vccd1 vccd1 _3408_/Y
+ sky130_fd_sc_hd__o41ai_4
X_4388_ _4388_/A vssd1 vssd1 vccd1 vccd1 _4396_/C sky130_fd_sc_hd__inv_2
X_3339_ _3339_/A _3339_/B vssd1 vssd1 vccd1 vccd1 _3339_/Y sky130_fd_sc_hd__nor2_1
XFILLER_65_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5009_ _5118_/CLK hold15/X vssd1 vssd1 vccd1 vccd1 _5009_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2710_ _2700_/A _5025_/Q _2966_/B _2802_/A vssd1 vssd1 vccd1 vccd1 _2710_/Y sky130_fd_sc_hd__a31oi_1
X_3690_ _3871_/B _5128_/Q vssd1 vssd1 vccd1 vccd1 _3691_/B sky130_fd_sc_hd__and2_1
X_2641_ _5019_/Q vssd1 vssd1 vccd1 vccd1 _3022_/B sky130_fd_sc_hd__inv_2
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2572_ _5035_/Q vssd1 vssd1 vccd1 vccd1 _4683_/A sky130_fd_sc_hd__inv_2
X_5291_ _5292_/CLK _5291_/D vssd1 vssd1 vccd1 vccd1 _5291_/Q sky130_fd_sc_hd__dfxtp_1
X_4311_ _5091_/Q _5059_/Q vssd1 vssd1 vccd1 vccd1 _4536_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4242_ _5080_/Q vssd1 vssd1 vccd1 vccd1 _4739_/B sky130_fd_sc_hd__buf_2
XFILLER_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4173_ _4180_/A _4180_/B _4173_/C vssd1 vssd1 vccd1 vccd1 _4174_/A sky130_fd_sc_hd__and3_1
X_3124_ _3758_/B _5170_/Q vssd1 vssd1 vccd1 vccd1 _3125_/B sky130_fd_sc_hd__and2_1
XFILLER_27_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3055_ _3055_/A _3064_/A vssd1 vssd1 vccd1 vccd1 _3056_/A sky130_fd_sc_hd__nor2_2
XFILLER_70_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_47_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5114_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3957_ _4145_/B vssd1 vssd1 vccd1 vccd1 _4149_/B sky130_fd_sc_hd__inv_2
X_2908_ _2908_/A _2908_/B vssd1 vssd1 vccd1 vccd1 _2930_/A sky130_fd_sc_hd__nor2_1
X_3888_ _4893_/A vssd1 vssd1 vccd1 vccd1 _4440_/A sky130_fd_sc_hd__clkbuf_2
X_2839_ _2995_/A _3713_/B vssd1 vssd1 vccd1 vccd1 _2839_/Y sky130_fd_sc_hd__nand2_1
X_4509_ _4492_/X _5066_/Q _4505_/X _4507_/Y _4508_/X vssd1 vssd1 vccd1 vccd1 _5066_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_73_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_38_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5280_/CLK sky130_fd_sc_hd__clkbuf_16
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_29_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5252_/CLK sky130_fd_sc_hd__clkbuf_16
X_4860_ _4865_/B _4865_/A vssd1 vssd1 vccd1 vccd1 _4862_/A sky130_fd_sc_hd__nand2_1
XFILLER_60_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3811_ _3820_/A _3811_/B vssd1 vssd1 vccd1 vccd1 _3811_/Y sky130_fd_sc_hd__nand2_1
X_4791_ _4688_/B _4806_/B _4690_/Y vssd1 vssd1 vccd1 vccd1 _4797_/B sky130_fd_sc_hd__o21ai_1
X_3742_ _3755_/A vssd1 vssd1 vccd1 vccd1 _3752_/A sky130_fd_sc_hd__buf_1
XFILLER_9_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3673_ _3673_/A vssd1 vssd1 vccd1 vccd1 _3677_/A sky130_fd_sc_hd__inv_2
X_2624_ _3767_/A vssd1 vssd1 vccd1 vccd1 _3613_/A sky130_fd_sc_hd__clkbuf_2
X_2555_ _5307_/Q _2548_/X _2544_/X _2554_/Y vssd1 vssd1 vccd1 vccd1 _5307_/D sky130_fd_sc_hd__o211a_1
X_5274_ _5274_/CLK _5274_/D vssd1 vssd1 vccd1 vccd1 _5274_/Q sky130_fd_sc_hd__dfxtp_1
X_4225_ _4217_/X _5085_/Q _4223_/Y _4224_/X _3695_/X vssd1 vssd1 vccd1 vccd1 _5085_/D
+ sky130_fd_sc_hd__o221a_1
X_4156_ _4352_/A _4356_/A _4156_/C vssd1 vssd1 vccd1 vccd1 _4160_/C sky130_fd_sc_hd__nor3_4
XFILLER_55_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3107_ _5262_/Q _5166_/Q vssd1 vssd1 vccd1 vccd1 _3318_/B sky130_fd_sc_hd__xor2_2
XFILLER_43_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4087_ _4165_/A _4087_/B _4190_/B vssd1 vssd1 vccd1 vccd1 _4105_/A sky130_fd_sc_hd__and3_2
XFILLER_70_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3038_ _3724_/B _5183_/Q vssd1 vssd1 vccd1 vccd1 _3175_/B sky130_fd_sc_hd__and2_1
XFILLER_62_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4989_ _4990_/CLK hold41/X vssd1 vssd1 vccd1 vccd1 _4990_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_11_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 hold4/X vssd1 vssd1 vccd1 vccd1 hold3/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_4010_ _4030_/A _4011_/A _4008_/X _4009_/Y vssd1 vssd1 vccd1 vccd1 _4037_/C sky130_fd_sc_hd__o2bb2ai_4
XFILLER_37_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4912_ _4912_/A _4912_/B vssd1 vssd1 vccd1 vccd1 _4913_/B sky130_fd_sc_hd__nand2_1
XFILLER_18_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4843_ _4842_/B _4842_/A _3907_/A vssd1 vssd1 vccd1 vccd1 _4843_/X sky130_fd_sc_hd__a21o_1
XFILLER_33_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4774_ _4780_/A _4774_/B vssd1 vssd1 vccd1 vccd1 _4775_/B sky130_fd_sc_hd__nand2_1
XFILLER_20_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3725_ _5183_/Q _3715_/X _3723_/X _3724_/Y vssd1 vssd1 vccd1 vccd1 _5183_/D sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_9_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5118_/CLK sky130_fd_sc_hd__clkbuf_16
X_3656_ _3655_/B _3655_/A _3642_/X vssd1 vssd1 vccd1 vccd1 _3656_/X sky130_fd_sc_hd__a21o_1
X_2607_ _2622_/A _4853_/A vssd1 vssd1 vccd1 vccd1 _2607_/Y sky130_fd_sc_hd__nand2_1
X_3587_ _3582_/B _3586_/Y _3306_/X vssd1 vssd1 vccd1 vccd1 _3587_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2538_ _2546_/A _4704_/A vssd1 vssd1 vccd1 vccd1 _2538_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5257_ _5267_/CLK _5257_/D vssd1 vssd1 vccd1 vccd1 _5257_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_57_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4208_ _4208_/A _4208_/B _4222_/A _4208_/D vssd1 vssd1 vccd1 vccd1 _4208_/X sky130_fd_sc_hd__and4_1
XFILLER_87_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5188_ _5283_/CLK _5188_/D vssd1 vssd1 vccd1 vccd1 _5188_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4139_ _4139_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4139_/Y sky130_fd_sc_hd__nand2_1
XFILLER_71_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3510_ _3408_/Y _3490_/Y _3509_/X vssd1 vssd1 vccd1 vccd1 _3572_/A sky130_fd_sc_hd__o21bai_2
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4490_ _4799_/A _5069_/Q vssd1 vssd1 vccd1 vccd1 _4490_/Y sky130_fd_sc_hd__nand2_1
X_3441_ _5227_/Q _3441_/B vssd1 vssd1 vccd1 vccd1 _3675_/A sky130_fd_sc_hd__nor2_2
X_3372_ _5252_/Q _5156_/Q vssd1 vssd1 vccd1 vccd1 _3539_/B sky130_fd_sc_hd__and2_1
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5111_ _5114_/CLK _5111_/D vssd1 vssd1 vccd1 vccd1 _5111_/Q sky130_fd_sc_hd__dfxtp_2
X_5042_ _5076_/CLK _5042_/D vssd1 vssd1 vccd1 vccd1 _5042_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_65_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4826_ _5032_/Q _4770_/X _4824_/Y _4825_/X _4785_/X vssd1 vssd1 vccd1 vccd1 _5032_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_21_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4757_ _4757_/A _4757_/B vssd1 vssd1 vccd1 vccd1 _4758_/C sky130_fd_sc_hd__and2_1
X_3708_ _5189_/Q _3668_/X _3646_/X _3707_/Y vssd1 vssd1 vccd1 vccd1 _5189_/D sky130_fd_sc_hd__o211a_1
X_4688_ _4688_/A _4688_/B vssd1 vssd1 vccd1 vccd1 _4688_/X sky130_fd_sc_hd__or2_1
X_3639_ _3647_/B _3647_/A vssd1 vssd1 vccd1 vccd1 _3640_/A sky130_fd_sc_hd__or2_1
XFILLER_0_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5309_ _5311_/CLK _5309_/D vssd1 vssd1 vccd1 vccd1 _5309_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold4 phase_in[2] vssd1 vssd1 vccd1 vccd1 hold4/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3990_ _3990_/A _3990_/B _3990_/C vssd1 vssd1 vccd1 vccd1 _3993_/A sky130_fd_sc_hd__or3_4
X_2941_ _2940_/X _2936_/A _2878_/X vssd1 vssd1 vccd1 vccd1 _2941_/X sky130_fd_sc_hd__a21o_1
X_2872_ _3642_/A vssd1 vssd1 vccd1 vccd1 _2901_/A sky130_fd_sc_hd__buf_2
XFILLER_30_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4611_ _4673_/B vssd1 vssd1 vccd1 vccd1 _4611_/Y sky130_fd_sc_hd__inv_2
X_4542_ _4542_/A vssd1 vssd1 vccd1 vccd1 _4542_/X sky130_fd_sc_hd__buf_2
X_4473_ _4807_/A vssd1 vssd1 vccd1 vccd1 _4473_/X sky130_fd_sc_hd__clkbuf_2
X_3424_ _3864_/B _5131_/Q _3677_/B vssd1 vssd1 vccd1 vccd1 _3424_/Y sky130_fd_sc_hd__o21ai_1
X_3355_ _5224_/Q _3321_/X _3353_/X _3354_/Y _3316_/X vssd1 vssd1 vccd1 vccd1 _5224_/D
+ sky130_fd_sc_hd__o221a_1
X_3286_ _5236_/Q _3253_/X _3246_/X _3285_/X vssd1 vssd1 vccd1 vccd1 _5236_/D sky130_fd_sc_hd__o211a_1
XFILLER_85_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5025_ _5027_/CLK _5025_/D vssd1 vssd1 vccd1 vccd1 _5025_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4809_ _3879_/X _4806_/X _4807_/X _4808_/Y vssd1 vssd1 vccd1 vccd1 _5035_/D sky130_fd_sc_hd__o211a_1
XFILLER_79_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140_ _3747_/B _5174_/Q vssd1 vssd1 vccd1 vccd1 _3141_/A sky130_fd_sc_hd__nand2_1
XFILLER_67_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_67_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3071_ _3125_/A _3123_/A _3287_/A vssd1 vssd1 vccd1 vccd1 _3278_/A sky130_fd_sc_hd__a21o_1
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3973_ _4017_/A vssd1 vssd1 vccd1 vccd1 _3973_/Y sky130_fd_sc_hd__inv_2
XFILLER_62_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2924_ _3321_/A vssd1 vssd1 vccd1 vccd1 _2924_/X sky130_fd_sc_hd__clkbuf_2
X_2855_ _2865_/B _2865_/C _2865_/A vssd1 vssd1 vccd1 vccd1 _2867_/C sky130_fd_sc_hd__o21ai_1
X_4525_ _4525_/A _4525_/B vssd1 vssd1 vccd1 vccd1 _4527_/B sky130_fd_sc_hd__nor2_1
X_2786_ _5316_/Q _5049_/Q vssd1 vssd1 vccd1 vccd1 _2787_/B sky130_fd_sc_hd__nand2_1
X_4456_ _4453_/X _5075_/Q _3911_/X _4455_/X vssd1 vssd1 vccd1 vccd1 _5075_/D sky130_fd_sc_hd__o211a_1
X_3407_ _3407_/A _3407_/B vssd1 vssd1 vccd1 vccd1 _3407_/Y sky130_fd_sc_hd__nor2_2
X_4387_ _4387_/A _4392_/A vssd1 vssd1 vccd1 vccd1 _4388_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3338_ _3338_/A vssd1 vssd1 vccd1 vccd1 _3339_/B sky130_fd_sc_hd__inv_2
XFILLER_65_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3269_ _3321_/A vssd1 vssd1 vccd1 vccd1 _3269_/X sky130_fd_sc_hd__clkbuf_2
X_5008_ _5118_/CLK hold28/X vssd1 vssd1 vccd1 vccd1 _5008_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2640_ _4631_/A _2634_/X _2619_/X _2639_/Y vssd1 vssd1 vccd1 vccd1 _5287_/D sky130_fd_sc_hd__o211a_1
XFILLER_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2571_ _5303_/Q _2567_/X _2563_/X _2570_/Y vssd1 vssd1 vccd1 vccd1 _5303_/D sky130_fd_sc_hd__o211a_1
X_5290_ _5292_/CLK _5290_/D vssd1 vssd1 vccd1 vccd1 _5290_/Q sky130_fd_sc_hd__dfxtp_1
X_4310_ _4310_/A _4648_/B vssd1 vssd1 vccd1 vccd1 _4312_/A sky130_fd_sc_hd__nand2_1
X_4241_ _4405_/B _4591_/B vssd1 vssd1 vccd1 vccd1 _4241_/Y sky130_fd_sc_hd__nor2_1
X_4172_ _4734_/A _4172_/B _4172_/C vssd1 vssd1 vccd1 vccd1 _5097_/D sky130_fd_sc_hd__nor3_1
XFILLER_67_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3123_ _3123_/A vssd1 vssd1 vccd1 vccd1 _3287_/B sky130_fd_sc_hd__inv_2
X_3054_ _3739_/B _5177_/Q vssd1 vssd1 vccd1 vccd1 _3064_/A sky130_fd_sc_hd__and2_1
XFILLER_48_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3956_ _4347_/A _4342_/A _4352_/A _4356_/A vssd1 vssd1 vccd1 vccd1 _4145_/B sky130_fd_sc_hd__or4_4
XFILLER_50_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2907_ _2901_/X _2903_/X _2892_/X _2906_/Y vssd1 vssd1 vccd1 vccd1 _5274_/D sky130_fd_sc_hd__o211a_1
XFILLER_50_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3887_ _3907_/A vssd1 vssd1 vccd1 vccd1 _3887_/X sky130_fd_sc_hd__clkbuf_2
X_2838_ _5283_/Q vssd1 vssd1 vccd1 vccd1 _3713_/B sky130_fd_sc_hd__inv_2
X_2769_ _2769_/A _2769_/B vssd1 vssd1 vccd1 vccd1 _2770_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4508_ _4785_/A vssd1 vssd1 vccd1 vccd1 _4508_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4439_ _4381_/A _4445_/C _4396_/C vssd1 vssd1 vccd1 vccd1 _4439_/X sky130_fd_sc_hd__o21a_1
XFILLER_58_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_89_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3810_ _3823_/A vssd1 vssd1 vccd1 vccd1 _3820_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_32_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4790_ _4790_/A _4790_/B vssd1 vssd1 vccd1 vccd1 _4806_/B sky130_fd_sc_hd__nor2_2
XFILLER_60_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3741_ _3754_/A vssd1 vssd1 vccd1 vccd1 _3741_/X sky130_fd_sc_hd__buf_1
XFILLER_9_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3672_ _5196_/Q _3668_/X _3646_/X _3671_/X vssd1 vssd1 vccd1 vccd1 _5196_/D sky130_fd_sc_hd__o211a_1
X_2623_ _5289_/Q _2604_/X _2619_/X _2622_/Y vssd1 vssd1 vccd1 vccd1 _5289_/D sky130_fd_sc_hd__o211a_1
X_2554_ _2565_/A _4601_/A vssd1 vssd1 vccd1 vccd1 _2554_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5273_ _5277_/CLK _5273_/D vssd1 vssd1 vccd1 vccd1 _5273_/Q sky130_fd_sc_hd__dfxtp_1
X_4224_ _4226_/A _4221_/Y _4222_/Y _3879_/A vssd1 vssd1 vccd1 vccd1 _4224_/X sky130_fd_sc_hd__a31o_1
X_4155_ _4155_/A _4155_/B vssd1 vssd1 vccd1 vccd1 _5102_/D sky130_fd_sc_hd__nor2_1
XFILLER_55_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3106_ _3103_/B _3324_/B _3103_/A vssd1 vssd1 vccd1 vccd1 _3310_/B sky130_fd_sc_hd__o21ba_1
XFILLER_46_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4086_ _4282_/A _4304_/A vssd1 vssd1 vccd1 vccd1 _4190_/B sky130_fd_sc_hd__nor2_4
XFILLER_55_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3037_ _3037_/A vssd1 vssd1 vccd1 vccd1 _3174_/A sky130_fd_sc_hd__inv_2
XFILLER_36_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4988_ _4992_/CLK hold46/X vssd1 vssd1 vccd1 vccd1 _4988_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3939_ _4940_/A _5009_/Q _5121_/Q _3923_/Y vssd1 vssd1 vccd1 vccd1 _3939_/X sky130_fd_sc_hd__a22o_1
XFILLER_87_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_74_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 hold8/X vssd1 vssd1 vccd1 vccd1 hold7/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4911_ _4913_/A _4911_/B vssd1 vssd1 vccd1 vccd1 _5004_/D sky130_fd_sc_hd__nor2_1
X_4842_ _4842_/A _4842_/B vssd1 vssd1 vccd1 vccd1 _4842_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4773_ _4779_/B _4779_/A vssd1 vssd1 vccd1 vccd1 _4780_/A sky130_fd_sc_hd__or2_1
X_3724_ _3726_/A _3724_/B vssd1 vssd1 vccd1 vccd1 _3724_/Y sky130_fd_sc_hd__nand2_1
X_3655_ _3655_/A _3655_/B vssd1 vssd1 vccd1 vccd1 _3655_/Y sky130_fd_sc_hd__nor2_1
X_2606_ _5026_/Q vssd1 vssd1 vccd1 vccd1 _4853_/A sky130_fd_sc_hd__inv_2
X_3586_ _3586_/A _3586_/B vssd1 vssd1 vccd1 vccd1 _3586_/Y sky130_fd_sc_hd__nand2_1
X_2537_ _5044_/Q vssd1 vssd1 vccd1 vccd1 _4704_/A sky130_fd_sc_hd__inv_2
X_5256_ _5267_/CLK _5256_/D vssd1 vssd1 vccd1 vccd1 _5256_/Q sky130_fd_sc_hd__dfxtp_1
X_4207_ _4207_/A vssd1 vssd1 vccd1 vccd1 _4208_/A sky130_fd_sc_hd__inv_2
XFILLER_57_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_68_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5187_ _5283_/CLK _5187_/D vssd1 vssd1 vccd1 vccd1 _5187_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4138_ _4149_/A _5105_/Q _4138_/C vssd1 vssd1 vccd1 vccd1 _4144_/B sky130_fd_sc_hd__nand3_1
X_4069_ _5086_/Q vssd1 vssd1 vccd1 vccd1 _4558_/A sky130_fd_sc_hd__inv_2
XFILLER_28_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_78_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3440_ _5131_/Q vssd1 vssd1 vccd1 vccd1 _3441_/B sky130_fd_sc_hd__inv_2
X_3371_ _3531_/A vssd1 vssd1 vccd1 vccd1 _3371_/Y sky130_fd_sc_hd__inv_2
X_5110_ _5112_/CLK _5110_/D vssd1 vssd1 vccd1 vccd1 _5110_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5041_ _5076_/CLK _5041_/D vssd1 vssd1 vccd1 vccd1 _5041_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_77_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4825_ _4824_/B _4824_/A _3907_/A vssd1 vssd1 vccd1 vccd1 _4825_/X sky130_fd_sc_hd__a21o_1
X_4756_ _4567_/X _4752_/X _4754_/X _4550_/X _4755_/Y vssd1 vssd1 vccd1 vccd1 _5046_/D
+ sky130_fd_sc_hd__o311a_1
X_3707_ _3713_/A _3707_/B vssd1 vssd1 vccd1 vccd1 _3707_/Y sky130_fd_sc_hd__nand2_1
X_4687_ _4801_/A _4801_/B _4806_/A vssd1 vssd1 vccd1 vccd1 _4688_/B sky130_fd_sc_hd__or3_1
X_3638_ _3638_/A _3638_/B vssd1 vssd1 vccd1 vccd1 _3647_/A sky130_fd_sc_hd__nor2_1
X_3569_ _3569_/A _3569_/B vssd1 vssd1 vccd1 vccd1 _3569_/Y sky130_fd_sc_hd__nor2_1
X_5308_ _5311_/CLK _5308_/D vssd1 vssd1 vccd1 vccd1 _5308_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_0_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5239_ _5268_/CLK _5239_/D vssd1 vssd1 vccd1 vccd1 _5239_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_83_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold5 hold5/A vssd1 vssd1 vccd1 vccd1 hold5/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ _2940_/A _2940_/B vssd1 vssd1 vccd1 vccd1 _2940_/X sky130_fd_sc_hd__or2_1
XFILLER_15_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2871_ _2871_/A _2874_/B _2871_/C vssd1 vssd1 vccd1 vccd1 _2874_/A sky130_fd_sc_hd__nand3_2
XPHY_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4610_ _4818_/A _4610_/B vssd1 vssd1 vccd1 vccd1 _4673_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4541_ _4541_/A _4541_/B vssd1 vssd1 vccd1 vccd1 _4541_/Y sky130_fd_sc_hd__nand2_1
XFILLER_7_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4472_ _4434_/X _4469_/Y _4470_/X _2915_/X _4471_/Y vssd1 vssd1 vccd1 vccd1 _5072_/D
+ sky130_fd_sc_hd__o311a_1
X_3423_ _5130_/Q _3866_/B vssd1 vssd1 vccd1 vccd1 _3677_/B sky130_fd_sc_hd__or2_2
X_3354_ _3346_/A _3350_/X _3352_/Y _2888_/X vssd1 vssd1 vccd1 vccd1 _3354_/Y sky130_fd_sc_hd__o31ai_1
X_3285_ _3279_/X _3284_/Y _2963_/X vssd1 vssd1 vccd1 vccd1 _3285_/X sky130_fd_sc_hd__a21o_1
X_5024_ _5027_/CLK _5024_/D vssd1 vssd1 vccd1 vccd1 _5024_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_26_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4808_ _4808_/A _4846_/B vssd1 vssd1 vccd1 vccd1 _4808_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4739_ _4739_/A _4739_/B vssd1 vssd1 vccd1 vccd1 _4741_/B sky130_fd_sc_hd__nor2_1
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_67_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3070_ _5171_/Q _3756_/B vssd1 vssd1 vccd1 vccd1 _3287_/A sky130_fd_sc_hd__nor2_1
XFILLER_85_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3972_ _4992_/D _3974_/A vssd1 vssd1 vccd1 vccd1 _4017_/A sky130_fd_sc_hd__nor2_4
XFILLER_50_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2923_ _3769_/A vssd1 vssd1 vccd1 vccd1 _3321_/A sky130_fd_sc_hd__clkbuf_2
X_2854_ _2871_/A _2854_/B vssd1 vssd1 vccd1 vccd1 _2865_/C sky130_fd_sc_hd__and2_1
X_2785_ _5316_/Q _5049_/Q vssd1 vssd1 vccd1 vccd1 _2787_/A sky130_fd_sc_hd__or2_1
X_4524_ _4531_/B _4531_/A vssd1 vssd1 vccd1 vccd1 _4527_/A sky130_fd_sc_hd__or2_1
X_4455_ _4454_/X _4449_/A _4204_/X vssd1 vssd1 vccd1 vccd1 _4455_/X sky130_fd_sc_hd__a21o_1
X_3406_ _3406_/A _3406_/B vssd1 vssd1 vccd1 vccd1 _3407_/B sky130_fd_sc_hd__nor2_1
X_4386_ _4386_/A _4713_/B vssd1 vssd1 vccd1 vccd1 _4392_/A sky130_fd_sc_hd__nor2_1
X_3337_ _3337_/A _3337_/B vssd1 vssd1 vccd1 vccd1 _3338_/A sky130_fd_sc_hd__nand2_1
X_3268_ _3265_/Y _3267_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _5240_/D sky130_fd_sc_hd__o21a_1
X_5007_ _5097_/CLK hold33/X vssd1 vssd1 vccd1 vccd1 _5007_/Q sky130_fd_sc_hd__dfxtp_1
X_3199_ _3199_/A _3199_/B _3199_/C vssd1 vssd1 vccd1 vccd1 _3199_/Y sky130_fd_sc_hd__nand3_2
XFILLER_45_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_76_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _2584_/A _4682_/A vssd1 vssd1 vccd1 vccd1 _2570_/Y sky130_fd_sc_hd__nand2_1
XFILLER_4_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4240_ _5081_/Q vssd1 vssd1 vccd1 vccd1 _4591_/B sky130_fd_sc_hd__inv_2
X_4171_ _4164_/A _4111_/X _4112_/X _4173_/C _5097_/Q vssd1 vssd1 vccd1 vccd1 _4172_/B
+ sky130_fd_sc_hd__a41oi_1
XFILLER_67_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3122_ _3118_/B _3300_/B _3118_/A vssd1 vssd1 vccd1 vccd1 _3288_/B sky130_fd_sc_hd__o21ba_1
X_3053_ _5177_/Q _3739_/B vssd1 vssd1 vccd1 vccd1 _3055_/A sky130_fd_sc_hd__nor2_1
XFILLER_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3955_ _4354_/A vssd1 vssd1 vccd1 vccd1 _4356_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2906_ _3276_/A _3737_/B vssd1 vssd1 vccd1 vccd1 _2906_/Y sky130_fd_sc_hd__nand2_1
XFILLER_31_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3886_ _4764_/A vssd1 vssd1 vccd1 vccd1 _3907_/A sky130_fd_sc_hd__buf_2
X_2837_ _4550_/A vssd1 vssd1 vccd1 vccd1 _2837_/X sky130_fd_sc_hd__buf_2
X_2768_ _2762_/Y _2753_/A _2764_/B vssd1 vssd1 vccd1 vccd1 _2769_/A sky130_fd_sc_hd__o21ai_1
X_2699_ _5292_/Q vssd1 vssd1 vccd1 vccd1 _2700_/A sky130_fd_sc_hd__inv_2
X_4507_ _4507_/A _4507_/B vssd1 vssd1 vccd1 vccd1 _4507_/Y sky130_fd_sc_hd__nor2_1
X_4438_ _4444_/B _4438_/B vssd1 vssd1 vccd1 vccd1 _4445_/C sky130_fd_sc_hd__nor2_1
XFILLER_86_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_76_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4369_ _5075_/Q vssd1 vssd1 vccd1 vccd1 _4701_/B sky130_fd_sc_hd__inv_2
XFILLER_86_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3740_ _5177_/Q _3728_/X _3736_/X _3739_/Y vssd1 vssd1 vccd1 vccd1 _5177_/D sky130_fd_sc_hd__o211a_1
X_3671_ _3669_/X _3670_/Y _2848_/X vssd1 vssd1 vccd1 vccd1 _3671_/X sky130_fd_sc_hd__a21o_1
X_2622_ _2622_/A _4872_/A vssd1 vssd1 vccd1 vccd1 _2622_/Y sky130_fd_sc_hd__nand2_1
X_2553_ _5040_/Q vssd1 vssd1 vccd1 vccd1 _4601_/A sky130_fd_sc_hd__inv_2
X_5272_ _5277_/CLK _5272_/D vssd1 vssd1 vccd1 vccd1 _5272_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4223_ _4226_/A _4221_/Y _4222_/Y vssd1 vssd1 vccd1 vccd1 _4223_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_68_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4154_ _4154_/A _4238_/B vssd1 vssd1 vccd1 vccd1 _4155_/B sky130_fd_sc_hd__nand2_1
X_4085_ _5089_/Q vssd1 vssd1 vccd1 vccd1 _4304_/A sky130_fd_sc_hd__inv_2
XFILLER_28_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3105_ _3079_/Y _3333_/A _3096_/Y _3104_/Y vssd1 vssd1 vccd1 vccd1 _3310_/A sky130_fd_sc_hd__o211ai_2
X_3036_ _5182_/Q _3726_/B vssd1 vssd1 vccd1 vccd1 _3037_/A sky130_fd_sc_hd__nor2_2
XFILLER_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4987_ _4987_/CLK hold45/X vssd1 vssd1 vccd1 vccd1 hold46/A sky130_fd_sc_hd__dfxtp_1
XFILLER_23_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3938_ _5009_/Q vssd1 vssd1 vccd1 vccd1 _3938_/Y sky130_fd_sc_hd__inv_2
X_3869_ _5129_/Q _3862_/X _3857_/X _3868_/Y vssd1 vssd1 vccd1 vccd1 _5129_/D sky130_fd_sc_hd__o211a_1
XFILLER_11_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput17 hold10/X vssd1 vssd1 vccd1 vccd1 hold9/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4910_ _4910_/A hold38/X vssd1 vssd1 vccd1 vccd1 hold39/A sky130_fd_sc_hd__or2_1
X_4841_ _4845_/B _4650_/A _4650_/B vssd1 vssd1 vccd1 vccd1 _4842_/B sky130_fd_sc_hd__a21bo_1
XFILLER_20_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4772_ _4697_/B _4787_/B _4604_/X vssd1 vssd1 vccd1 vccd1 _4779_/A sky130_fd_sc_hd__o21ba_1
XFILLER_20_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3723_ _3762_/A vssd1 vssd1 vccd1 vccd1 _3723_/X sky130_fd_sc_hd__buf_1
X_3654_ _3855_/B _5134_/Q _3653_/X vssd1 vssd1 vccd1 vccd1 _3655_/B sky130_fd_sc_hd__o21a_1
X_2605_ _2605_/A vssd1 vssd1 vccd1 vccd1 _2622_/A sky130_fd_sc_hd__buf_1
X_3585_ _3646_/A vssd1 vssd1 vccd1 vccd1 _3585_/X sky130_fd_sc_hd__clkbuf_2
X_2536_ _5312_/Q _2528_/X _2522_/X _2535_/Y vssd1 vssd1 vccd1 vccd1 _5312_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5255_ _5283_/CLK _5255_/D vssd1 vssd1 vccd1 vccd1 _5255_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4206_ _4206_/A _4238_/B _4206_/C vssd1 vssd1 vccd1 vccd1 _5087_/D sky130_fd_sc_hd__and3_1
XFILLER_3_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5186_ _5250_/CLK _5186_/D vssd1 vssd1 vccd1 vccd1 _5186_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4137_ _4137_/A vssd1 vssd1 vccd1 vccd1 _4138_/C sky130_fd_sc_hd__inv_2
XFILLER_83_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4068_ _4070_/A _4053_/C _5085_/Q vssd1 vssd1 vccd1 vccd1 _4222_/A sky130_fd_sc_hd__a21o_2
XFILLER_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3019_ _3023_/B _3018_/X _2888_/X vssd1 vssd1 vccd1 vccd1 _3019_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3370_ _5156_/Q _3798_/B vssd1 vssd1 vccd1 vccd1 _3531_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5040_ _5040_/CLK _5040_/D vssd1 vssd1 vccd1 vccd1 _5040_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4824_ _4824_/A _4824_/B vssd1 vssd1 vccd1 vccd1 _4824_/Y sky130_fd_sc_hd__nor2_1
X_4755_ _4755_/A _4799_/A vssd1 vssd1 vccd1 vccd1 _4755_/Y sky130_fd_sc_hd__nand2_1
XFILLER_21_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3706_ _5190_/Q _2524_/A _3704_/Y _3705_/Y _3695_/X vssd1 vssd1 vccd1 vccd1 _5190_/D
+ sky130_fd_sc_hd__o221a_1
X_4686_ _4686_/A _4686_/B vssd1 vssd1 vccd1 vccd1 _4806_/A sky130_fd_sc_hd__nand2_1
X_3637_ _5202_/Q _3613_/X _3585_/X _3636_/X vssd1 vssd1 vccd1 vccd1 _5202_/D sky130_fd_sc_hd__o211a_1
X_3568_ _3568_/A _3568_/B vssd1 vssd1 vccd1 vccd1 _3569_/B sky130_fd_sc_hd__nor2_1
X_2519_ _5315_/Q _2506_/X _2510_/X _2518_/Y vssd1 vssd1 vccd1 vccd1 _5315_/D sky130_fd_sc_hd__o211a_1
X_5307_ _5311_/CLK _5307_/D vssd1 vssd1 vccd1 vccd1 _5307_/Q sky130_fd_sc_hd__dfxtp_1
X_3499_ _3582_/C _3499_/B vssd1 vssd1 vccd1 vccd1 _3586_/B sky130_fd_sc_hd__nand2_1
X_5238_ _5252_/CLK _5238_/D vssd1 vssd1 vccd1 vccd1 _5238_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5169_ _5171_/CLK _5169_/D vssd1 vssd1 vccd1 vccd1 _5169_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_79_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold6 phase_in[5] vssd1 vssd1 vccd1 vccd1 hold6/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_47_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_74_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2870_ _2864_/Y _2867_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _5280_/D sky130_fd_sc_hd__o21a_1
XPHY_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_10_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5124_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_11_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4540_ _4807_/A vssd1 vssd1 vccd1 vccd1 _4540_/X sky130_fd_sc_hd__buf_2
XFILLER_7_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4471_ _4528_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4471_/Y sky130_fd_sc_hd__nand2_1
X_3422_ _5226_/Q vssd1 vssd1 vccd1 vccd1 _3866_/B sky130_fd_sc_hd__inv_2
X_3353_ _3346_/A _3350_/X _3352_/Y vssd1 vssd1 vccd1 vccd1 _3353_/X sky130_fd_sc_hd__o21a_1
X_3284_ _3284_/A _3284_/B vssd1 vssd1 vccd1 vccd1 _3284_/Y sky130_fd_sc_hd__nand2_1
X_5023_ _5085_/CLK _5023_/D vssd1 vssd1 vccd1 vccd1 _5023_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_65_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_70_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4807_ _4807_/A vssd1 vssd1 vccd1 vccd1 _4807_/X sky130_fd_sc_hd__clkbuf_2
X_2999_ _5258_/Q _2939_/X _2961_/X _2998_/Y vssd1 vssd1 vccd1 vccd1 _5258_/D sky130_fd_sc_hd__o211a_1
X_4738_ _4736_/X _4737_/Y _4116_/A vssd1 vssd1 vccd1 vccd1 _5049_/D sky130_fd_sc_hd__a21oi_1
X_4669_ _4821_/A _4821_/B _4668_/Y vssd1 vssd1 vccd1 vccd1 _4810_/A sky130_fd_sc_hd__o21bai_1
XFILLER_88_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_85_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3971_ _4992_/Q vssd1 vssd1 vccd1 vccd1 _3974_/A sky130_fd_sc_hd__inv_2
X_2922_ _2920_/X _2921_/Y _4913_/A vssd1 vssd1 vccd1 vccd1 _5272_/D sky130_fd_sc_hd__a21oi_1
X_2853_ _2853_/A _2853_/B vssd1 vssd1 vccd1 vccd1 _2871_/A sky130_fd_sc_hd__nand2_1
X_2784_ _2836_/A _2836_/B _2834_/B vssd1 vssd1 vccd1 vccd1 _2784_/Y sky130_fd_sc_hd__a21oi_1
X_4523_ _4523_/A _4523_/B vssd1 vssd1 vccd1 vccd1 _4531_/A sky130_fd_sc_hd__and2_1
X_4454_ _4454_/A _4454_/B _4378_/A vssd1 vssd1 vccd1 vccd1 _4454_/X sky130_fd_sc_hd__or3b_2
X_3405_ _3608_/A _3485_/A vssd1 vssd1 vccd1 vccd1 _3405_/Y sky130_fd_sc_hd__nor2_2
X_4385_ _5078_/Q vssd1 vssd1 vccd1 vccd1 _4713_/B sky130_fd_sc_hd__inv_2
XFILLER_58_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3336_ _3337_/A _3337_/B _3339_/A _2901_/A vssd1 vssd1 vccd1 vccd1 _3336_/X sky130_fd_sc_hd__a31o_1
XFILLER_85_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5006_ _5118_/CLK hold37/X vssd1 vssd1 vccd1 vccd1 _5006_/Q sky130_fd_sc_hd__dfxtp_1
X_3267_ _3267_/A _3862_/A _3267_/C vssd1 vssd1 vccd1 vccd1 _3267_/X sky130_fd_sc_hd__and3_1
X_3198_ _3204_/A _3198_/B _3198_/C vssd1 vssd1 vccd1 vccd1 _3199_/A sky130_fd_sc_hd__nand3b_1
XFILLER_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4170_ _5098_/Q _4172_/C _4169_/Y vssd1 vssd1 vccd1 vccd1 _5098_/D sky130_fd_sc_hd__o21a_1
XFILLER_67_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3121_ _3298_/A _3298_/B _3120_/X vssd1 vssd1 vccd1 vccd1 _3288_/A sky130_fd_sc_hd__o21bai_1
XFILLER_67_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3052_ _3064_/B _3052_/B vssd1 vssd1 vccd1 vccd1 _3266_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3954_ _5099_/Q vssd1 vssd1 vccd1 vccd1 _4354_/A sky130_fd_sc_hd__inv_2
X_3885_ _4199_/A vssd1 vssd1 vccd1 vccd1 _4764_/A sky130_fd_sc_hd__clkbuf_2
X_2905_ _5274_/Q vssd1 vssd1 vccd1 vccd1 _3737_/B sky130_fd_sc_hd__inv_2
X_2836_ _2836_/A _2836_/B _2836_/C vssd1 vssd1 vccd1 vccd1 _2836_/X sky130_fd_sc_hd__and3_1
X_2767_ _2885_/A vssd1 vssd1 vccd1 vccd1 _2767_/Y sky130_fd_sc_hd__inv_2
X_2698_ _2698_/A _5291_/Q vssd1 vssd1 vccd1 vccd1 _2798_/A sky130_fd_sc_hd__nand2_1
X_4506_ _4506_/A _4506_/B vssd1 vssd1 vccd1 vccd1 _4507_/B sky130_fd_sc_hd__and2_1
X_4437_ _4444_/B _4438_/B _4388_/A _4383_/A vssd1 vssd1 vccd1 vccd1 _4437_/X sky130_fd_sc_hd__o211a_1
XFILLER_86_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4368_ _4474_/A _4474_/B _4367_/Y vssd1 vssd1 vccd1 vccd1 _4454_/B sky130_fd_sc_hd__a21oi_4
XFILLER_86_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4299_ _4568_/A _4571_/B _4576_/B vssd1 vssd1 vccd1 vccd1 _4559_/A sky130_fd_sc_hd__nand3_4
X_3319_ _3311_/X _3318_/Y _3306_/X vssd1 vssd1 vccd1 vccd1 _3319_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3670_ _3670_/A _3670_/B vssd1 vssd1 vccd1 vccd1 _3670_/Y sky130_fd_sc_hd__nand2_1
X_2621_ _3000_/A vssd1 vssd1 vccd1 vccd1 _4872_/A sky130_fd_sc_hd__inv_2
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2552_ _5308_/Q _2548_/X _2544_/X _2551_/Y vssd1 vssd1 vccd1 vccd1 _5308_/D sky130_fd_sc_hd__o211a_1
X_5271_ _5288_/CLK _5271_/D vssd1 vssd1 vccd1 vccd1 _5271_/Q sky130_fd_sc_hd__dfxtp_1
X_4222_ _4222_/A _4222_/B vssd1 vssd1 vccd1 vccd1 _4222_/Y sky130_fd_sc_hd__nand2_1
XFILLER_68_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4153_ _4169_/B _4152_/X _5102_/Q vssd1 vssd1 vccd1 vccd1 _4155_/A sky130_fd_sc_hd__a21oi_1
XFILLER_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4084_ _5090_/Q vssd1 vssd1 vccd1 vccd1 _4282_/A sky130_fd_sc_hd__inv_2
X_3104_ _3330_/B _3325_/A vssd1 vssd1 vccd1 vccd1 _3104_/Y sky130_fd_sc_hd__nor2_1
XFILLER_83_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3035_ _5278_/Q vssd1 vssd1 vccd1 vccd1 _3726_/B sky130_fd_sc_hd__inv_2
XFILLER_36_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4986_ _4990_/CLK _4986_/D vssd1 vssd1 vccd1 vccd1 _4986_/Q sky130_fd_sc_hd__dfxtp_1
XPHY_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3937_ _5014_/Q vssd1 vssd1 vccd1 vccd1 _3937_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3868_ _3873_/A _3868_/B vssd1 vssd1 vccd1 vccd1 _3868_/Y sky130_fd_sc_hd__nand2_1
X_2819_ _2793_/C _2793_/B _2793_/A _2818_/Y vssd1 vssd1 vccd1 vccd1 _2819_/Y sky130_fd_sc_hd__o22ai_1
X_3799_ _5156_/Q _3796_/X _3791_/X _3798_/Y vssd1 vssd1 vccd1 vccd1 _5156_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput18 hold6/X vssd1 vssd1 vccd1 vccd1 hold5/A sky130_fd_sc_hd__clkbuf_1
XFILLER_10_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_65_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4840_ _4840_/A _4840_/B vssd1 vssd1 vccd1 vccd1 _4845_/B sky130_fd_sc_hd__or2_1
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4771_ _4771_/A _4771_/B vssd1 vssd1 vccd1 vccd1 _4787_/B sky130_fd_sc_hd__and2_1
X_3722_ _5184_/Q _3715_/X _3710_/X _3721_/Y vssd1 vssd1 vccd1 vccd1 _5184_/D sky130_fd_sc_hd__o211a_1
XFILLER_9_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3653_ _3658_/B _3658_/A vssd1 vssd1 vccd1 vccd1 _3653_/X sky130_fd_sc_hd__or2_1
X_2604_ _2604_/A vssd1 vssd1 vccd1 vccd1 _2604_/X sky130_fd_sc_hd__clkbuf_2
X_3584_ _3581_/X _2506_/X _3582_/Y _3583_/Y vssd1 vssd1 vccd1 vccd1 _5213_/D sky130_fd_sc_hd__a31oi_1
X_2535_ _2546_/A _4710_/A vssd1 vssd1 vccd1 vccd1 _2535_/Y sky130_fd_sc_hd__nand2_1
X_5254_ _5288_/CLK _5254_/D vssd1 vssd1 vccd1 vccd1 _5254_/Q sky130_fd_sc_hd__dfxtp_2
X_4205_ _4204_/X _4201_/C _4289_/A vssd1 vssd1 vccd1 vccd1 _4206_/C sky130_fd_sc_hd__o21ai_1
X_5185_ _5250_/CLK _5185_/D vssd1 vssd1 vccd1 vccd1 _5185_/Q sky130_fd_sc_hd__dfxtp_1
X_4136_ _4149_/B _4136_/B vssd1 vssd1 vccd1 vccd1 _4137_/A sky130_fd_sc_hd__nand2_1
XFILLER_83_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_68_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4067_ _4222_/B _4226_/B _4067_/C vssd1 vssd1 vccd1 vccd1 _4208_/D sky130_fd_sc_hd__nand3_4
X_3018_ _3017_/Y _3018_/B vssd1 vssd1 vccd1 vccd1 _3018_/X sky130_fd_sc_hd__and2b_1
XPHY_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4969_ _5317_/Q _2841_/X _4197_/B _4968_/Y vssd1 vssd1 vccd1 vccd1 _5317_/D sky130_fd_sc_hd__o211a_1
XPHY_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4823_ _4823_/A _4823_/B vssd1 vssd1 vccd1 vccd1 _4824_/B sky130_fd_sc_hd__nand2_1
XFILLER_21_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4754_ _4709_/A _4758_/B _4716_/B vssd1 vssd1 vccd1 vccd1 _4754_/X sky130_fd_sc_hd__o21a_1
X_3705_ _3705_/A _3705_/B vssd1 vssd1 vccd1 vccd1 _3705_/Y sky130_fd_sc_hd__nand2_1
X_4685_ _4808_/A _4685_/B vssd1 vssd1 vccd1 vccd1 _4686_/B sky130_fd_sc_hd__nand2_1
X_3636_ _3630_/X _3635_/Y _3615_/X vssd1 vssd1 vccd1 vccd1 _3636_/X sky130_fd_sc_hd__a21o_1
X_3567_ _3572_/B _3567_/B vssd1 vssd1 vccd1 vccd1 _3568_/B sky130_fd_sc_hd__nor2_1
X_2518_ _2524_/A _4725_/A vssd1 vssd1 vccd1 vccd1 _2518_/Y sky130_fd_sc_hd__nand2_1
X_5306_ _5311_/CLK _5306_/D vssd1 vssd1 vccd1 vccd1 _5306_/Q sky130_fd_sc_hd__dfxtp_1
X_3498_ _3818_/B _5148_/Q vssd1 vssd1 vccd1 vccd1 _3499_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5237_ _5268_/CLK _5237_/D vssd1 vssd1 vccd1 vccd1 _5237_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_84_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5168_ _5171_/CLK _5168_/D vssd1 vssd1 vccd1 vccd1 _5168_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4119_ _4382_/A _4119_/B _4119_/C vssd1 vssd1 vccd1 vccd1 _4125_/C sky130_fd_sc_hd__nor3_4
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5099_ _5109_/CLK _5099_/D vssd1 vssd1 vccd1 vccd1 _5099_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_83_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_79_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xhold7 hold7/A vssd1 vssd1 vccd1 vccd1 hold7/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4470_ _4470_/A _4470_/B vssd1 vssd1 vccd1 vccd1 _4470_/X sky130_fd_sc_hd__and2_1
X_3421_ _5227_/Q vssd1 vssd1 vccd1 vccd1 _3864_/B sky130_fd_sc_hd__inv_2
X_3352_ _3352_/A vssd1 vssd1 vccd1 vccd1 _3352_/Y sky130_fd_sc_hd__inv_2
X_3283_ _5237_/Q _3269_/X _3281_/Y _3282_/X _3262_/X vssd1 vssd1 vccd1 vccd1 _5237_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_85_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5022_ _5027_/CLK _5022_/D vssd1 vssd1 vccd1 vccd1 _5022_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4806_ _4806_/A _4806_/B vssd1 vssd1 vccd1 vccd1 _4806_/X sky130_fd_sc_hd__xor2_1
X_2998_ _2989_/A _2997_/X _2951_/X vssd1 vssd1 vccd1 vccd1 _2998_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4737_ _4799_/A _5049_/Q vssd1 vssd1 vccd1 vccd1 _4737_/Y sky130_fd_sc_hd__nand2_1
X_4668_ _4827_/A _4820_/A vssd1 vssd1 vccd1 vccd1 _4668_/Y sky130_fd_sc_hd__nand2_1
X_3619_ _3625_/B _3625_/A vssd1 vssd1 vccd1 vccd1 _3622_/A sky130_fd_sc_hd__or2_1
X_4599_ _4599_/A vssd1 vssd1 vccd1 vccd1 _4775_/A sky130_fd_sc_hd__inv_2
XFILLER_48_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_85_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3970_ _4988_/Q _3970_/B vssd1 vssd1 vccd1 vccd1 _4023_/A sky130_fd_sc_hd__nor2_2
XFILLER_62_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2921_ _3542_/A _5272_/Q vssd1 vssd1 vccd1 vccd1 _2921_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2852_ _5282_/Q _2841_/X _2846_/Y _2849_/X _4902_/A vssd1 vssd1 vccd1 vccd1 _5282_/D
+ sky130_fd_sc_hd__o221a_1
X_2783_ _4739_/A _2783_/B vssd1 vssd1 vccd1 vccd1 _2834_/B sky130_fd_sc_hd__nor2_1
X_4522_ _4453_/X _5063_/Q _4473_/X _4521_/Y vssd1 vssd1 vccd1 vccd1 _5063_/D sky130_fd_sc_hd__o211a_1
XFILLER_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4453_ _4742_/B vssd1 vssd1 vccd1 vccd1 _4453_/X sky130_fd_sc_hd__clkbuf_2
X_3404_ _5142_/Q _3833_/B vssd1 vssd1 vccd1 vccd1 _3485_/A sky130_fd_sc_hd__nor2_2
X_4384_ _5110_/Q _5078_/Q vssd1 vssd1 vccd1 vccd1 _4387_/A sky130_fd_sc_hd__nor2_1
X_3335_ _3335_/A _3335_/B vssd1 vssd1 vccd1 vccd1 _3339_/A sky130_fd_sc_hd__nor2_1
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3266_ _3266_/A _3266_/B vssd1 vssd1 vccd1 vccd1 _3267_/C sky130_fd_sc_hd__nand2_1
XFILLER_85_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5005_ _5097_/CLK hold39/X vssd1 vssd1 vccd1 vccd1 _5005_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_38_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3197_ _3197_/A _3197_/B vssd1 vssd1 vccd1 vccd1 _3198_/C sky130_fd_sc_hd__nor2_1
XFILLER_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120_ _3305_/B _3301_/A vssd1 vssd1 vccd1 vccd1 _3120_/X sky130_fd_sc_hd__or2_1
X_3051_ _3743_/B _5176_/Q vssd1 vssd1 vccd1 vccd1 _3052_/B sky130_fd_sc_hd__nand2_1
XFILLER_82_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3953_ _5100_/Q vssd1 vssd1 vccd1 vccd1 _4352_/A sky130_fd_sc_hd__inv_2
X_3884_ _4970_/X _3879_/X _3870_/X _3883_/Y vssd1 vssd1 vccd1 vccd1 _5125_/D sky130_fd_sc_hd__o211a_1
X_2904_ _3604_/A vssd1 vssd1 vccd1 vccd1 _3276_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_50_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2835_ _2836_/A _2836_/B _2836_/C vssd1 vssd1 vccd1 vccd1 _2835_/Y sky130_fd_sc_hd__a21oi_1
X_2766_ _2811_/A _2751_/Y _2765_/X vssd1 vssd1 vccd1 vccd1 _2853_/A sky130_fd_sc_hd__o21bai_2
X_2697_ _2997_/A _2997_/C _2997_/B vssd1 vssd1 vccd1 vccd1 _2989_/A sky130_fd_sc_hd__a21oi_4
X_4505_ _4506_/A _4507_/A _4506_/B _3879_/A vssd1 vssd1 vccd1 vccd1 _4505_/X sky130_fd_sc_hd__a31o_1
X_4436_ _4444_/A _4444_/C vssd1 vssd1 vccd1 vccd1 _4438_/B sky130_fd_sc_hd__and2_1
X_4367_ _4367_/A _4367_/B vssd1 vssd1 vccd1 vccd1 _4367_/Y sky130_fd_sc_hd__nand2_1
X_3318_ _3318_/A _3318_/B vssd1 vssd1 vccd1 vccd1 _3318_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4298_ _5085_/Q _5053_/Q vssd1 vssd1 vccd1 vccd1 _4576_/B sky130_fd_sc_hd__nand2_2
XFILLER_58_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3249_ _5244_/Q _2939_/X _3246_/X _3248_/X vssd1 vssd1 vccd1 vccd1 _5244_/D sky130_fd_sc_hd__o211a_1
XFILLER_54_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _5022_/Q vssd1 vssd1 vccd1 vccd1 _3000_/A sky130_fd_sc_hd__clkbuf_4
X_2551_ _2565_/A _4778_/B vssd1 vssd1 vccd1 vccd1 _2551_/Y sky130_fd_sc_hd__nand2_1
X_5270_ _5288_/CLK _5270_/D vssd1 vssd1 vccd1 vccd1 _5270_/Q sky130_fd_sc_hd__dfxtp_1
X_4221_ _4226_/B _4221_/B vssd1 vssd1 vccd1 vccd1 _4221_/Y sky130_fd_sc_hd__nand2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_68_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4152_ _5101_/Q _5100_/Q _5099_/Q vssd1 vssd1 vccd1 vccd1 _4152_/X sky130_fd_sc_hd__and3_1
X_3103_ _3103_/A _3103_/B vssd1 vssd1 vccd1 vccd1 _3325_/A sky130_fd_sc_hd__or2_1
X_4083_ _4164_/A _5098_/Q _5097_/Q vssd1 vssd1 vccd1 vccd1 _4087_/B sky130_fd_sc_hd__and3_1
XFILLER_83_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3034_ _3175_/A vssd1 vssd1 vccd1 vccd1 _3034_/Y sky130_fd_sc_hd__inv_2
XFILLER_36_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4985_ _4987_/CLK hold43/X vssd1 vssd1 vccd1 vccd1 _4986_/D sky130_fd_sc_hd__dfxtp_1
X_3936_ _3934_/B _5010_/Q _5122_/Q _3935_/Y vssd1 vssd1 vccd1 vccd1 _3936_/X sky130_fd_sc_hd__a22o_1
X_3867_ _5130_/Q _3862_/X _3857_/X _3866_/Y vssd1 vssd1 vccd1 vccd1 _5130_/D sky130_fd_sc_hd__o211a_1
X_2818_ _2787_/B _2787_/A _2826_/B _2826_/C vssd1 vssd1 vccd1 vccd1 _2818_/Y sky130_fd_sc_hd__a22oi_1
X_3798_ _3807_/A _3798_/B vssd1 vssd1 vccd1 vccd1 _3798_/Y sky130_fd_sc_hd__nand2_1
XFILLER_11_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2749_ _2926_/B _2749_/B vssd1 vssd1 vccd1 vccd1 _2930_/B sky130_fd_sc_hd__nand2_1
XFILLER_11_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4419_ _4415_/Y _4418_/X _2869_/X vssd1 vssd1 vccd1 vccd1 _5081_/D sky130_fd_sc_hd__o21a_1
Xinput19 phase_in[6] vssd1 vssd1 vccd1 vccd1 hold41/A sky130_fd_sc_hd__clkbuf_1
XFILLER_52_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4770_ _4770_/A vssd1 vssd1 vccd1 vccd1 _4770_/X sky130_fd_sc_hd__clkbuf_2
X_3721_ _3726_/A _3721_/B vssd1 vssd1 vccd1 vccd1 _3721_/Y sky130_fd_sc_hd__nand2_1
X_3652_ _3652_/A _3652_/B vssd1 vssd1 vccd1 vccd1 _3658_/A sky130_fd_sc_hd__and2_1
X_2603_ _5294_/Q _2586_/X _2600_/X _2602_/Y vssd1 vssd1 vccd1 vccd1 _5294_/D sky130_fd_sc_hd__o211a_1
X_3583_ _5213_/Q _3705_/A _2889_/X vssd1 vssd1 vccd1 vccd1 _3583_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2534_ _5045_/Q vssd1 vssd1 vccd1 vccd1 _4710_/A sky130_fd_sc_hd__inv_2
X_5253_ _5285_/CLK _5253_/D vssd1 vssd1 vccd1 vccd1 _5253_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_87_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5184_ _5247_/CLK _5184_/D vssd1 vssd1 vccd1 vccd1 _5184_/Q sky130_fd_sc_hd__dfxtp_1
X_4204_ _4764_/A vssd1 vssd1 vccd1 vccd1 _4204_/X sky130_fd_sc_hd__buf_2
X_4135_ _5106_/Q vssd1 vssd1 vccd1 vccd1 _4250_/A sky130_fd_sc_hd__inv_2
XFILLER_28_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_83_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4066_ _4580_/A _4062_/X _4234_/B _4220_/A vssd1 vssd1 vccd1 vccd1 _4067_/C sky130_fd_sc_hd__o211ai_4
X_3017_ _4631_/A _3017_/B vssd1 vssd1 vccd1 vccd1 _3017_/Y sky130_fd_sc_hd__nor2_1
XPHY_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4968_ _4968_/A _4968_/B vssd1 vssd1 vccd1 vccd1 _4968_/Y sky130_fd_sc_hd__nand2_1
XFILLER_51_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3919_ _5116_/Q vssd1 vssd1 vccd1 vccd1 _3920_/A sky130_fd_sc_hd__inv_2
X_4899_ _4896_/Y _4899_/B _4899_/C vssd1 vssd1 vccd1 vccd1 _5016_/D sky130_fd_sc_hd__and3b_1
XFILLER_3_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_80_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4822_ _4827_/B _4827_/A vssd1 vssd1 vccd1 vccd1 _4823_/A sky130_fd_sc_hd__nand2_1
XFILLER_33_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4753_ _4757_/B _4757_/A vssd1 vssd1 vccd1 vccd1 _4758_/B sky130_fd_sc_hd__nor2_1
X_3704_ _5126_/Q _3875_/B vssd1 vssd1 vccd1 vccd1 _3704_/Y sky130_fd_sc_hd__nor2_1
X_4684_ _4684_/A vssd1 vssd1 vccd1 vccd1 _4686_/A sky130_fd_sc_hd__inv_2
X_3635_ _3635_/A _3635_/B vssd1 vssd1 vccd1 vccd1 _3635_/Y sky130_fd_sc_hd__nand2_1
X_3566_ _3566_/A _3566_/B vssd1 vssd1 vccd1 vccd1 _3569_/A sky130_fd_sc_hd__nor2_1
X_3497_ _3511_/A vssd1 vssd1 vccd1 vccd1 _3582_/C sky130_fd_sc_hd__inv_2
X_2517_ _5048_/Q vssd1 vssd1 vccd1 vccd1 _4725_/A sky130_fd_sc_hd__inv_2
X_5305_ _5311_/CLK _5305_/D vssd1 vssd1 vccd1 vccd1 _5305_/Q sky130_fd_sc_hd__dfxtp_1
X_5236_ _5236_/CLK _5236_/D vssd1 vssd1 vccd1 vccd1 _5236_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_75_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5167_ _5171_/CLK _5167_/D vssd1 vssd1 vccd1 vccd1 _5167_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4118_ _4118_/A vssd1 vssd1 vccd1 vccd1 _4119_/B sky130_fd_sc_hd__inv_2
X_5098_ _5098_/CLK _5098_/D vssd1 vssd1 vccd1 vccd1 _5098_/Q sky130_fd_sc_hd__dfxtp_1
X_4049_ _4018_/X _4048_/Y _4064_/A _4063_/A _4059_/B vssd1 vssd1 vccd1 vccd1 _4052_/A
+ sky130_fd_sc_hd__o2111ai_4
XFILLER_17_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_83_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold8 phase_in[3] vssd1 vssd1 vccd1 vccd1 hold8/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_87_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3420_ _3420_/A _3455_/A vssd1 vssd1 vccd1 vccd1 _3638_/A sky130_fd_sc_hd__nand2_1
X_3351_ _3351_/A _3359_/B vssd1 vssd1 vccd1 vccd1 _3352_/A sky130_fd_sc_hd__and2_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3282_ _3281_/B _3281_/A _2969_/X vssd1 vssd1 vccd1 vccd1 _3282_/X sky130_fd_sc_hd__a21o_1
XFILLER_85_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5021_ _5027_/CLK _5021_/D vssd1 vssd1 vccd1 vccd1 _5021_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_80_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4805_ _5036_/Q _4770_/X _4803_/Y _4804_/X _4785_/X vssd1 vssd1 vccd1 vccd1 _5036_/D
+ sky130_fd_sc_hd__o221a_1
X_2997_ _2997_/A _2997_/B _2997_/C vssd1 vssd1 vccd1 vccd1 _2997_/X sky130_fd_sc_hd__and3_1
X_4736_ _4798_/A _4736_/B _4736_/C vssd1 vssd1 vccd1 vccd1 _4736_/X sky130_fd_sc_hd__or3_2
X_4667_ _4667_/A _4667_/B vssd1 vssd1 vccd1 vccd1 _4820_/A sky130_fd_sc_hd__nor2_1
X_3618_ _3618_/A _3618_/B vssd1 vssd1 vccd1 vccd1 _3625_/A sky130_fd_sc_hd__nor2_1
X_4598_ _4606_/A _4598_/B vssd1 vssd1 vccd1 vccd1 _4599_/A sky130_fd_sc_hd__nor2_1
XFILLER_88_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3549_ _5250_/Q _3549_/B vssd1 vssd1 vccd1 vccd1 _3550_/B sky130_fd_sc_hd__nor2_1
XFILLER_88_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_76_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5219_ _5219_/CLK _5219_/D vssd1 vssd1 vccd1 vccd1 _5219_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2920_ _2911_/Y _2910_/Y _2909_/X _2919_/Y vssd1 vssd1 vccd1 vccd1 _2920_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2851_ _4785_/A vssd1 vssd1 vccd1 vccd1 _4902_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_79_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2782_ _5315_/Q vssd1 vssd1 vccd1 vccd1 _2783_/B sky130_fd_sc_hd__inv_2
XPHY_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4521_ _4519_/Y _4520_/X _4475_/X vssd1 vssd1 vccd1 vccd1 _4521_/Y sky130_fd_sc_hd__o21ai_1
X_4452_ _4420_/X _5076_/Q _4450_/Y _4451_/X _4432_/X vssd1 vssd1 vccd1 vccd1 _5076_/D
+ sky130_fd_sc_hd__o221a_1
X_3403_ _5143_/Q _3831_/B vssd1 vssd1 vccd1 vccd1 _3608_/A sky130_fd_sc_hd__nor2_2
X_4383_ _4383_/A _4383_/B vssd1 vssd1 vccd1 vccd1 _4444_/B sky130_fd_sc_hd__nand2_2
X_3334_ _5163_/Q _3779_/B vssd1 vssd1 vccd1 vccd1 _3335_/B sky130_fd_sc_hd__nor2_1
XFILLER_58_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3265_ _3828_/B _4968_/A vssd1 vssd1 vccd1 vccd1 _3265_/Y sky130_fd_sc_hd__nor2_1
X_5004_ _5114_/CLK _5004_/D vssd1 vssd1 vccd1 vccd1 _5004_/Q sky130_fd_sc_hd__dfxtp_1
X_3196_ _3180_/Y _3183_/Y _3204_/B vssd1 vssd1 vccd1 vccd1 _3198_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4719_ _4705_/B _4700_/A _4705_/A vssd1 vssd1 vccd1 vccd1 _4719_/X sky130_fd_sc_hd__o21ba_1
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_72_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3050_ _5176_/Q _3743_/B vssd1 vssd1 vccd1 vccd1 _3064_/B sky130_fd_sc_hd__or2_2
XFILLER_48_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3952_ _5101_/Q vssd1 vssd1 vccd1 vccd1 _4342_/A sky130_fd_sc_hd__inv_2
X_3883_ _3933_/B _4846_/B vssd1 vssd1 vccd1 vccd1 _3883_/Y sky130_fd_sc_hd__nand2_1
X_2903_ _2902_/X _2903_/B vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__and2b_1
X_2834_ _2834_/A _2834_/B vssd1 vssd1 vccd1 vccd1 _2836_/C sky130_fd_sc_hd__nor2_1
XFILLER_31_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4504_ _4504_/A _4504_/B vssd1 vssd1 vccd1 vccd1 _4507_/A sky130_fd_sc_hd__nor2_1
X_2765_ _2902_/C _2769_/B _2764_/X vssd1 vssd1 vccd1 vccd1 _2765_/X sky130_fd_sc_hd__or3b_1
X_2696_ _2993_/B _2696_/B vssd1 vssd1 vccd1 vccd1 _2997_/B sky130_fd_sc_hd__nand2_2
X_4435_ _4454_/A _4454_/B _4390_/A vssd1 vssd1 vccd1 vccd1 _4444_/A sky130_fd_sc_hd__o21ai_1
X_4366_ _4470_/B _4457_/A _4457_/B vssd1 vssd1 vccd1 vccd1 _4367_/B sky130_fd_sc_hd__and3_1
X_3317_ _5231_/Q _3269_/X _3313_/Y _3314_/X _3316_/X vssd1 vssd1 vccd1 vccd1 _5231_/D
+ sky130_fd_sc_hd__o221a_1
X_4297_ _5086_/Q _5054_/Q vssd1 vssd1 vccd1 vccd1 _4571_/B sky130_fd_sc_hd__nand2_2
XFILLER_58_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3248_ _3243_/A _3247_/Y _2963_/X vssd1 vssd1 vccd1 vccd1 _3248_/X sky130_fd_sc_hd__a21o_1
XFILLER_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3179_ _3231_/A _3231_/C _3178_/X vssd1 vssd1 vccd1 vccd1 _3179_/Y sky130_fd_sc_hd__a21oi_4
XFILLER_54_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_82_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_72_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _5041_/Q vssd1 vssd1 vccd1 vccd1 _4778_/B sky130_fd_sc_hd__inv_2
X_4220_ _4220_/A _4234_/B vssd1 vssd1 vccd1 vccd1 _4221_/B sky130_fd_sc_hd__nand2_1
X_4151_ _4365_/A _4154_/A _4150_/Y vssd1 vssd1 vccd1 vccd1 _5103_/D sky130_fd_sc_hd__a21oi_1
XFILLER_83_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3102_ _3773_/B _5165_/Q vssd1 vssd1 vccd1 vccd1 _3103_/B sky130_fd_sc_hd__and2_1
X_4082_ _4331_/A _4326_/A vssd1 vssd1 vccd1 vccd1 _4164_/A sky130_fd_sc_hd__nor2_2
XFILLER_83_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3033_ _5183_/Q _3724_/B vssd1 vssd1 vccd1 vccd1 _3175_/A sky130_fd_sc_hd__nor2_1
XFILLER_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4984_ _5002_/CLK _4984_/D vssd1 vssd1 vccd1 vccd1 _4984_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_23_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3935_ _5012_/Q vssd1 vssd1 vccd1 vccd1 _3935_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3866_ _3873_/A _3866_/B vssd1 vssd1 vccd1 vccd1 _3866_/Y sky130_fd_sc_hd__nand2_1
X_3797_ _3823_/A vssd1 vssd1 vccd1 vccd1 _3807_/A sky130_fd_sc_hd__clkbuf_2
X_2817_ _2834_/A vssd1 vssd1 vccd1 vccd1 _2826_/C sky130_fd_sc_hd__inv_2
XFILLER_11_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2748_ _4808_/A _5302_/Q vssd1 vssd1 vccd1 vccd1 _2749_/B sky130_fd_sc_hd__nand2_1
X_4418_ _4423_/A _4416_/Y _4742_/B _4411_/B vssd1 vssd1 vccd1 vccd1 _4418_/X sky130_fd_sc_hd__o211a_1
X_2679_ _2728_/B _2729_/A _5031_/Q _2678_/Y vssd1 vssd1 vccd1 vccd1 _2808_/A sky130_fd_sc_hd__a31o_1
X_4349_ _4487_/A _4478_/A vssd1 vssd1 vccd1 vccd1 _4359_/A sky130_fd_sc_hd__nand2_1
XFILLER_27_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3720_ _5185_/Q _3715_/X _3710_/X _3719_/Y vssd1 vssd1 vccd1 vccd1 _5185_/D sky130_fd_sc_hd__o211a_1
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_40_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5311_/CLK sky130_fd_sc_hd__clkbuf_16
X_3651_ _3651_/A vssd1 vssd1 vccd1 vccd1 _3655_/A sky130_fd_sc_hd__inv_2
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2602_ _2602_/A _4846_/A vssd1 vssd1 vccd1 vccd1 _2602_/Y sky130_fd_sc_hd__nand2_1
X_3582_ _3504_/B _3582_/B _3582_/C vssd1 vssd1 vccd1 vccd1 _3582_/Y sky130_fd_sc_hd__nand3b_1
X_2533_ _5313_/Q _2528_/X _2522_/X _2532_/Y vssd1 vssd1 vccd1 vccd1 _5313_/D sky130_fd_sc_hd__o211a_1
XFILLER_87_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5252_ _5252_/CLK _5252_/D vssd1 vssd1 vccd1 vccd1 _5252_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4203_ _4286_/A _4206_/A _4202_/X vssd1 vssd1 vccd1 vccd1 _5088_/D sky130_fd_sc_hd__a21oi_1
X_5183_ _5247_/CLK _5183_/D vssd1 vssd1 vccd1 vccd1 _5183_/Q sky130_fd_sc_hd__dfxtp_1
X_4134_ _4370_/A _4139_/A _4133_/Y vssd1 vssd1 vccd1 vccd1 _5107_/D sky130_fd_sc_hd__a21oi_1
XFILLER_28_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4065_ _4233_/A _4233_/B _5083_/Q vssd1 vssd1 vccd1 vccd1 _4220_/A sky130_fd_sc_hd__a21boi_4
XFILLER_83_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3016_ _3022_/B _5286_/Q vssd1 vssd1 vccd1 vccd1 _3023_/B sky130_fd_sc_hd__nand2_1
XPHY_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4967_ _5003_/Q _5004_/Q vssd1 vssd1 vccd1 vccd1 _4967_/X sky130_fd_sc_hd__and2_1
X_3918_ _4440_/A vssd1 vssd1 vccd1 vccd1 _4446_/A sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_31_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5219_/CLK sky130_fd_sc_hd__clkbuf_16
X_4898_ _4898_/A _4898_/B vssd1 vssd1 vccd1 vccd1 _4899_/C sky130_fd_sc_hd__nand2_1
XFILLER_22_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3849_ _3862_/A vssd1 vssd1 vccd1 vccd1 _3849_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_59_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 _5171_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_6_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4821_ _4821_/A _4821_/B vssd1 vssd1 vccd1 vccd1 _4827_/B sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_13_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5125_/CLK sky130_fd_sc_hd__clkbuf_16
X_4752_ _4757_/B _4757_/A _4715_/A _4720_/B vssd1 vssd1 vccd1 vccd1 _4752_/X sky130_fd_sc_hd__o211a_1
X_3703_ _5191_/Q _2524_/A _3701_/Y _3702_/X _3695_/X vssd1 vssd1 vccd1 vccd1 _5191_/D
+ sky130_fd_sc_hd__o221a_1
X_4683_ _4683_/A _4685_/B vssd1 vssd1 vccd1 vccd1 _4684_/A sky130_fd_sc_hd__nor2_1
X_3634_ _5203_/Q _3596_/X _3632_/Y _3633_/X _3591_/X vssd1 vssd1 vccd1 vccd1 _5203_/D
+ sky130_fd_sc_hd__o221a_1
X_3565_ _3563_/Y _3564_/Y _3202_/X vssd1 vssd1 vccd1 vccd1 _5216_/D sky130_fd_sc_hd__a21oi_1
X_3496_ _5148_/Q _3818_/B vssd1 vssd1 vccd1 vccd1 _3511_/A sky130_fd_sc_hd__nor2_1
X_2516_ _5316_/Q _2506_/X _2510_/X _2515_/Y vssd1 vssd1 vccd1 vccd1 _5316_/D sky130_fd_sc_hd__o211a_1
X_5304_ _5311_/CLK _5304_/D vssd1 vssd1 vccd1 vccd1 _5304_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_88_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5235_ _5268_/CLK _5235_/D vssd1 vssd1 vccd1 vccd1 _5235_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_56_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_5166_ _5288_/CLK _5166_/D vssd1 vssd1 vccd1 vccd1 _5166_/Q sky130_fd_sc_hd__dfxtp_1
X_4117_ _4131_/B _5108_/Q _5107_/Q vssd1 vssd1 vccd1 vccd1 _4118_/A sky130_fd_sc_hd__and3_1
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5097_ _5097_/CLK _5097_/D vssd1 vssd1 vccd1 vccd1 _5097_/Q sky130_fd_sc_hd__dfxtp_1
X_4048_ _4056_/C _4048_/B vssd1 vssd1 vccd1 vccd1 _4048_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold9 hold9/A vssd1 vssd1 vccd1 vccd1 hold9/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_58_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3350_ _3787_/B _5160_/Q vssd1 vssd1 vccd1 vccd1 _3350_/X sky130_fd_sc_hd__and2_1
X_5020_ _5301_/CLK _5020_/D vssd1 vssd1 vccd1 vccd1 _5020_/Q sky130_fd_sc_hd__dfxtp_1
X_3281_ _3281_/A _3281_/B vssd1 vssd1 vccd1 vccd1 _3281_/Y sky130_fd_sc_hd__nor2_1
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_2_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5098_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_65_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_80_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4804_ _4803_/B _4803_/A _4764_/X vssd1 vssd1 vccd1 vccd1 _4804_/X sky130_fd_sc_hd__a21o_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4735_ _4735_/A _4735_/B _4735_/C vssd1 vssd1 vccd1 vccd1 _4736_/C sky130_fd_sc_hd__and3_1
XFILLER_21_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2996_ _2634_/X _2992_/Y _2993_/X _2915_/X _2995_/Y vssd1 vssd1 vccd1 vccd1 _5259_/D
+ sky130_fd_sc_hd__o311a_1
X_4666_ _4666_/A _4666_/B vssd1 vssd1 vccd1 vccd1 _4667_/B sky130_fd_sc_hd__nor2_1
X_3617_ _5206_/Q _3613_/X _3585_/X _3616_/X vssd1 vssd1 vccd1 vccd1 _5206_/D sky130_fd_sc_hd__o211a_1
X_4597_ _4597_/A _4597_/B vssd1 vssd1 vccd1 vccd1 _4598_/B sky130_fd_sc_hd__nor2_2
X_3548_ _5219_/Q _3365_/X _3546_/Y _3547_/X _3363_/X vssd1 vssd1 vccd1 vccd1 _5219_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_76_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3479_ _5140_/Q _3839_/B vssd1 vssd1 vccd1 vccd1 _3622_/B sky130_fd_sc_hd__or2_2
X_5218_ _5219_/CLK _5218_/D vssd1 vssd1 vccd1 vccd1 _5218_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_69_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5149_ _5221_/CLK _5149_/D vssd1 vssd1 vccd1 vccd1 _5149_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_71_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_90_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2850_ _3315_/A vssd1 vssd1 vccd1 vccd1 _4785_/A sky130_fd_sc_hd__buf_1
XPHY_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2781_ _5048_/Q vssd1 vssd1 vccd1 vccd1 _4739_/A sky130_fd_sc_hd__clkbuf_2
XPHY_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4520_ _4520_/A _4520_/B vssd1 vssd1 vccd1 vccd1 _4520_/X sky130_fd_sc_hd__and2_1
X_4451_ _4450_/B _4450_/A _4588_/A vssd1 vssd1 vccd1 vccd1 _4451_/X sky130_fd_sc_hd__a21o_1
X_3402_ _3831_/B _5143_/Q vssd1 vssd1 vccd1 vccd1 _3608_/B sky130_fd_sc_hd__and2_2
X_4382_ _4382_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4383_/B sky130_fd_sc_hd__nand2_1
X_3333_ _3333_/A vssd1 vssd1 vccd1 vccd1 _3337_/A sky130_fd_sc_hd__inv_2
X_3264_ _5240_/Q vssd1 vssd1 vccd1 vccd1 _3828_/B sky130_fd_sc_hd__inv_2
X_5003_ _5114_/CLK _5003_/D vssd1 vssd1 vccd1 vccd1 _5003_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3195_ _5283_/Q _3195_/B vssd1 vssd1 vccd1 vccd1 _3204_/B sky130_fd_sc_hd__nor2_1
XFILLER_81_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2979_ _2979_/A _2979_/B vssd1 vssd1 vccd1 vccd1 _2980_/A sky130_fd_sc_hd__nor2_1
X_4718_ _4767_/A _4767_/B _4717_/Y vssd1 vssd1 vccd1 vccd1 _4746_/A sky130_fd_sc_hd__o21bai_1
X_4649_ _5027_/Q _5059_/Q vssd1 vssd1 vccd1 vccd1 _4650_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_72_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_71_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_67_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3951_ _5102_/Q vssd1 vssd1 vccd1 vccd1 _4347_/A sky130_fd_sc_hd__inv_2
X_2902_ _2902_/A _2902_/B _2902_/C vssd1 vssd1 vccd1 vccd1 _2902_/X sky130_fd_sc_hd__and3_1
XFILLER_50_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3882_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4846_/B sky130_fd_sc_hd__buf_2
X_2833_ _2827_/Y _2829_/Y _4913_/A vssd1 vssd1 vccd1 vccd1 _5284_/D sky130_fd_sc_hd__a21oi_1
X_2764_ _2762_/Y _2764_/B vssd1 vssd1 vccd1 vccd1 _2764_/X sky130_fd_sc_hd__and2b_1
X_4503_ _4510_/B _4510_/A vssd1 vssd1 vccd1 vccd1 _4506_/A sky130_fd_sc_hd__or2_1
X_2695_ _4628_/A _5290_/Q vssd1 vssd1 vccd1 vccd1 _2696_/B sky130_fd_sc_hd__nand2_1
XFILLER_6_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4434_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4434_/X sky130_fd_sc_hd__buf_2
X_4365_ _4365_/A _4602_/B vssd1 vssd1 vccd1 vccd1 _4457_/B sky130_fd_sc_hd__nand2_1
X_3316_ _3695_/A vssd1 vssd1 vccd1 vccd1 _3316_/X sky130_fd_sc_hd__clkbuf_2
X_4296_ _4581_/B _4575_/B _4576_/A vssd1 vssd1 vccd1 vccd1 _4568_/A sky130_fd_sc_hd__o21ai_2
X_3247_ _3247_/A _3247_/B vssd1 vssd1 vccd1 vccd1 _3247_/Y sky130_fd_sc_hd__nand2_1
X_3178_ _3178_/A _3218_/A vssd1 vssd1 vccd1 vccd1 _3178_/X sky130_fd_sc_hd__or2_2
XFILLER_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_66_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4150_ _4150_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4150_/Y sky130_fd_sc_hd__nand2_1
X_3101_ _5165_/Q _3773_/B vssd1 vssd1 vccd1 vccd1 _3103_/A sky130_fd_sc_hd__nor2_1
X_4081_ _5095_/Q vssd1 vssd1 vccd1 vccd1 _4326_/A sky130_fd_sc_hd__inv_2
X_3032_ _5279_/Q vssd1 vssd1 vccd1 vccd1 _3724_/B sky130_fd_sc_hd__inv_2
X_4983_ _4992_/CLK hold21/X vssd1 vssd1 vccd1 vccd1 _4984_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3934_ _5010_/Q _3934_/B vssd1 vssd1 vccd1 vccd1 _3934_/Y sky130_fd_sc_hd__nor2_1
X_3865_ _5131_/Q _3862_/X _3857_/X _3864_/Y vssd1 vssd1 vccd1 vccd1 _5131_/D sky130_fd_sc_hd__o211a_1
X_2816_ _2783_/B _4739_/A _2843_/A _2815_/Y vssd1 vssd1 vccd1 vccd1 _2826_/B sky130_fd_sc_hd__o22ai_2
X_3796_ _3822_/A vssd1 vssd1 vccd1 vccd1 _3796_/X sky130_fd_sc_hd__clkbuf_2
X_2747_ _2747_/A _2747_/B vssd1 vssd1 vccd1 vccd1 _2927_/A sky130_fd_sc_hd__or2_1
X_2678_ _5299_/Q _4666_/A vssd1 vssd1 vccd1 vccd1 _2678_/Y sky130_fd_sc_hd__nor2_1
X_4417_ _4417_/A vssd1 vssd1 vccd1 vccd1 _4742_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_59_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4348_ _4362_/B _4348_/B vssd1 vssd1 vccd1 vccd1 _4478_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4279_ _5090_/Q _5058_/Q vssd1 vssd1 vccd1 vccd1 _4306_/A sky130_fd_sc_hd__nor2_1
XFILLER_27_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3650_ _3650_/A vssd1 vssd1 vccd1 vccd1 _3650_/X sky130_fd_sc_hd__clkbuf_2
X_2601_ _5027_/Q vssd1 vssd1 vccd1 vccd1 _4846_/A sky130_fd_sc_hd__inv_2
X_3581_ _3582_/B _3582_/C _3504_/B vssd1 vssd1 vccd1 vccd1 _3581_/X sky130_fd_sc_hd__a21bo_1
X_2532_ _2546_/A _4755_/A vssd1 vssd1 vccd1 vccd1 _2532_/Y sky130_fd_sc_hd__nand2_1
X_5251_ _5251_/CLK _5251_/D vssd1 vssd1 vccd1 vccd1 _5251_/Q sky130_fd_sc_hd__dfxtp_1
X_4202_ _4589_/A _4202_/B vssd1 vssd1 vccd1 vccd1 _4202_/X sky130_fd_sc_hd__or2_1
XFILLER_68_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5182_ _5247_/CLK _5182_/D vssd1 vssd1 vccd1 vccd1 _5182_/Q sky130_fd_sc_hd__dfxtp_1
X_4133_ _4133_/A _4183_/B vssd1 vssd1 vccd1 vccd1 _4133_/Y sky130_fd_sc_hd__nand2_1
X_4064_ _4064_/A vssd1 vssd1 vccd1 vccd1 _4233_/B sky130_fd_sc_hd__inv_2
X_3015_ _3789_/B _4968_/A vssd1 vssd1 vccd1 vccd1 _3015_/Y sky130_fd_sc_hd__nor2_1
XFILLER_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4966_ _4966_/A _4966_/B vssd1 vssd1 vccd1 vccd1 _4966_/X sky130_fd_sc_hd__and2_1
XFILLER_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3917_ _3907_/X _4978_/X _3911_/X _3916_/Y vssd1 vssd1 vccd1 vccd1 _5117_/D sky130_fd_sc_hd__o211a_1
X_4897_ _5017_/Q _4896_/Y _4891_/A _4899_/B vssd1 vssd1 vccd1 vccd1 _5017_/D sky130_fd_sc_hd__o211a_1
X_3848_ _5137_/Q _3835_/X _3844_/X _3847_/Y vssd1 vssd1 vccd1 vccd1 _5137_/D sky130_fd_sc_hd__o211a_1
XFILLER_22_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3779_ _3781_/A _3779_/B vssd1 vssd1 vccd1 vccd1 _3779_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_86_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_80_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_73_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4820_ _4820_/A vssd1 vssd1 vccd1 vccd1 _4824_/A sky130_fd_sc_hd__inv_2
XFILLER_21_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4751_ _4750_/X _4717_/A _4719_/X vssd1 vssd1 vccd1 vccd1 _4757_/A sky130_fd_sc_hd__a21oi_2
X_3702_ _3705_/B _3701_/B _3642_/X vssd1 vssd1 vccd1 vccd1 _3702_/X sky130_fd_sc_hd__a21o_1
X_4682_ _4682_/A _4682_/B vssd1 vssd1 vccd1 vccd1 _4801_/B sky130_fd_sc_hd__nor2_1
X_3633_ _3632_/B _3632_/A _3361_/X vssd1 vssd1 vccd1 vccd1 _3633_/X sky130_fd_sc_hd__a21o_1
X_3564_ _3605_/A _5216_/Q vssd1 vssd1 vccd1 vccd1 _3564_/Y sky130_fd_sc_hd__nand2_1
X_3495_ _5244_/Q vssd1 vssd1 vccd1 vccd1 _3818_/B sky130_fd_sc_hd__inv_2
X_2515_ _2524_/A _4591_/A vssd1 vssd1 vccd1 vccd1 _2515_/Y sky130_fd_sc_hd__nand2_1
X_5303_ _5303_/CLK _5303_/D vssd1 vssd1 vccd1 vccd1 _5303_/Q sky130_fd_sc_hd__dfxtp_1
X_5234_ _5251_/CLK _5234_/D vssd1 vssd1 vccd1 vccd1 _5234_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5165_ _5288_/CLK _5165_/D vssd1 vssd1 vccd1 vccd1 _5165_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4116_ _4116_/A _4116_/B _4116_/C vssd1 vssd1 vccd1 vccd1 _5111_/D sky130_fd_sc_hd__nor3_1
XFILLER_68_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5096_ _5096_/CLK _5096_/D vssd1 vssd1 vccd1 vccd1 _5096_/Q sky130_fd_sc_hd__dfxtp_1
X_4047_ _4047_/A _4051_/B _4059_/B vssd1 vssd1 vccd1 vccd1 _4070_/A sky130_fd_sc_hd__nand3_4
XFILLER_37_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4949_ _5121_/Q _4949_/B vssd1 vssd1 vccd1 vccd1 _4950_/B sky130_fd_sc_hd__nor2_1
XFILLER_33_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_74_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3280_ _3752_/B _5172_/Q _3279_/X vssd1 vssd1 vccd1 vccd1 _3281_/B sky130_fd_sc_hd__o21a_1
XFILLER_65_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4803_ _4803_/A _4803_/B vssd1 vssd1 vccd1 vccd1 _4803_/Y sky130_fd_sc_hd__nor2_1
XFILLER_61_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4734_ _4734_/A _4734_/B _4734_/C vssd1 vssd1 vccd1 vccd1 _5050_/D sky130_fd_sc_hd__nor3_1
X_2995_ _2995_/A _3779_/B vssd1 vssd1 vccd1 vccd1 _2995_/Y sky130_fd_sc_hd__nand2_1
X_4665_ _5032_/Q _5064_/Q vssd1 vssd1 vccd1 vccd1 _4667_/A sky130_fd_sc_hd__nor2_1
X_3616_ _3610_/A _3614_/Y _3615_/X vssd1 vssd1 vccd1 vccd1 _3616_/X sky130_fd_sc_hd__a21o_1
X_4596_ _5042_/Q _5074_/Q vssd1 vssd1 vccd1 vccd1 _4606_/A sky130_fd_sc_hd__nor2_1
X_3547_ _3521_/Y _3524_/Y _3545_/Y _3206_/X vssd1 vssd1 vccd1 vccd1 _3547_/X sky130_fd_sc_hd__a31o_1
XFILLER_88_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_88_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3478_ _5236_/Q vssd1 vssd1 vccd1 vccd1 _3839_/B sky130_fd_sc_hd__inv_2
X_5217_ _5221_/CLK _5217_/D vssd1 vssd1 vccd1 vccd1 _5217_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_5148_ _5236_/CLK _5148_/D vssd1 vssd1 vccd1 vccd1 _5148_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5079_ _5108_/CLK _5079_/D vssd1 vssd1 vccd1 vccd1 _5079_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2780_ _2843_/A vssd1 vssd1 vccd1 vccd1 _2836_/B sky130_fd_sc_hd__inv_2
XPHY_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4450_ _4450_/A _4450_/B vssd1 vssd1 vccd1 vccd1 _4450_/Y sky130_fd_sc_hd__nor2_1
X_3401_ _5239_/Q vssd1 vssd1 vccd1 vccd1 _3831_/B sky130_fd_sc_hd__inv_2
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4381_ _4381_/A vssd1 vssd1 vccd1 vccd1 _4383_/A sky130_fd_sc_hd__inv_2
X_3332_ _5228_/Q _3328_/X _3304_/X _3331_/X vssd1 vssd1 vccd1 vccd1 _5228_/D sky130_fd_sc_hd__o211a_1
X_3263_ _5241_/Q _3210_/X _3260_/Y _3261_/X _3262_/X vssd1 vssd1 vccd1 vccd1 _5241_/D
+ sky130_fd_sc_hd__o221a_1
X_5002_ _5002_/CLK _5002_/D vssd1 vssd1 vccd1 vccd1 _5002_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_66_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3194_ _5187_/Q vssd1 vssd1 vccd1 vccd1 _3195_/B sky130_fd_sc_hd__inv_2
XFILLER_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_81_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2978_ _2978_/A vssd1 vssd1 vccd1 vccd1 _2979_/B sky130_fd_sc_hd__inv_2
X_4717_ _4717_/A _4717_/B vssd1 vssd1 vccd1 vccd1 _4717_/Y sky130_fd_sc_hd__nand2_1
X_4648_ _4846_/A _4648_/B vssd1 vssd1 vccd1 vccd1 _4650_/A sky130_fd_sc_hd__nand2_1
XFILLER_89_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4579_ _4574_/X _5053_/Q _4577_/Y _4578_/X _4508_/X vssd1 vssd1 vccd1 vccd1 _5053_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_76_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_84_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3950_ _4386_/A _4382_/A _4375_/A _4370_/A vssd1 vssd1 vccd1 vccd1 _4100_/C sky130_fd_sc_hd__or4_4
XFILLER_35_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2901_ _2901_/A vssd1 vssd1 vccd1 vccd1 _2901_/X sky130_fd_sc_hd__clkbuf_2
X_3881_ _4893_/A vssd1 vssd1 vccd1 vccd1 _4814_/A sky130_fd_sc_hd__buf_1
X_2832_ _4169_/A vssd1 vssd1 vccd1 vccd1 _4913_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_31_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2763_ _4601_/A _5307_/Q vssd1 vssd1 vccd1 vccd1 _2764_/B sky130_fd_sc_hd__nand2_1
X_4502_ _4502_/A _4502_/B vssd1 vssd1 vccd1 vccd1 _4510_/A sky130_fd_sc_hd__and2_1
X_2694_ _3000_/B _3000_/A vssd1 vssd1 vccd1 vccd1 _2997_/C sky130_fd_sc_hd__nand2_2
X_4433_ _4420_/X _5079_/Q _4430_/X _4431_/Y _4432_/X vssd1 vssd1 vccd1 vccd1 _5079_/D
+ sky130_fd_sc_hd__o221a_1
X_4364_ _4364_/A _4364_/B vssd1 vssd1 vccd1 vccd1 _4470_/B sky130_fd_sc_hd__nor2_2
X_4295_ _5085_/Q _5053_/Q vssd1 vssd1 vccd1 vccd1 _4576_/A sky130_fd_sc_hd__or2_1
X_3315_ _3315_/A vssd1 vssd1 vccd1 vccd1 _3695_/A sky130_fd_sc_hd__buf_2
X_3246_ _3646_/A vssd1 vssd1 vccd1 vccd1 _3246_/X sky130_fd_sc_hd__clkbuf_2
X_3177_ _3231_/B _3177_/B vssd1 vssd1 vccd1 vccd1 _3218_/A sky130_fd_sc_hd__or2_1
XFILLER_39_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3100_ _5261_/Q vssd1 vssd1 vccd1 vccd1 _3773_/B sky130_fd_sc_hd__inv_2
X_4080_ _5096_/Q vssd1 vssd1 vccd1 vccd1 _4331_/A sky130_fd_sc_hd__inv_2
X_3031_ _5186_/Q vssd1 vssd1 vccd1 vccd1 _3211_/B sky130_fd_sc_hd__inv_2
XFILLER_48_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4982_ _4990_/CLK _4982_/D vssd1 vssd1 vccd1 vccd1 _4982_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_63_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3933_ _3933_/A _3933_/B _3933_/C _3933_/D vssd1 vssd1 vccd1 vccd1 _3933_/X sky130_fd_sc_hd__and4_1
X_3864_ _3873_/A _3864_/B vssd1 vssd1 vccd1 vccd1 _3864_/Y sky130_fd_sc_hd__nand2_1
X_2815_ _5314_/Q _4592_/A _2845_/A _2845_/B vssd1 vssd1 vccd1 vccd1 _2815_/Y sky130_fd_sc_hd__a22oi_2
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3795_ _5157_/Q _3783_/X _3791_/X _3794_/Y vssd1 vssd1 vccd1 vccd1 _5157_/D sky130_fd_sc_hd__o211a_1
X_2746_ _2908_/A vssd1 vssd1 vccd1 vccd1 _2746_/Y sky130_fd_sc_hd__inv_2
X_2677_ _5298_/Q vssd1 vssd1 vccd1 vccd1 _2729_/A sky130_fd_sc_hd__inv_2
X_4416_ _4416_/A _4416_/B vssd1 vssd1 vccd1 vccd1 _4416_/Y sky130_fd_sc_hd__nand2_1
XFILLER_59_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4347_ _4347_/A _4677_/B vssd1 vssd1 vccd1 vccd1 _4348_/B sky130_fd_sc_hd__nor2_1
X_4278_ _4525_/A _4527_/C _4525_/B vssd1 vssd1 vccd1 vccd1 _4513_/A sky130_fd_sc_hd__o21bai_1
X_3229_ _3177_/B _3037_/A _3232_/B _2888_/X vssd1 vssd1 vccd1 vccd1 _3229_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_27_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2600_ _2892_/A vssd1 vssd1 vccd1 vccd1 _2600_/X sky130_fd_sc_hd__clkbuf_2
X_3580_ _3586_/B _3586_/A vssd1 vssd1 vccd1 vccd1 _3582_/B sky130_fd_sc_hd__or2_1
X_2531_ _5046_/Q vssd1 vssd1 vccd1 vccd1 _4755_/A sky130_fd_sc_hd__inv_2
X_5250_ _5250_/CLK _5250_/D vssd1 vssd1 vccd1 vccd1 _5250_/Q sky130_fd_sc_hd__dfxtp_2
X_4201_ _4542_/A _4289_/A _4201_/C vssd1 vssd1 vccd1 vccd1 _4206_/A sky130_fd_sc_hd__or3_1
X_5181_ _5247_/CLK _5181_/D vssd1 vssd1 vccd1 vccd1 _5181_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4132_ _4132_/A vssd1 vssd1 vccd1 vccd1 _4183_/B sky130_fd_sc_hd__clkbuf_2
X_4063_ _4063_/A _4063_/B vssd1 vssd1 vccd1 vccd1 _4233_/A sky130_fd_sc_hd__nand2_2
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3014_ _5255_/Q vssd1 vssd1 vccd1 vccd1 _3789_/B sky130_fd_sc_hd__inv_2
XFILLER_36_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4965_ _5125_/Q _4965_/B vssd1 vssd1 vccd1 vccd1 _4966_/A sky130_fd_sc_hd__xor2_1
XPHY_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3916_ _3916_/A _4930_/A vssd1 vssd1 vccd1 vccd1 _3916_/Y sky130_fd_sc_hd__nand2_1
X_4896_ _4898_/A _4898_/B vssd1 vssd1 vccd1 vccd1 _4896_/Y sky130_fd_sc_hd__nor2_1
X_3847_ _3847_/A _3847_/B vssd1 vssd1 vccd1 vccd1 _3847_/Y sky130_fd_sc_hd__nand2_1
X_3778_ _3830_/A vssd1 vssd1 vccd1 vccd1 _3778_/X sky130_fd_sc_hd__clkbuf_2
X_2729_ _2729_/A _5031_/Q vssd1 vssd1 vccd1 vccd1 _2731_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_70_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_65_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4750_ _4767_/A _4767_/B vssd1 vssd1 vccd1 vccd1 _4750_/X sky130_fd_sc_hd__or2_1
X_3701_ _3705_/B _3701_/B vssd1 vssd1 vccd1 vccd1 _3701_/Y sky130_fd_sc_hd__nor2_1
X_4681_ _5036_/Q _5068_/Q vssd1 vssd1 vccd1 vccd1 _4801_/A sky130_fd_sc_hd__nor2_1
X_3632_ _3632_/A _3632_/B vssd1 vssd1 vccd1 vccd1 _3632_/Y sky130_fd_sc_hd__nor2_1
X_3563_ _3563_/A _3563_/B _3563_/C vssd1 vssd1 vccd1 vccd1 _3563_/Y sky130_fd_sc_hd__nand3_1
X_5302_ _5303_/CLK _5302_/D vssd1 vssd1 vccd1 vccd1 _5302_/Q sky130_fd_sc_hd__dfxtp_1
X_3494_ _3494_/A _3494_/B vssd1 vssd1 vccd1 vccd1 _3577_/A sky130_fd_sc_hd__nand2_1
X_2514_ _5049_/Q vssd1 vssd1 vccd1 vccd1 _4591_/A sky130_fd_sc_hd__inv_2
XFILLER_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5233_ _5268_/CLK _5233_/D vssd1 vssd1 vccd1 vccd1 _5233_/Q sky130_fd_sc_hd__dfxtp_2
X_5164_ _5288_/CLK _5164_/D vssd1 vssd1 vccd1 vccd1 _5164_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4115_ _4244_/A _4115_/B _4115_/C vssd1 vssd1 vccd1 vccd1 _4116_/C sky130_fd_sc_hd__nor3_2
XFILLER_68_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5095_ _5097_/CLK _5095_/D vssd1 vssd1 vccd1 vccd1 _5095_/Q sky130_fd_sc_hd__dfxtp_1
X_4046_ _4056_/B _4054_/A _4028_/A _4028_/B vssd1 vssd1 vccd1 vccd1 _4059_/B sky130_fd_sc_hd__o2bb2ai_4
XFILLER_17_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4948_ _4948_/A _4948_/B vssd1 vssd1 vccd1 vccd1 _4953_/A sky130_fd_sc_hd__nor2_1
XFILLER_12_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4879_ _5021_/Q _4475_/X _4876_/X _4878_/X _2837_/X vssd1 vssd1 vccd1 vccd1 _5021_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_59_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_74_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_65_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2994_ _5259_/Q vssd1 vssd1 vccd1 vccd1 _3779_/B sky130_fd_sc_hd__inv_2
X_4802_ _4806_/A _4806_/B _4686_/A vssd1 vssd1 vccd1 vccd1 _4803_/B sky130_fd_sc_hd__o21a_1
XFILLER_9_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4733_ _4733_/A _4733_/B _4733_/C vssd1 vssd1 vccd1 vccd1 _4734_/C sky130_fd_sc_hd__and3_1
X_4664_ _4664_/A vssd1 vssd1 vccd1 vccd1 _4827_/A sky130_fd_sc_hd__inv_2
X_3615_ _3615_/A vssd1 vssd1 vccd1 vccd1 _3615_/X sky130_fd_sc_hd__clkbuf_2
X_4595_ _4595_/A _4605_/A vssd1 vssd1 vccd1 vccd1 _4779_/B sky130_fd_sc_hd__or2_2
X_3546_ _3521_/Y _3524_/Y _3545_/Y vssd1 vssd1 vccd1 vccd1 _3546_/Y sky130_fd_sc_hd__a21oi_1
X_3477_ _3837_/B _5141_/Q vssd1 vssd1 vccd1 vccd1 _3620_/B sky130_fd_sc_hd__and2_1
X_5216_ _5221_/CLK _5216_/D vssd1 vssd1 vccd1 vccd1 _5216_/Q sky130_fd_sc_hd__dfxtp_1
X_5147_ _5221_/CLK _5147_/D vssd1 vssd1 vccd1 vccd1 _5147_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5078_ _5108_/CLK _5078_/D vssd1 vssd1 vccd1 vccd1 _5078_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4029_ _4029_/A _4029_/B vssd1 vssd1 vccd1 vccd1 _4036_/A sky130_fd_sc_hd__or2_2
XFILLER_71_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3400_ _3406_/B _3400_/B vssd1 vssd1 vccd1 vccd1 _3603_/B sky130_fd_sc_hd__nand2_2
X_4380_ _4382_/A _4710_/B vssd1 vssd1 vccd1 vccd1 _4381_/A sky130_fd_sc_hd__nor2_1
X_3331_ _3329_/X _3330_/Y _3306_/X vssd1 vssd1 vccd1 vccd1 _3331_/X sky130_fd_sc_hd__a21o_1
X_3262_ _3262_/A vssd1 vssd1 vccd1 vccd1 _3262_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_5001_ _5001_/CLK hold11/X vssd1 vssd1 vccd1 vccd1 _5002_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_85_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3193_ _3189_/Y _3191_/Y _3192_/Y vssd1 vssd1 vccd1 vccd1 _5253_/D sky130_fd_sc_hd__a21oi_1
XFILLER_38_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2977_ _3321_/A vssd1 vssd1 vccd1 vccd1 _2977_/X sky130_fd_sc_hd__buf_2
X_4716_ _4757_/B _4716_/B vssd1 vssd1 vccd1 vccd1 _4717_/B sky130_fd_sc_hd__nor2_2
X_4647_ _4849_/A _4849_/B _4646_/Y vssd1 vssd1 vccd1 vccd1 _4840_/B sky130_fd_sc_hd__a21oi_1
X_4578_ _4578_/A _4578_/B vssd1 vssd1 vccd1 vccd1 _4578_/X sky130_fd_sc_hd__and2_1
X_3529_ _3794_/B _5157_/Q vssd1 vssd1 vccd1 vccd1 _3531_/C sky130_fd_sc_hd__and2_1
XFILLER_39_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2900_ _5275_/Q _2841_/X _2896_/Y _2898_/X _2899_/X vssd1 vssd1 vccd1 vccd1 _5275_/D
+ sky130_fd_sc_hd__o221a_1
X_3880_ _5125_/Q vssd1 vssd1 vccd1 vccd1 _3933_/B sky130_fd_sc_hd__inv_2
XFILLER_31_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2831_ _4589_/A vssd1 vssd1 vccd1 vccd1 _4169_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2762_ _5307_/Q _4601_/A vssd1 vssd1 vccd1 vccd1 _2762_/Y sky130_fd_sc_hd__nor2_1
XFILLER_8_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4501_ _4453_/X _5067_/Q _4473_/X _4500_/X vssd1 vssd1 vccd1 vccd1 _5067_/D sky130_fd_sc_hd__o211a_1
XANTENNA_0 enable_in vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2693_ _3000_/B _3000_/A _3010_/A _3002_/B vssd1 vssd1 vccd1 vccd1 _2997_/A sky130_fd_sc_hd__o22ai_4
X_4432_ _4785_/A vssd1 vssd1 vccd1 vccd1 _4432_/X sky130_fd_sc_hd__clkbuf_2
X_4363_ _4347_/A _4677_/B _4361_/Y _4359_/A _4362_/X vssd1 vssd1 vccd1 vccd1 _4474_/B
+ sky130_fd_sc_hd__o221a_2
X_4294_ _5084_/Q _4634_/B _5083_/Q _5051_/Q vssd1 vssd1 vccd1 vccd1 _4575_/B sky130_fd_sc_hd__o211a_1
X_3314_ _3313_/B _3313_/A _3292_/X vssd1 vssd1 vccd1 vccd1 _3314_/X sky130_fd_sc_hd__a21o_1
X_3245_ _3242_/X _2506_/X _3243_/Y _3244_/Y vssd1 vssd1 vccd1 vccd1 _5245_/D sky130_fd_sc_hd__a31oi_1
X_3176_ _3176_/A vssd1 vssd1 vccd1 vccd1 _3177_/B sky130_fd_sc_hd__inv_2
XFILLER_81_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_81_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_77_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_66_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3030_ _5187_/Q _3713_/B vssd1 vssd1 vccd1 vccd1 _3204_/A sky130_fd_sc_hd__nor2_4
XFILLER_36_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4981_ _4990_/CLK hold42/X vssd1 vssd1 vccd1 vccd1 _4982_/D sky130_fd_sc_hd__dfxtp_1
XFILLER_63_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3932_ _5118_/Q _3931_/Y _4930_/A _5007_/Q vssd1 vssd1 vccd1 vccd1 _3933_/D sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_43_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5199_/CLK sky130_fd_sc_hd__clkbuf_16
X_3863_ _3863_/A vssd1 vssd1 vccd1 vccd1 _3873_/A sky130_fd_sc_hd__clkbuf_2
X_2814_ _2814_/A vssd1 vssd1 vccd1 vccd1 _2845_/B sky130_fd_sc_hd__inv_2
X_3794_ _3794_/A _3794_/B vssd1 vssd1 vccd1 vccd1 _3794_/Y sky130_fd_sc_hd__nand2_1
X_2745_ _2737_/B _2739_/A _5033_/Q _2735_/Y vssd1 vssd1 vccd1 vccd1 _2908_/A sky130_fd_sc_hd__a31o_1
X_2676_ _4666_/A _5299_/Q vssd1 vssd1 vccd1 vccd1 _2728_/B sky130_fd_sc_hd__nand2_1
X_4415_ _4778_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _4415_/Y sky130_fd_sc_hd__nor2_1
X_4346_ _5070_/Q vssd1 vssd1 vccd1 vccd1 _4677_/B sky130_fd_sc_hd__inv_2
XFILLER_86_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4277_ _4277_/A _4617_/B vssd1 vssd1 vccd1 vccd1 _4525_/B sky130_fd_sc_hd__nor2_1
X_3228_ _3037_/A _3232_/B _3177_/B vssd1 vssd1 vccd1 vccd1 _3228_/X sky130_fd_sc_hd__o21a_1
XFILLER_54_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3159_ _5180_/Q _3732_/B vssd1 vssd1 vccd1 vccd1 _3167_/A sky130_fd_sc_hd__nor2_1
XFILLER_54_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_34_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5251_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_50_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_25_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 _5274_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_41_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2530_ _2605_/A vssd1 vssd1 vccd1 vccd1 _2546_/A sky130_fd_sc_hd__buf_1
X_4200_ _5087_/Q vssd1 vssd1 vccd1 vccd1 _4289_/A sky130_fd_sc_hd__inv_2
XFILLER_5_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5180_ _5247_/CLK _5180_/D vssd1 vssd1 vccd1 vccd1 _5180_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4131_ _4149_/A _4131_/B vssd1 vssd1 vccd1 vccd1 _4139_/A sky130_fd_sc_hd__nand2_1
X_4062_ _4057_/A _4057_/B _4059_/B vssd1 vssd1 vccd1 vccd1 _4062_/X sky130_fd_sc_hd__o21a_1
X_3013_ _5256_/Q _2977_/X _3009_/X _3012_/Y _2971_/X vssd1 vssd1 vccd1 vccd1 _5256_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_36_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_16_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5085_/CLK sky130_fd_sc_hd__clkbuf_16
X_4964_ _4964_/A _4966_/B vssd1 vssd1 vccd1 vccd1 _4964_/X sky130_fd_sc_hd__and2_1
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3915_ _5117_/Q vssd1 vssd1 vccd1 vccd1 _4930_/A sky130_fd_sc_hd__inv_2
XFILLER_51_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4895_ _4890_/Y _4891_/X _4899_/B vssd1 vssd1 vccd1 vccd1 _5018_/D sky130_fd_sc_hd__o21a_1
XFILLER_32_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3846_ _5138_/Q _3835_/X _3844_/X _3845_/Y vssd1 vssd1 vccd1 vccd1 _5138_/D sky130_fd_sc_hd__o211a_1
X_3777_ _3843_/A vssd1 vssd1 vccd1 vccd1 _3830_/A sky130_fd_sc_hd__clkbuf_2
X_2728_ _2678_/Y _2728_/B vssd1 vssd1 vccd1 vccd1 _2946_/A sky130_fd_sc_hd__and2b_1
X_2659_ _2772_/A _2657_/Y _2772_/B vssd1 vssd1 vccd1 vccd1 _2865_/B sky130_fd_sc_hd__o21ba_1
XFILLER_59_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4329_ _5096_/Q _5064_/Q vssd1 vssd1 vccd1 vccd1 _4332_/A sky130_fd_sc_hd__nor2_1
XFILLER_59_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_70_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_88_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_77_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3700_ _3700_/A _3700_/B vssd1 vssd1 vccd1 vccd1 _3701_/B sky130_fd_sc_hd__nand2_1
X_4680_ _4794_/A _4797_/A vssd1 vssd1 vccd1 vccd1 _4688_/A sky130_fd_sc_hd__nand2_1
X_3631_ _3845_/B _5138_/Q _3630_/X vssd1 vssd1 vccd1 vccd1 _3632_/B sky130_fd_sc_hd__o21a_1
X_3562_ _3562_/A _3562_/B vssd1 vssd1 vccd1 vccd1 _3563_/C sky130_fd_sc_hd__nand2_1
X_2513_ _3863_/A vssd1 vssd1 vccd1 vccd1 _2524_/A sky130_fd_sc_hd__clkbuf_2
X_5301_ _5301_/CLK _5301_/D vssd1 vssd1 vccd1 vccd1 _5301_/Q sky130_fd_sc_hd__dfxtp_1
X_3493_ _3824_/B _5146_/Q vssd1 vssd1 vccd1 vccd1 _3494_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5232_ _5236_/CLK _5232_/D vssd1 vssd1 vccd1 vccd1 _5232_/Q sky130_fd_sc_hd__dfxtp_1
Xclkbuf_leaf_5_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5303_/CLK sky130_fd_sc_hd__clkbuf_16
X_5163_ _5274_/CLK _5163_/D vssd1 vssd1 vccd1 vccd1 _5163_/Q sky130_fd_sc_hd__dfxtp_1
X_4114_ _4156_/C vssd1 vssd1 vccd1 vccd1 _4115_/C sky130_fd_sc_hd__clkbuf_2
X_5094_ _5096_/CLK _5094_/D vssd1 vssd1 vccd1 vccd1 _5094_/Q sky130_fd_sc_hd__dfxtp_1
X_4045_ _4056_/B _4045_/B _4045_/C vssd1 vssd1 vccd1 vccd1 _4051_/B sky130_fd_sc_hd__nand3_4
XFILLER_52_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_4947_ _4951_/A _4947_/B vssd1 vssd1 vccd1 vccd1 _4947_/X sky130_fd_sc_hd__and2_1
XFILLER_33_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4878_ _4878_/A _4878_/B _4878_/C vssd1 vssd1 vccd1 vccd1 _4878_/X sky130_fd_sc_hd__and3_1
X_3829_ _5144_/Q _3822_/X _3817_/X _3828_/Y vssd1 vssd1 vccd1 vccd1 _5144_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4801_ _4801_/A _4801_/B vssd1 vssd1 vccd1 vccd1 _4803_/A sky130_fd_sc_hd__nor2_1
X_2993_ _2993_/A _2993_/B _2993_/C vssd1 vssd1 vccd1 vccd1 _2993_/X sky130_fd_sc_hd__and3_1
XFILLER_21_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4732_ _4733_/A _4733_/B _4733_/C vssd1 vssd1 vccd1 vccd1 _4734_/B sky130_fd_sc_hd__a21oi_1
XFILLER_21_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4663_ _4663_/A _4823_/B vssd1 vssd1 vccd1 vccd1 _4664_/A sky130_fd_sc_hd__nand2_1
X_3614_ _3614_/A _3614_/B vssd1 vssd1 vccd1 vccd1 _3614_/Y sky130_fd_sc_hd__nand2_1
X_4594_ _4778_/B _4594_/B vssd1 vssd1 vccd1 vccd1 _4605_/A sky130_fd_sc_hd__nor2_1
X_3545_ _3545_/A vssd1 vssd1 vccd1 vccd1 _3545_/Y sky130_fd_sc_hd__inv_2
X_3476_ _5141_/Q _3837_/B vssd1 vssd1 vccd1 vccd1 _3620_/A sky130_fd_sc_hd__nor2_1
X_5215_ _5221_/CLK _5215_/D vssd1 vssd1 vccd1 vccd1 _5215_/Q sky130_fd_sc_hd__dfxtp_1
X_5146_ _5251_/CLK _5146_/D vssd1 vssd1 vccd1 vccd1 _5146_/Q sky130_fd_sc_hd__dfxtp_1
X_5077_ _5108_/CLK _5077_/D vssd1 vssd1 vccd1 vccd1 _5077_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4028_ _4028_/A _4028_/B vssd1 vssd1 vccd1 vccd1 _4043_/A sky130_fd_sc_hd__nor2_2
XFILLER_71_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_79_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3330_ _3330_/A _3330_/B vssd1 vssd1 vccd1 vccd1 _3330_/Y sky130_fd_sc_hd__nand2_1
X_5000_ _5001_/CLK _5000_/D vssd1 vssd1 vccd1 vccd1 _5000_/Q sky130_fd_sc_hd__dfxtp_1
X_3261_ _3267_/A _3056_/A _3064_/B _3206_/X vssd1 vssd1 vccd1 vccd1 _3261_/X sky130_fd_sc_hd__a31o_1
X_3192_ _5253_/Q _3199_/C _4238_/B vssd1 vssd1 vccd1 vccd1 _3192_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_78_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_81_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2976_ _2901_/X _2973_/X _2961_/X _2975_/Y vssd1 vssd1 vccd1 vccd1 _5262_/D sky130_fd_sc_hd__o211a_1
X_4715_ _4715_/A vssd1 vssd1 vccd1 vccd1 _4716_/B sky130_fd_sc_hd__inv_2
X_4646_ _4848_/A _4852_/B vssd1 vssd1 vccd1 vccd1 _4646_/Y sky130_fd_sc_hd__nand2_1
X_4577_ _4578_/B _4578_/A _4912_/B vssd1 vssd1 vccd1 vccd1 _4577_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_30_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3528_ _5157_/Q _3794_/B vssd1 vssd1 vccd1 vccd1 _3531_/B sky130_fd_sc_hd__nor2_1
X_3459_ _5136_/Q _3851_/B vssd1 vssd1 vccd1 vccd1 _3640_/B sky130_fd_sc_hd__or2_1
XFILLER_57_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_69_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5129_ _5197_/CLK _5129_/D vssd1 vssd1 vccd1 vccd1 _5129_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2830_ hold44/X vssd1 vssd1 vccd1 vccd1 _4589_/A sky130_fd_sc_hd__clkbuf_2
XPHY_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2761_ _2885_/B _2885_/A _2893_/B vssd1 vssd1 vccd1 vccd1 _2769_/B sky130_fd_sc_hd__or3_1
X_4500_ _4496_/A _4499_/Y _4204_/X vssd1 vssd1 vccd1 vccd1 _4500_/X sky130_fd_sc_hd__a21o_1
X_2692_ _5288_/Q _4633_/A _3008_/A _3018_/B vssd1 vssd1 vccd1 vccd1 _3002_/B sky130_fd_sc_hd__a22oi_4
XANTENNA_1 oversample_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4431_ _4427_/Y _4429_/X _4428_/Y _4742_/B vssd1 vssd1 vccd1 vccd1 _4431_/Y sky130_fd_sc_hd__o31ai_1
XFILLER_6_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4362_ _4482_/B _4362_/B vssd1 vssd1 vccd1 vccd1 _4362_/X sky130_fd_sc_hd__or2_1
X_4293_ _5052_/Q vssd1 vssd1 vccd1 vccd1 _4634_/B sky130_fd_sc_hd__clkbuf_2
X_3313_ _3313_/A _3313_/B vssd1 vssd1 vccd1 vccd1 _3313_/Y sky130_fd_sc_hd__nor2_1
X_3244_ _5245_/Q _3563_/B _2889_/X vssd1 vssd1 vccd1 vccd1 _3244_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_39_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3175_ _3175_/A _3175_/B vssd1 vssd1 vccd1 vccd1 _3176_/A sky130_fd_sc_hd__nor2_1
XFILLER_39_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2959_ _5265_/Q _2924_/X _2956_/X _2958_/Y _2899_/X vssd1 vssd1 vccd1 vccd1 _5265_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_22_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4629_ _5023_/Q _5055_/Q vssd1 vssd1 vccd1 vccd1 _4862_/C sky130_fd_sc_hd__nand2_1
XFILLER_89_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_89_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_85_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4980_ _4913_/B _5004_/Q _4980_/S vssd1 vssd1 vccd1 vccd1 _4980_/X sky130_fd_sc_hd__mux2_1
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3931_ _5008_/Q vssd1 vssd1 vccd1 vccd1 _3931_/Y sky130_fd_sc_hd__inv_2
XFILLER_51_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3862_ _3862_/A vssd1 vssd1 vccd1 vccd1 _3862_/X sky130_fd_sc_hd__clkbuf_2
X_2813_ _2796_/Y _2812_/Y _2776_/Y vssd1 vssd1 vccd1 vccd1 _2845_/A sky130_fd_sc_hd__o21bai_2
XFILLER_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3793_ _5158_/Q _3783_/X _3791_/X _3792_/Y vssd1 vssd1 vccd1 vccd1 _5158_/D sky130_fd_sc_hd__o211a_1
XFILLER_8_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2744_ _2808_/A _2734_/Y _2743_/Y vssd1 vssd1 vccd1 vccd1 _2744_/Y sky130_fd_sc_hd__o21bai_1
X_2675_ _2675_/A _2675_/B _2674_/Y vssd1 vssd1 vccd1 vccd1 _2811_/A sky130_fd_sc_hd__or3b_4
X_4414_ _4412_/Y _4733_/B _4214_/X vssd1 vssd1 vccd1 vccd1 _5082_/D sky130_fd_sc_hd__a21oi_1
X_4345_ _5102_/Q _5070_/Q vssd1 vssd1 vccd1 vccd1 _4362_/B sky130_fd_sc_hd__nor2_1
X_4276_ _5062_/Q vssd1 vssd1 vccd1 vccd1 _4617_/B sky130_fd_sc_hd__inv_2
XFILLER_67_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3227_ _3231_/B _3227_/B vssd1 vssd1 vccd1 vccd1 _3232_/B sky130_fd_sc_hd__nor2_2
X_3158_ _5276_/Q vssd1 vssd1 vccd1 vccd1 _3732_/B sky130_fd_sc_hd__inv_2
XFILLER_36_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3089_ _5161_/Q _3785_/B vssd1 vssd1 vccd1 vccd1 _3090_/A sky130_fd_sc_hd__nor2_1
XFILLER_42_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_77_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_68_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4130_ _4133_/A _4375_/A _4129_/Y vssd1 vssd1 vccd1 vccd1 _5108_/D sky130_fd_sc_hd__a21oi_1
XFILLER_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4061_ _4057_/Y _4052_/A _4580_/A _4060_/Y vssd1 vssd1 vccd1 vccd1 _4226_/B sky130_fd_sc_hd__o211ai_4
XFILLER_68_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3012_ _3012_/A _3705_/A vssd1 vssd1 vccd1 vccd1 _3012_/Y sky130_fd_sc_hd__nand2_1
X_4963_ _4963_/A _4965_/B vssd1 vssd1 vccd1 vccd1 _4964_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3914_ _3907_/X _4977_/X _3911_/X _3913_/Y vssd1 vssd1 vccd1 vccd1 _5118_/D sky130_fd_sc_hd__o211a_1
XFILLER_32_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4894_ _4898_/A _4980_/S _4132_/A vssd1 vssd1 vccd1 vccd1 _4899_/B sky130_fd_sc_hd__o21a_1
XFILLER_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3845_ _3847_/A _3845_/B vssd1 vssd1 vccd1 vccd1 _3845_/Y sky130_fd_sc_hd__nand2_1
X_3776_ _5164_/Q _3768_/X _3762_/X _3775_/Y vssd1 vssd1 vccd1 vccd1 _5164_/D sky130_fd_sc_hd__o211a_1
X_2727_ _2723_/B _2957_/B _2726_/Y vssd1 vssd1 vccd1 vccd1 _2943_/B sky130_fd_sc_hd__o21a_1
X_2658_ _4704_/A _5311_/Q vssd1 vssd1 vccd1 vccd1 _2772_/B sky130_fd_sc_hd__and2_1
X_2589_ _2602_/A _4661_/A vssd1 vssd1 vccd1 vccd1 _2589_/Y sky130_fd_sc_hd__nand2_1
XFILLER_86_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4328_ _4328_/A _4328_/B vssd1 vssd1 vccd1 vccd1 _4520_/B sky130_fd_sc_hd__nand2_1
XFILLER_86_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_74_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4259_ _4364_/B vssd1 vssd1 vccd1 vccd1 _4259_/Y sky130_fd_sc_hd__inv_2
XFILLER_86_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_86_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_67_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_88_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_88_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3630_ _3635_/B _3635_/A vssd1 vssd1 vccd1 vccd1 _3630_/X sky130_fd_sc_hd__or2_1
X_3561_ _3558_/X _3559_/Y _3560_/Y vssd1 vssd1 vccd1 vccd1 _5217_/D sky130_fd_sc_hd__a21oi_1
X_2512_ _3769_/A vssd1 vssd1 vccd1 vccd1 _3863_/A sky130_fd_sc_hd__clkbuf_2
X_5300_ _5303_/CLK _5300_/D vssd1 vssd1 vccd1 vccd1 _5300_/Q sky130_fd_sc_hd__dfxtp_1
X_3492_ _5146_/Q _3824_/B vssd1 vssd1 vccd1 vccd1 _3494_/A sky130_fd_sc_hd__or2_2
X_5231_ _5268_/CLK _5231_/D vssd1 vssd1 vccd1 vccd1 _5231_/Q sky130_fd_sc_hd__dfxtp_2
X_5162_ _5274_/CLK _5162_/D vssd1 vssd1 vccd1 vccd1 _5162_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5093_ _5096_/CLK _5093_/D vssd1 vssd1 vccd1 vccd1 _5093_/Q sky130_fd_sc_hd__dfxtp_1
X_4113_ _4111_/X _4112_/X _4094_/X _4095_/X _5111_/Q vssd1 vssd1 vccd1 vccd1 _4116_/B
+ sky130_fd_sc_hd__a41oi_1
XFILLER_29_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4044_ _4234_/B _4059_/A vssd1 vssd1 vccd1 vccd1 _4047_/A sky130_fd_sc_hd__nand2_1
XFILLER_64_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4946_ _4946_/A _4949_/B vssd1 vssd1 vccd1 vccd1 _4947_/B sky130_fd_sc_hd__nor2_1
X_4877_ _4881_/A _4877_/B vssd1 vssd1 vccd1 vccd1 _4878_/A sky130_fd_sc_hd__nand2_1
X_3828_ _3833_/A _3828_/B vssd1 vssd1 vccd1 vccd1 _3828_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3759_ _5170_/Q _3754_/X _3749_/X _3758_/Y vssd1 vssd1 vccd1 vccd1 _5170_/D sky130_fd_sc_hd__o211a_1
XFILLER_59_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4800_ _4798_/X _4799_/Y _4116_/A vssd1 vssd1 vccd1 vccd1 _5037_/D sky130_fd_sc_hd__a21oi_1
X_2992_ _2993_/A _2993_/B _2993_/C vssd1 vssd1 vccd1 vccd1 _2992_/Y sky130_fd_sc_hd__a21oi_2
XFILLER_61_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4731_ _5050_/Q _5082_/Q vssd1 vssd1 vccd1 vccd1 _4733_/C sky130_fd_sc_hd__xnor2_1
X_4662_ _5031_/Q _5063_/Q vssd1 vssd1 vccd1 vccd1 _4823_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3613_ _3613_/A vssd1 vssd1 vccd1 vccd1 _3613_/X sky130_fd_sc_hd__clkbuf_2
X_4593_ _5041_/Q _5073_/Q vssd1 vssd1 vccd1 vccd1 _4595_/A sky130_fd_sc_hd__nor2_1
X_3544_ _3544_/A _3544_/B vssd1 vssd1 vccd1 vccd1 _3545_/A sky130_fd_sc_hd__or2_1
X_3475_ _5237_/Q vssd1 vssd1 vccd1 vccd1 _3837_/B sky130_fd_sc_hd__inv_2
X_5214_ _5221_/CLK _5214_/D vssd1 vssd1 vccd1 vccd1 _5214_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_5145_ _5251_/CLK _5145_/D vssd1 vssd1 vccd1 vccd1 _5145_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_28_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5076_ _5076_/CLK _5076_/D vssd1 vssd1 vccd1 vccd1 _5076_/Q sky130_fd_sc_hd__dfxtp_1
X_4027_ _4022_/A _4022_/B _4022_/C _4048_/B vssd1 vssd1 vccd1 vccd1 _4028_/B sky130_fd_sc_hd__a31oi_4
XFILLER_25_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4929_ _5117_/Q _5116_/Q vssd1 vssd1 vccd1 vccd1 _4931_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_90_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3260_ _3267_/A _3064_/B _3056_/A vssd1 vssd1 vccd1 vccd1 _3260_/Y sky130_fd_sc_hd__a21oi_1
X_3191_ _3199_/B _3190_/Y _3605_/A vssd1 vssd1 vccd1 vccd1 _3191_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_78_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_81_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4714_ _4720_/A _4714_/B vssd1 vssd1 vccd1 vccd1 _4715_/A sky130_fd_sc_hd__nor2_1
X_2975_ _3276_/A _3771_/B vssd1 vssd1 vccd1 vccd1 _2975_/Y sky130_fd_sc_hd__nand2_1
X_4645_ _4645_/A _4645_/B vssd1 vssd1 vccd1 vccd1 _4852_/B sky130_fd_sc_hd__nor2_1
X_4576_ _4576_/A _4576_/B vssd1 vssd1 vccd1 vccd1 _4578_/A sky130_fd_sc_hd__and2_1
X_3527_ _5253_/Q vssd1 vssd1 vccd1 vccd1 _3794_/B sky130_fd_sc_hd__inv_2
XFILLER_89_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3458_ _5232_/Q vssd1 vssd1 vccd1 vccd1 _3851_/B sky130_fd_sc_hd__inv_2
XFILLER_57_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3389_ _3805_/B _5153_/Q vssd1 vssd1 vccd1 vccd1 _3391_/A sky130_fd_sc_hd__and2_1
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5128_ _5195_/CLK _5128_/D vssd1 vssd1 vccd1 vccd1 _5128_/Q sky130_fd_sc_hd__dfxtp_2
XFILLER_55_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5059_ _5062_/CLK _5059_/D vssd1 vssd1 vccd1 vccd1 _5059_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_55_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2760_ _2760_/A _2760_/B vssd1 vssd1 vccd1 vccd1 _2893_/B sky130_fd_sc_hd__nand2_1
XFILLER_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2691_ _3017_/B _4631_/A vssd1 vssd1 vccd1 vccd1 _3018_/B sky130_fd_sc_hd__nand2_2
XANTENNA_2 oversample_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4430_ _4427_/Y _4428_/Y _4429_/X vssd1 vssd1 vccd1 vccd1 _4430_/X sky130_fd_sc_hd__o21a_1
XFILLER_6_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4361_ _4494_/B _4355_/A _4494_/A vssd1 vssd1 vccd1 vccd1 _4361_/Y sky130_fd_sc_hd__o21bai_1
X_4292_ _5084_/Q _5052_/Q vssd1 vssd1 vccd1 vccd1 _4581_/B sky130_fd_sc_hd__and2_1
XFILLER_3_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3312_ _3771_/B _5166_/Q _3311_/X vssd1 vssd1 vccd1 vccd1 _3313_/B sky130_fd_sc_hd__o21a_1
X_3243_ _3243_/A _3243_/B _3243_/C vssd1 vssd1 vccd1 vccd1 _3243_/Y sky130_fd_sc_hd__nand3_1
XFILLER_66_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3174_ _3174_/A _3174_/B vssd1 vssd1 vccd1 vccd1 _3231_/B sky130_fd_sc_hd__nand2_1
XFILLER_54_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2958_ _2958_/A _2958_/B vssd1 vssd1 vccd1 vccd1 _2958_/Y sky130_fd_sc_hd__nor2_1
X_4628_ _4628_/A _4628_/B vssd1 vssd1 vccd1 vccd1 _4630_/A sky130_fd_sc_hd__nand2_1
X_2889_ _4132_/A vssd1 vssd1 vccd1 vccd1 _2889_/X sky130_fd_sc_hd__clkbuf_4
X_4559_ _4559_/A _4571_/C _4559_/C vssd1 vssd1 vccd1 vccd1 _4559_/X sky130_fd_sc_hd__and3_1
XFILLER_1_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_89_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_66_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput50 _5194_/Q vssd1 vssd1 vccd1 vccd1 data_out[4] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3930_ _4962_/A _5014_/Q vssd1 vssd1 vccd1 vccd1 _3933_/C sky130_fd_sc_hd__nand2_1
XFILLER_63_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3861_ _5132_/Q _3849_/X _3857_/X _3860_/Y vssd1 vssd1 vccd1 vccd1 _5132_/D sky130_fd_sc_hd__o211a_1
XFILLER_82_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3792_ _3794_/A _3792_/B vssd1 vssd1 vccd1 vccd1 _3792_/Y sky130_fd_sc_hd__nand2_1
X_2812_ _2902_/A _2902_/B _2765_/X vssd1 vssd1 vccd1 vccd1 _2812_/Y sky130_fd_sc_hd__a21oi_2
X_2743_ _2937_/A _2940_/A vssd1 vssd1 vccd1 vccd1 _2743_/Y sky130_fd_sc_hd__nand2_1
X_2674_ _2674_/A _2910_/A vssd1 vssd1 vccd1 vccd1 _2674_/Y sky130_fd_sc_hd__nand2_1
X_4413_ _4542_/A _5082_/Q vssd1 vssd1 vccd1 vccd1 _4733_/B sky130_fd_sc_hd__nand2_1
X_4344_ _4344_/A _4482_/B vssd1 vssd1 vccd1 vccd1 _4487_/A sky130_fd_sc_hd__and2_1
XFILLER_86_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4275_ _5093_/Q _5061_/Q vssd1 vssd1 vccd1 vccd1 _4527_/C sky130_fd_sc_hd__nand2_1
X_3226_ _3224_/Y _3225_/Y _3202_/X vssd1 vssd1 vccd1 vccd1 _5248_/D sky130_fd_sc_hd__a21oi_1
XFILLER_82_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3157_ _5181_/Q _3730_/B vssd1 vssd1 vccd1 vccd1 _3241_/A sky130_fd_sc_hd__nor2_1
XFILLER_36_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3088_ _5257_/Q vssd1 vssd1 vccd1 vccd1 _3785_/B sky130_fd_sc_hd__inv_2
XFILLER_42_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_68_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4060_ _4060_/A _4234_/B vssd1 vssd1 vccd1 vccd1 _4060_/Y sky130_fd_sc_hd__nand2_2
XFILLER_64_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3011_ _3011_/A vssd1 vssd1 vccd1 vccd1 _3705_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4962_ _4962_/A _4962_/B vssd1 vssd1 vccd1 vccd1 _4965_/B sky130_fd_sc_hd__nor2_1
XFILLER_17_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3913_ _3916_/A _3913_/B vssd1 vssd1 vccd1 vccd1 _3913_/Y sky130_fd_sc_hd__nand2_1
X_4893_ _4893_/A _4912_/A vssd1 vssd1 vccd1 vccd1 _4980_/S sky130_fd_sc_hd__nor2_1
X_3844_ _3911_/A vssd1 vssd1 vccd1 vccd1 _3844_/X sky130_fd_sc_hd__clkbuf_2
X_3775_ _3781_/A _3775_/B vssd1 vssd1 vccd1 vccd1 _3775_/Y sky130_fd_sc_hd__nand2_1
X_2726_ _2726_/A vssd1 vssd1 vccd1 vccd1 _2726_/Y sky130_fd_sc_hd__inv_2
X_2657_ _5310_/Q _4701_/A vssd1 vssd1 vccd1 vccd1 _2657_/Y sky130_fd_sc_hd__nor2_1
X_2588_ _5031_/Q vssd1 vssd1 vccd1 vccd1 _4661_/A sky130_fd_sc_hd__inv_2
XFILLER_59_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4327_ _5095_/Q _5063_/Q vssd1 vssd1 vccd1 vccd1 _4328_/B sky130_fd_sc_hd__nand2_1
X_4258_ _4258_/A _4601_/B vssd1 vssd1 vccd1 vccd1 _4364_/B sky130_fd_sc_hd__nor2_2
XFILLER_86_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3209_ _5251_/Q _2977_/X _3205_/Y _3207_/X _3208_/X vssd1 vssd1 vccd1 vccd1 _5251_/D
+ sky130_fd_sc_hd__o221a_1
X_4189_ _5092_/Q _4185_/A _4188_/Y vssd1 vssd1 vccd1 vccd1 _5092_/D sky130_fd_sc_hd__o21a_1
XFILLER_82_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_88_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_77_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_77_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3560_ _5217_/Q _3199_/C _3533_/X vssd1 vssd1 vccd1 vccd1 _3560_/Y sky130_fd_sc_hd__o21ai_1
X_2511_ _2888_/A vssd1 vssd1 vccd1 vccd1 _3769_/A sky130_fd_sc_hd__buf_2
X_3491_ _5242_/Q vssd1 vssd1 vccd1 vccd1 _3824_/B sky130_fd_sc_hd__inv_2
XFILLER_5_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5230_ _5251_/CLK _5230_/D vssd1 vssd1 vccd1 vccd1 _5230_/Q sky130_fd_sc_hd__dfxtp_2
X_5161_ _5274_/CLK _5161_/D vssd1 vssd1 vccd1 vccd1 _5161_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_68_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5092_ _5097_/CLK _5092_/D vssd1 vssd1 vccd1 vccd1 _5092_/Q sky130_fd_sc_hd__dfxtp_1
X_4112_ _4180_/B vssd1 vssd1 vccd1 vccd1 _4112_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_83_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4043_ _4043_/A _4056_/B _4054_/A vssd1 vssd1 vccd1 vccd1 _4059_/A sky130_fd_sc_hd__nand3_4
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4945_ _4948_/B vssd1 vssd1 vccd1 vccd1 _4949_/B sky130_fd_sc_hd__inv_2
X_4876_ _4874_/Y _4881_/A _4877_/B _3879_/A vssd1 vssd1 vccd1 vccd1 _4876_/X sky130_fd_sc_hd__a31o_1
X_3827_ _5145_/Q _3822_/X _3817_/X _3826_/Y vssd1 vssd1 vccd1 vccd1 _5145_/D sky130_fd_sc_hd__o211a_1
XFILLER_20_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3758_ _3765_/A _3758_/B vssd1 vssd1 vccd1 vccd1 _3758_/Y sky130_fd_sc_hd__nand2_1
X_2709_ _2709_/A vssd1 vssd1 vccd1 vccd1 _2802_/A sky130_fd_sc_hd__inv_2
X_3689_ _5193_/Q _3650_/X _3687_/Y _3688_/X _3644_/X vssd1 vssd1 vccd1 vccd1 _5193_/D
+ sky130_fd_sc_hd__o221a_1
XFILLER_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_74_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_82_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_78_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_65_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2991_ _2991_/A _2991_/B vssd1 vssd1 vccd1 vccd1 _2993_/C sky130_fd_sc_hd__nor2_1
XFILLER_61_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_4730_ _4728_/B _4736_/B _4417_/A vssd1 vssd1 vccd1 vccd1 _4733_/A sky130_fd_sc_hd__o21ai_1
XFILLER_14_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4661_ _4661_/A _4661_/B vssd1 vssd1 vccd1 vccd1 _4663_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3612_ _5207_/Q _3596_/X _3609_/X _3611_/Y _3591_/X vssd1 vssd1 vccd1 vccd1 _5207_/D
+ sky130_fd_sc_hd__o221a_1
X_4592_ _4592_/A _4592_/B vssd1 vssd1 vccd1 vccd1 _4744_/B sky130_fd_sc_hd__nor2_2
X_3543_ _3541_/Y _3542_/Y _3202_/X vssd1 vssd1 vccd1 vccd1 _5220_/D sky130_fd_sc_hd__a21oi_1
X_3474_ _3629_/A _3629_/B _3473_/X vssd1 vssd1 vccd1 vccd1 _3618_/B sky130_fd_sc_hd__a21oi_2
X_5213_ _5251_/CLK _5213_/D vssd1 vssd1 vccd1 vccd1 _5213_/Q sky130_fd_sc_hd__dfxtp_1
X_5144_ _5251_/CLK _5144_/D vssd1 vssd1 vccd1 vccd1 _5144_/Q sky130_fd_sc_hd__dfxtp_1
X_5075_ _5109_/CLK _5075_/D vssd1 vssd1 vccd1 vccd1 _5075_/Q sky130_fd_sc_hd__dfxtp_1
X_4026_ _4063_/A _4064_/A _4063_/B vssd1 vssd1 vccd1 vccd1 _4234_/B sky130_fd_sc_hd__nand3_4
XFILLER_37_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4928_ _5116_/Q _4932_/A vssd1 vssd1 vccd1 vccd1 _4928_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4859_ _4859_/A _4871_/C vssd1 vssd1 vccd1 vccd1 _4865_/B sky130_fd_sc_hd__and2_1
XFILLER_60_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_79_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_69_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_75_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_90_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3190_ _3190_/A _3190_/B _3190_/C vssd1 vssd1 vccd1 vccd1 _3190_/Y sky130_fd_sc_hd__nor3_1
XFILLER_38_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2974_ _5262_/Q vssd1 vssd1 vccd1 vccd1 _3771_/B sky130_fd_sc_hd__inv_2
X_4713_ _4755_/A _4713_/B vssd1 vssd1 vccd1 vccd1 _4714_/B sky130_fd_sc_hd__nor2_2
X_4644_ _4644_/A _4852_/C vssd1 vssd1 vccd1 vccd1 _4848_/A sky130_fd_sc_hd__and2_1
X_4575_ _4581_/B _4575_/B vssd1 vssd1 vccd1 vccd1 _4578_/B sky130_fd_sc_hd__nor2_1
X_3526_ _3539_/B _3539_/A _3544_/A _3525_/Y vssd1 vssd1 vccd1 vccd1 _3541_/B sky130_fd_sc_hd__o22ai_4
XFILLER_89_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3457_ _3652_/A _3652_/B _3456_/X vssd1 vssd1 vccd1 vccd1 _3638_/B sky130_fd_sc_hd__a21oi_1
X_3388_ _5153_/Q _3805_/B vssd1 vssd1 vccd1 vccd1 _3390_/A sky130_fd_sc_hd__nor2_1
XFILLER_69_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_69_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5127_ _5195_/CLK _5127_/D vssd1 vssd1 vccd1 vccd1 _5127_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_29_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5058_ _5062_/CLK _5058_/D vssd1 vssd1 vccd1 vccd1 _5058_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4009_ _4984_/Q _4009_/B vssd1 vssd1 vccd1 vccd1 _4009_/Y sky130_fd_sc_hd__nor2_2
XFILLER_84_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_90_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_90_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_75_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_90_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_71_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2690_ _5286_/Q _3022_/B _5020_/Q _3017_/B vssd1 vssd1 vccd1 vccd1 _3008_/A sky130_fd_sc_hd__o2bb2ai_2
XFILLER_6_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_3 _5003_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_4360_ _4479_/A _4479_/B _4359_/Y vssd1 vssd1 vccd1 vccd1 _4474_/A sky130_fd_sc_hd__o21ai_4
XFILLER_6_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3311_ _3318_/B _3318_/A vssd1 vssd1 vccd1 vccd1 _3311_/X sky130_fd_sc_hd__or2_1
X_4291_ _4291_/A _4301_/A vssd1 vssd1 vccd1 vccd1 _4559_/C sky130_fd_sc_hd__and2_1
XFILLER_3_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3242_ _3243_/A _3243_/B _3243_/C vssd1 vssd1 vccd1 vccd1 _3242_/X sky130_fd_sc_hd__a21o_1
X_3173_ _3726_/B _5182_/Q vssd1 vssd1 vccd1 vccd1 _3174_/B sky130_fd_sc_hd__nand2_1
XFILLER_66_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_66_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_81_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_clk clkbuf_2_0_0_clk/X vssd1 vssd1 vccd1 vccd1 _5195_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_26_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2957_ _2957_/A _2957_/B vssd1 vssd1 vccd1 vccd1 _2958_/B sky130_fd_sc_hd__and2_1
X_2888_ _2888_/A vssd1 vssd1 vccd1 vccd1 _2888_/X sky130_fd_sc_hd__buf_2
X_4627_ _4627_/A _4627_/B vssd1 vssd1 vccd1 vccd1 _4862_/B sky130_fd_sc_hd__nor2_4
X_4558_ _4558_/A _4858_/B vssd1 vssd1 vccd1 vccd1 _4571_/C sky130_fd_sc_hd__nand2_1
X_3509_ _3577_/A _3509_/B _3508_/Y vssd1 vssd1 vccd1 vccd1 _3509_/X sky130_fd_sc_hd__or3b_2
X_4489_ _4814_/A vssd1 vssd1 vccd1 vccd1 _4799_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_89_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_72_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_37_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5283_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_53_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput51 _5195_/Q vssd1 vssd1 vccd1 vccd1 data_out[5] sky130_fd_sc_hd__clkbuf_2
Xoutput40 _5214_/Q vssd1 vssd1 vccd1 vccd1 data_out[24] sky130_fd_sc_hd__clkbuf_2
XFILLER_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_28_clk clkbuf_2_2_0_clk/X vssd1 vssd1 vccd1 vccd1 _5247_/CLK sky130_fd_sc_hd__clkbuf_16
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_72_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3860_ _3860_/A _3860_/B vssd1 vssd1 vccd1 vccd1 _3860_/Y sky130_fd_sc_hd__nand2_1
X_3791_ _3830_/A vssd1 vssd1 vccd1 vccd1 _3791_/X sky130_fd_sc_hd__clkbuf_2
X_2811_ _2811_/A vssd1 vssd1 vccd1 vccd1 _2902_/B sky130_fd_sc_hd__inv_2
XPHY_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2742_ _2742_/A vssd1 vssd1 vccd1 vccd1 _2940_/A sky130_fd_sc_hd__inv_2
XFILLER_8_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4412_ _4412_/A _4412_/B _4778_/A vssd1 vssd1 vccd1 vccd1 _4412_/Y sky130_fd_sc_hd__nand3_1
X_2673_ _2670_/Y _2926_/B _2747_/B vssd1 vssd1 vccd1 vccd1 _2910_/A sky130_fd_sc_hd__a21oi_2
X_4343_ _5101_/Q _5069_/Q vssd1 vssd1 vccd1 vccd1 _4482_/B sky130_fd_sc_hd__nand2_1
X_4274_ _5094_/Q _5062_/Q vssd1 vssd1 vccd1 vccd1 _4525_/A sky130_fd_sc_hd__nor2_1
XFILLER_86_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3225_ _3542_/A _5248_/Q vssd1 vssd1 vccd1 vccd1 _3225_/Y sky130_fd_sc_hd__nand2_1
X_3156_ _3730_/B _5181_/Q vssd1 vssd1 vccd1 vccd1 _3241_/B sky130_fd_sc_hd__and2_1
XFILLER_39_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_82_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xclkbuf_leaf_19_clk clkbuf_opt_0_clk/A vssd1 vssd1 vccd1 vccd1 _5292_/CLK sky130_fd_sc_hd__clkbuf_16
X_3087_ _5257_/Q _3080_/Y _3346_/A _3346_/B vssd1 vssd1 vccd1 vccd1 _3341_/A sky130_fd_sc_hd__o22ai_4
XFILLER_27_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_82_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3989_ _5000_/Q _5000_/D vssd1 vssd1 vccd1 vccd1 _3990_/C sky130_fd_sc_hd__xnor2_2
XFILLER_77_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3010_ _3010_/A _3010_/B _3010_/C vssd1 vssd1 vccd1 vccd1 _3012_/A sky130_fd_sc_hd__or3_2
XFILLER_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4961_ _5124_/Q _4961_/B vssd1 vssd1 vccd1 vccd1 _4963_/A sky130_fd_sc_hd__nor2_1
XFILLER_17_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3912_ _5118_/Q vssd1 vssd1 vccd1 vccd1 _3913_/B sky130_fd_sc_hd__inv_2
X_4892_ _4892_/A _4898_/B _5018_/Q vssd1 vssd1 vccd1 vccd1 _4912_/A sky130_fd_sc_hd__and3_1
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3843_ _3843_/A vssd1 vssd1 vccd1 vccd1 _3911_/A sky130_fd_sc_hd__clkbuf_4
X_3774_ _5165_/Q _3768_/X _3762_/X _3773_/Y vssd1 vssd1 vccd1 vccd1 _5165_/D sky130_fd_sc_hd__o211a_1
X_2725_ _2685_/Y _2716_/Y _2724_/Y vssd1 vssd1 vccd1 vccd1 _2943_/A sky130_fd_sc_hd__o21bai_1
X_2656_ _5311_/Q _4704_/A vssd1 vssd1 vccd1 vccd1 _2772_/A sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_8_clk clkbuf_2_1_0_clk/X vssd1 vssd1 vccd1 vccd1 _5097_/CLK sky130_fd_sc_hd__clkbuf_16
X_2587_ _2605_/A vssd1 vssd1 vccd1 vccd1 _2602_/A sky130_fd_sc_hd__buf_1
X_4326_ _4326_/A _4661_/B vssd1 vssd1 vccd1 vccd1 _4328_/A sky130_fd_sc_hd__nand2_1
X_4257_ _5072_/Q vssd1 vssd1 vccd1 vccd1 _4601_/B sky130_fd_sc_hd__inv_2
X_3208_ _3262_/A vssd1 vssd1 vccd1 vccd1 _3208_/X sky130_fd_sc_hd__clkbuf_2
X_4188_ _4194_/A _5092_/Q _4180_/C _4169_/A vssd1 vssd1 vccd1 vccd1 _4188_/Y sky130_fd_sc_hd__a31oi_1
X_3139_ _3138_/Y _3132_/A _3133_/A vssd1 vssd1 vccd1 vccd1 _3257_/B sky130_fd_sc_hd__a21oi_2
XFILLER_82_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_82_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3490_ _3575_/A _3575_/B _3489_/X vssd1 vssd1 vccd1 vccd1 _3490_/Y sky130_fd_sc_hd__a21oi_2
X_2510_ _4807_/A vssd1 vssd1 vccd1 vccd1 _2510_/X sky130_fd_sc_hd__buf_2
XFILLER_5_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5160_ _5274_/CLK _5160_/D vssd1 vssd1 vccd1 vccd1 _5160_/Q sky130_fd_sc_hd__dfxtp_2
X_5091_ _5097_/CLK _5091_/D vssd1 vssd1 vccd1 vccd1 _5091_/Q sky130_fd_sc_hd__dfxtp_1
X_4111_ _4180_/A vssd1 vssd1 vccd1 vccd1 _4111_/X sky130_fd_sc_hd__clkbuf_2
X_4042_ _4045_/C _4041_/A _4040_/A _4040_/B vssd1 vssd1 vccd1 vccd1 _4054_/A sky130_fd_sc_hd__o2bb2ai_4
XFILLER_68_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_83_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4944_ _4944_/A _5120_/Q vssd1 vssd1 vccd1 vccd1 _4948_/B sky130_fd_sc_hd__nand2_1
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4875_ _4875_/A vssd1 vssd1 vccd1 vccd1 _4881_/A sky130_fd_sc_hd__inv_2
X_3826_ _3833_/A _3826_/B vssd1 vssd1 vccd1 vccd1 _3826_/Y sky130_fd_sc_hd__nand2_1
X_3757_ _5171_/Q _3754_/X _3749_/X _3756_/Y vssd1 vssd1 vccd1 vccd1 _5171_/D sky130_fd_sc_hd__o211a_1
X_2708_ _2687_/Y _2989_/A _2798_/A _2707_/Y vssd1 vssd1 vccd1 vccd1 _2708_/Y sky130_fd_sc_hd__o211ai_1
X_3688_ _3687_/B _3687_/A _3642_/X vssd1 vssd1 vccd1 vccd1 _3688_/X sky130_fd_sc_hd__a21o_1
XFILLER_3_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2639_ _2995_/A _3017_/B vssd1 vssd1 vccd1 vccd1 _2639_/Y sky130_fd_sc_hd__nand2_1
XFILLER_87_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_4309_ _5059_/Q vssd1 vssd1 vccd1 vccd1 _4648_/B sky130_fd_sc_hd__inv_2
X_5289_ _5292_/CLK _5289_/D vssd1 vssd1 vccd1 vccd1 _5289_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_47_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_67_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2990_ _5291_/Q _4863_/A vssd1 vssd1 vccd1 vccd1 _2991_/A sky130_fd_sc_hd__nor2_1
XFILLER_61_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4660_ _4830_/A _4830_/B _4659_/X vssd1 vssd1 vccd1 vccd1 _4821_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3611_ _3611_/A _3611_/B vssd1 vssd1 vccd1 vccd1 _3611_/Y sky130_fd_sc_hd__nor2_1
X_4591_ _4591_/A _4591_/B vssd1 vssd1 vccd1 vccd1 _4728_/B sky130_fd_sc_hd__nor2_1
X_3542_ _3542_/A _5220_/Q vssd1 vssd1 vccd1 vccd1 _3542_/Y sky130_fd_sc_hd__nand2_1
X_3473_ _3628_/A _3628_/B _3635_/B vssd1 vssd1 vccd1 vccd1 _3473_/X sky130_fd_sc_hd__or3_1
XFILLER_69_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5212_ _5236_/CLK _5212_/D vssd1 vssd1 vccd1 vccd1 _5212_/Q sky130_fd_sc_hd__dfxtp_1
X_5143_ _5228_/CLK _5143_/D vssd1 vssd1 vccd1 vccd1 _5143_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_56_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_5074_ _5076_/CLK _5074_/D vssd1 vssd1 vccd1 vccd1 _5074_/Q sky130_fd_sc_hd__dfxtp_1
X_4025_ _4056_/C _4055_/A _4048_/B vssd1 vssd1 vccd1 vccd1 _4063_/B sky130_fd_sc_hd__nand3_4
XFILLER_37_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_71_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_4927_ _4927_/A _4927_/B vssd1 vssd1 vccd1 vccd1 _4932_/A sky130_fd_sc_hd__and2_1
XFILLER_52_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4858_ _4872_/A _4858_/B vssd1 vssd1 vccd1 vccd1 _4871_/C sky130_fd_sc_hd__nand2_1
XFILLER_60_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3809_ _3822_/A vssd1 vssd1 vccd1 vccd1 _3809_/X sky130_fd_sc_hd__clkbuf_2
X_4789_ _3879_/X _4787_/Y _4540_/X _4788_/Y vssd1 vssd1 vccd1 vccd1 _5039_/D sky130_fd_sc_hd__o211a_1
XFILLER_4_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_87_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_87_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_85_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_75_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_70_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_78_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2973_ _2973_/A _2973_/B vssd1 vssd1 vccd1 vccd1 _2973_/X sky130_fd_sc_hd__xor2_1
X_4712_ _5046_/Q _5078_/Q vssd1 vssd1 vccd1 vccd1 _4720_/A sky130_fd_sc_hd__nor2_1
X_4643_ _4643_/A _4643_/B vssd1 vssd1 vccd1 vccd1 _4644_/A sky130_fd_sc_hd__nand2_1
X_4574_ _4770_/A vssd1 vssd1 vccd1 vccd1 _4574_/X sky130_fd_sc_hd__buf_2
X_3525_ _3800_/B _5155_/Q _3521_/Y _3524_/Y vssd1 vssd1 vccd1 vccd1 _3525_/Y sky130_fd_sc_hd__a22oi_4
X_3456_ _3658_/B _3651_/A vssd1 vssd1 vccd1 vccd1 _3456_/X sky130_fd_sc_hd__or2_1
XFILLER_69_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3387_ _5249_/Q vssd1 vssd1 vccd1 vccd1 _3805_/B sky130_fd_sc_hd__inv_2
XFILLER_57_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_5126_ _5197_/CLK _5126_/D vssd1 vssd1 vccd1 vccd1 _5126_/Q sky130_fd_sc_hd__dfxtp_1
X_5057_ _5062_/CLK _5057_/D vssd1 vssd1 vccd1 vccd1 _5057_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_4008_ _4009_/B _4984_/Q vssd1 vssd1 vccd1 vccd1 _4008_/X sky130_fd_sc_hd__and2_1
XFILLER_44_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold40 input1/X vssd1 vssd1 vccd1 vccd1 hold40/X sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_75_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_4 _5003_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3310_ _3310_/A _3310_/B vssd1 vssd1 vccd1 vccd1 _3318_/A sky130_fd_sc_hd__and2_1
X_4290_ _5087_/Q _5055_/Q vssd1 vssd1 vccd1 vccd1 _4301_/A sky130_fd_sc_hd__nand2_1
XFILLER_3_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_79_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3241_ _3241_/A _3241_/B vssd1 vssd1 vccd1 vccd1 _3243_/C sky130_fd_sc_hd__nor2_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3172_ _3223_/A _3172_/B vssd1 vssd1 vccd1 vccd1 _3178_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_81_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2956_ _2957_/A _2958_/A _2957_/B _2901_/A vssd1 vssd1 vccd1 vccd1 _2956_/X sky130_fd_sc_hd__a31o_1
XFILLER_22_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2887_ _2884_/X _2760_/A _2885_/Y _2848_/X vssd1 vssd1 vccd1 vccd1 _2887_/X sky130_fd_sc_hd__a31o_1
XFILLER_30_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_4626_ _4863_/A _4626_/B vssd1 vssd1 vccd1 vccd1 _4627_/B sky130_fd_sc_hd__nor2_2
X_4557_ _5054_/Q vssd1 vssd1 vccd1 vccd1 _4858_/B sky130_fd_sc_hd__inv_2
X_3508_ _3512_/A _3508_/B vssd1 vssd1 vccd1 vccd1 _3508_/Y sky130_fd_sc_hd__nor2_1
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4488_ _4798_/A _4488_/B _4482_/A vssd1 vssd1 vccd1 vccd1 _4488_/X sky130_fd_sc_hd__or3b_1
X_3439_ _3681_/A _3685_/A _3681_/B vssd1 vssd1 vccd1 vccd1 _3673_/A sky130_fd_sc_hd__a21oi_4
XFILLER_57_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_5109_ _5109_/CLK _5109_/D vssd1 vssd1 vccd1 vccd1 _5109_/Q sky130_fd_sc_hd__dfxtp_1
XFILLER_57_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_72_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput30 _5205_/Q vssd1 vssd1 vccd1 vccd1 data_out[15] sky130_fd_sc_hd__clkbuf_2
Xoutput52 _5196_/Q vssd1 vssd1 vccd1 vccd1 data_out[6] sky130_fd_sc_hd__clkbuf_2
Xoutput41 _5215_/Q vssd1 vssd1 vccd1 vccd1 data_out[25] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3790_ _5159_/Q _3783_/X _3778_/X _3789_/Y vssd1 vssd1 vccd1 vccd1 _5159_/D sky130_fd_sc_hd__o211a_1
X_2810_ _2908_/A _2908_/B _2750_/X vssd1 vssd1 vccd1 vccd1 _2902_/A sky130_fd_sc_hd__o21bai_2
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2741_ _2936_/B _2741_/B vssd1 vssd1 vccd1 vccd1 _2742_/A sky130_fd_sc_hd__nand2_1
XFILLER_8_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_4411_ _4241_/Y _4411_/B _4411_/C vssd1 vssd1 vccd1 vccd1 _4412_/B sky130_fd_sc_hd__nand3b_1
X_2672_ _4682_/A _5303_/Q vssd1 vssd1 vccd1 vccd1 _2747_/B sky130_fd_sc_hd__and2_1
X_4342_ _4342_/A _4691_/B vssd1 vssd1 vccd1 vccd1 _4344_/A sky130_fd_sc_hd__nand2_1
X_4273_ _4504_/A _4506_/B _4504_/B vssd1 vssd1 vccd1 vccd1 _4479_/A sky130_fd_sc_hd__o21bai_2
XFILLER_86_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3224_ _3224_/A _3563_/B _3224_/C vssd1 vssd1 vccd1 vccd1 _3224_/Y sky130_fd_sc_hd__nand3_1
.ends

