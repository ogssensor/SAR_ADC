magic
tech sky130A
magscale 1 2
timestamp 1622831649
<< obsli1 >>
rect 1104 1853 178848 117521
<< obsm1 >>
rect 658 892 179294 119672
<< metal2 >>
rect 662 119200 718 120000
rect 2042 119200 2098 120000
rect 3422 119200 3478 120000
rect 4894 119200 4950 120000
rect 6274 119200 6330 120000
rect 7746 119200 7802 120000
rect 9126 119200 9182 120000
rect 10506 119200 10562 120000
rect 11978 119200 12034 120000
rect 13358 119200 13414 120000
rect 14830 119200 14886 120000
rect 16210 119200 16266 120000
rect 17590 119200 17646 120000
rect 19062 119200 19118 120000
rect 20442 119200 20498 120000
rect 21914 119200 21970 120000
rect 23294 119200 23350 120000
rect 24674 119200 24730 120000
rect 26146 119200 26202 120000
rect 27526 119200 27582 120000
rect 28998 119200 29054 120000
rect 30378 119200 30434 120000
rect 31850 119200 31906 120000
rect 33230 119200 33286 120000
rect 34610 119200 34666 120000
rect 36082 119200 36138 120000
rect 37462 119200 37518 120000
rect 38934 119200 38990 120000
rect 40314 119200 40370 120000
rect 41694 119200 41750 120000
rect 43166 119200 43222 120000
rect 44546 119200 44602 120000
rect 46018 119200 46074 120000
rect 47398 119200 47454 120000
rect 48778 119200 48834 120000
rect 50250 119200 50306 120000
rect 51630 119200 51686 120000
rect 53102 119200 53158 120000
rect 54482 119200 54538 120000
rect 55862 119200 55918 120000
rect 57334 119200 57390 120000
rect 58714 119200 58770 120000
rect 60186 119200 60242 120000
rect 61566 119200 61622 120000
rect 63038 119200 63094 120000
rect 64418 119200 64474 120000
rect 65798 119200 65854 120000
rect 67270 119200 67326 120000
rect 68650 119200 68706 120000
rect 70122 119200 70178 120000
rect 71502 119200 71558 120000
rect 72882 119200 72938 120000
rect 74354 119200 74410 120000
rect 75734 119200 75790 120000
rect 77206 119200 77262 120000
rect 78586 119200 78642 120000
rect 79966 119200 80022 120000
rect 81438 119200 81494 120000
rect 82818 119200 82874 120000
rect 84290 119200 84346 120000
rect 85670 119200 85726 120000
rect 87050 119200 87106 120000
rect 88522 119200 88578 120000
rect 89902 119200 89958 120000
rect 91374 119200 91430 120000
rect 92754 119200 92810 120000
rect 94226 119200 94282 120000
rect 95606 119200 95662 120000
rect 96986 119200 97042 120000
rect 98458 119200 98514 120000
rect 99838 119200 99894 120000
rect 101310 119200 101366 120000
rect 102690 119200 102746 120000
rect 104070 119200 104126 120000
rect 105542 119200 105598 120000
rect 106922 119200 106978 120000
rect 108394 119200 108450 120000
rect 109774 119200 109830 120000
rect 111154 119200 111210 120000
rect 112626 119200 112682 120000
rect 114006 119200 114062 120000
rect 115478 119200 115534 120000
rect 116858 119200 116914 120000
rect 118238 119200 118294 120000
rect 119710 119200 119766 120000
rect 121090 119200 121146 120000
rect 122562 119200 122618 120000
rect 123942 119200 123998 120000
rect 125414 119200 125470 120000
rect 126794 119200 126850 120000
rect 128174 119200 128230 120000
rect 129646 119200 129702 120000
rect 131026 119200 131082 120000
rect 132498 119200 132554 120000
rect 133878 119200 133934 120000
rect 135258 119200 135314 120000
rect 136730 119200 136786 120000
rect 138110 119200 138166 120000
rect 139582 119200 139638 120000
rect 140962 119200 141018 120000
rect 142342 119200 142398 120000
rect 143814 119200 143870 120000
rect 145194 119200 145250 120000
rect 146666 119200 146722 120000
rect 148046 119200 148102 120000
rect 149426 119200 149482 120000
rect 150898 119200 150954 120000
rect 152278 119200 152334 120000
rect 153750 119200 153806 120000
rect 155130 119200 155186 120000
rect 156602 119200 156658 120000
rect 157982 119200 158038 120000
rect 159362 119200 159418 120000
rect 160834 119200 160890 120000
rect 162214 119200 162270 120000
rect 163686 119200 163742 120000
rect 165066 119200 165122 120000
rect 166446 119200 166502 120000
rect 167918 119200 167974 120000
rect 169298 119200 169354 120000
rect 170770 119200 170826 120000
rect 172150 119200 172206 120000
rect 173530 119200 173586 120000
rect 175002 119200 175058 120000
rect 176382 119200 176438 120000
rect 177854 119200 177910 120000
rect 179234 119200 179290 120000
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5906 0 5962 800
rect 7562 0 7618 800
rect 9310 0 9366 800
rect 10966 0 11022 800
rect 12714 0 12770 800
rect 14370 0 14426 800
rect 16118 0 16174 800
rect 17774 0 17830 800
rect 19522 0 19578 800
rect 21178 0 21234 800
rect 22926 0 22982 800
rect 24582 0 24638 800
rect 26238 0 26294 800
rect 27986 0 28042 800
rect 29642 0 29698 800
rect 31390 0 31446 800
rect 33046 0 33102 800
rect 34794 0 34850 800
rect 36450 0 36506 800
rect 38198 0 38254 800
rect 39854 0 39910 800
rect 41602 0 41658 800
rect 43258 0 43314 800
rect 45006 0 45062 800
rect 46662 0 46718 800
rect 48318 0 48374 800
rect 50066 0 50122 800
rect 51722 0 51778 800
rect 53470 0 53526 800
rect 55126 0 55182 800
rect 56874 0 56930 800
rect 58530 0 58586 800
rect 60278 0 60334 800
rect 61934 0 61990 800
rect 63682 0 63738 800
rect 65338 0 65394 800
rect 67086 0 67142 800
rect 68742 0 68798 800
rect 70398 0 70454 800
rect 72146 0 72202 800
rect 73802 0 73858 800
rect 75550 0 75606 800
rect 77206 0 77262 800
rect 78954 0 79010 800
rect 80610 0 80666 800
rect 82358 0 82414 800
rect 84014 0 84070 800
rect 85762 0 85818 800
rect 87418 0 87474 800
rect 89166 0 89222 800
rect 90822 0 90878 800
rect 92478 0 92534 800
rect 94226 0 94282 800
rect 95882 0 95938 800
rect 97630 0 97686 800
rect 99286 0 99342 800
rect 101034 0 101090 800
rect 102690 0 102746 800
rect 104438 0 104494 800
rect 106094 0 106150 800
rect 107842 0 107898 800
rect 109498 0 109554 800
rect 111246 0 111302 800
rect 112902 0 112958 800
rect 114558 0 114614 800
rect 116306 0 116362 800
rect 117962 0 118018 800
rect 119710 0 119766 800
rect 121366 0 121422 800
rect 123114 0 123170 800
rect 124770 0 124826 800
rect 126518 0 126574 800
rect 128174 0 128230 800
rect 129922 0 129978 800
rect 131578 0 131634 800
rect 133326 0 133382 800
rect 134982 0 135038 800
rect 136638 0 136694 800
rect 138386 0 138442 800
rect 140042 0 140098 800
rect 141790 0 141846 800
rect 143446 0 143502 800
rect 145194 0 145250 800
rect 146850 0 146906 800
rect 148598 0 148654 800
rect 150254 0 150310 800
rect 152002 0 152058 800
rect 153658 0 153714 800
rect 155406 0 155462 800
rect 157062 0 157118 800
rect 158718 0 158774 800
rect 160466 0 160522 800
rect 162122 0 162178 800
rect 163870 0 163926 800
rect 165526 0 165582 800
rect 167274 0 167330 800
rect 168930 0 168986 800
rect 170678 0 170734 800
rect 172334 0 172390 800
rect 174082 0 174138 800
rect 175738 0 175794 800
rect 177486 0 177542 800
rect 179142 0 179198 800
<< obsm2 >>
rect 774 119144 1986 119785
rect 2154 119144 3366 119785
rect 3534 119144 4838 119785
rect 5006 119144 6218 119785
rect 6386 119144 7690 119785
rect 7858 119144 9070 119785
rect 9238 119144 10450 119785
rect 10618 119144 11922 119785
rect 12090 119144 13302 119785
rect 13470 119144 14774 119785
rect 14942 119144 16154 119785
rect 16322 119144 17534 119785
rect 17702 119144 19006 119785
rect 19174 119144 20386 119785
rect 20554 119144 21858 119785
rect 22026 119144 23238 119785
rect 23406 119144 24618 119785
rect 24786 119144 26090 119785
rect 26258 119144 27470 119785
rect 27638 119144 28942 119785
rect 29110 119144 30322 119785
rect 30490 119144 31794 119785
rect 31962 119144 33174 119785
rect 33342 119144 34554 119785
rect 34722 119144 36026 119785
rect 36194 119144 37406 119785
rect 37574 119144 38878 119785
rect 39046 119144 40258 119785
rect 40426 119144 41638 119785
rect 41806 119144 43110 119785
rect 43278 119144 44490 119785
rect 44658 119144 45962 119785
rect 46130 119144 47342 119785
rect 47510 119144 48722 119785
rect 48890 119144 50194 119785
rect 50362 119144 51574 119785
rect 51742 119144 53046 119785
rect 53214 119144 54426 119785
rect 54594 119144 55806 119785
rect 55974 119144 57278 119785
rect 57446 119144 58658 119785
rect 58826 119144 60130 119785
rect 60298 119144 61510 119785
rect 61678 119144 62982 119785
rect 63150 119144 64362 119785
rect 64530 119144 65742 119785
rect 65910 119144 67214 119785
rect 67382 119144 68594 119785
rect 68762 119144 70066 119785
rect 70234 119144 71446 119785
rect 71614 119144 72826 119785
rect 72994 119144 74298 119785
rect 74466 119144 75678 119785
rect 75846 119144 77150 119785
rect 77318 119144 78530 119785
rect 78698 119144 79910 119785
rect 80078 119144 81382 119785
rect 81550 119144 82762 119785
rect 82930 119144 84234 119785
rect 84402 119144 85614 119785
rect 85782 119144 86994 119785
rect 87162 119144 88466 119785
rect 88634 119144 89846 119785
rect 90014 119144 91318 119785
rect 91486 119144 92698 119785
rect 92866 119144 94170 119785
rect 94338 119144 95550 119785
rect 95718 119144 96930 119785
rect 97098 119144 98402 119785
rect 98570 119144 99782 119785
rect 99950 119144 101254 119785
rect 101422 119144 102634 119785
rect 102802 119144 104014 119785
rect 104182 119144 105486 119785
rect 105654 119144 106866 119785
rect 107034 119144 108338 119785
rect 108506 119144 109718 119785
rect 109886 119144 111098 119785
rect 111266 119144 112570 119785
rect 112738 119144 113950 119785
rect 114118 119144 115422 119785
rect 115590 119144 116802 119785
rect 116970 119144 118182 119785
rect 118350 119144 119654 119785
rect 119822 119144 121034 119785
rect 121202 119144 122506 119785
rect 122674 119144 123886 119785
rect 124054 119144 125358 119785
rect 125526 119144 126738 119785
rect 126906 119144 128118 119785
rect 128286 119144 129590 119785
rect 129758 119144 130970 119785
rect 131138 119144 132442 119785
rect 132610 119144 133822 119785
rect 133990 119144 135202 119785
rect 135370 119144 136674 119785
rect 136842 119144 138054 119785
rect 138222 119144 139526 119785
rect 139694 119144 140906 119785
rect 141074 119144 142286 119785
rect 142454 119144 143758 119785
rect 143926 119144 145138 119785
rect 145306 119144 146610 119785
rect 146778 119144 147990 119785
rect 148158 119144 149370 119785
rect 149538 119144 150842 119785
rect 151010 119144 152222 119785
rect 152390 119144 153694 119785
rect 153862 119144 155074 119785
rect 155242 119144 156546 119785
rect 156714 119144 157926 119785
rect 158094 119144 159306 119785
rect 159474 119144 160778 119785
rect 160946 119144 162158 119785
rect 162326 119144 163630 119785
rect 163798 119144 165010 119785
rect 165178 119144 166390 119785
rect 166558 119144 167862 119785
rect 168030 119144 169242 119785
rect 169410 119144 170714 119785
rect 170882 119144 172094 119785
rect 172262 119144 173474 119785
rect 173642 119144 174946 119785
rect 175114 119144 176326 119785
rect 176494 119144 177798 119785
rect 177966 119144 179178 119785
rect 664 856 179288 119144
rect 664 167 790 856
rect 958 167 2446 856
rect 2614 167 4102 856
rect 4270 167 5850 856
rect 6018 167 7506 856
rect 7674 167 9254 856
rect 9422 167 10910 856
rect 11078 167 12658 856
rect 12826 167 14314 856
rect 14482 167 16062 856
rect 16230 167 17718 856
rect 17886 167 19466 856
rect 19634 167 21122 856
rect 21290 167 22870 856
rect 23038 167 24526 856
rect 24694 167 26182 856
rect 26350 167 27930 856
rect 28098 167 29586 856
rect 29754 167 31334 856
rect 31502 167 32990 856
rect 33158 167 34738 856
rect 34906 167 36394 856
rect 36562 167 38142 856
rect 38310 167 39798 856
rect 39966 167 41546 856
rect 41714 167 43202 856
rect 43370 167 44950 856
rect 45118 167 46606 856
rect 46774 167 48262 856
rect 48430 167 50010 856
rect 50178 167 51666 856
rect 51834 167 53414 856
rect 53582 167 55070 856
rect 55238 167 56818 856
rect 56986 167 58474 856
rect 58642 167 60222 856
rect 60390 167 61878 856
rect 62046 167 63626 856
rect 63794 167 65282 856
rect 65450 167 67030 856
rect 67198 167 68686 856
rect 68854 167 70342 856
rect 70510 167 72090 856
rect 72258 167 73746 856
rect 73914 167 75494 856
rect 75662 167 77150 856
rect 77318 167 78898 856
rect 79066 167 80554 856
rect 80722 167 82302 856
rect 82470 167 83958 856
rect 84126 167 85706 856
rect 85874 167 87362 856
rect 87530 167 89110 856
rect 89278 167 90766 856
rect 90934 167 92422 856
rect 92590 167 94170 856
rect 94338 167 95826 856
rect 95994 167 97574 856
rect 97742 167 99230 856
rect 99398 167 100978 856
rect 101146 167 102634 856
rect 102802 167 104382 856
rect 104550 167 106038 856
rect 106206 167 107786 856
rect 107954 167 109442 856
rect 109610 167 111190 856
rect 111358 167 112846 856
rect 113014 167 114502 856
rect 114670 167 116250 856
rect 116418 167 117906 856
rect 118074 167 119654 856
rect 119822 167 121310 856
rect 121478 167 123058 856
rect 123226 167 124714 856
rect 124882 167 126462 856
rect 126630 167 128118 856
rect 128286 167 129866 856
rect 130034 167 131522 856
rect 131690 167 133270 856
rect 133438 167 134926 856
rect 135094 167 136582 856
rect 136750 167 138330 856
rect 138498 167 139986 856
rect 140154 167 141734 856
rect 141902 167 143390 856
rect 143558 167 145138 856
rect 145306 167 146794 856
rect 146962 167 148542 856
rect 148710 167 150198 856
rect 150366 167 151946 856
rect 152114 167 153602 856
rect 153770 167 155350 856
rect 155518 167 157006 856
rect 157174 167 158662 856
rect 158830 167 160410 856
rect 160578 167 162066 856
rect 162234 167 163814 856
rect 163982 167 165470 856
rect 165638 167 167218 856
rect 167386 167 168874 856
rect 169042 167 170622 856
rect 170790 167 172278 856
rect 172446 167 174026 856
rect 174194 167 175682 856
rect 175850 167 177430 856
rect 177598 167 179086 856
rect 179254 167 179288 856
<< metal3 >>
rect 0 119688 800 119808
rect 0 119416 800 119536
rect 0 119144 800 119264
rect 0 118736 800 118856
rect 0 118464 800 118584
rect 0 118192 800 118312
rect 0 117784 800 117904
rect 0 117512 800 117632
rect 0 117240 800 117360
rect 0 116968 800 117088
rect 0 116560 800 116680
rect 0 116288 800 116408
rect 0 116016 800 116136
rect 0 115608 800 115728
rect 0 115336 800 115456
rect 0 115064 800 115184
rect 0 114656 800 114776
rect 0 114384 800 114504
rect 0 114112 800 114232
rect 0 113840 800 113960
rect 0 113432 800 113552
rect 0 113160 800 113280
rect 0 112888 800 113008
rect 0 112480 800 112600
rect 0 112208 800 112328
rect 0 111936 800 112056
rect 0 111528 800 111648
rect 0 111256 800 111376
rect 0 110984 800 111104
rect 0 110712 800 110832
rect 0 110304 800 110424
rect 0 110032 800 110152
rect 0 109760 800 109880
rect 0 109352 800 109472
rect 0 109080 800 109200
rect 0 108808 800 108928
rect 0 108536 800 108656
rect 0 108128 800 108248
rect 0 107856 800 107976
rect 0 107584 800 107704
rect 0 107176 800 107296
rect 0 106904 800 107024
rect 0 106632 800 106752
rect 0 106224 800 106344
rect 0 105952 800 106072
rect 0 105680 800 105800
rect 0 105408 800 105528
rect 0 105000 800 105120
rect 0 104728 800 104848
rect 0 104456 800 104576
rect 0 104048 800 104168
rect 0 103776 800 103896
rect 0 103504 800 103624
rect 0 103096 800 103216
rect 0 102824 800 102944
rect 0 102552 800 102672
rect 0 102280 800 102400
rect 0 101872 800 101992
rect 0 101600 800 101720
rect 0 101328 800 101448
rect 0 100920 800 101040
rect 0 100648 800 100768
rect 0 100376 800 100496
rect 0 100104 800 100224
rect 0 99696 800 99816
rect 0 99424 800 99544
rect 0 99152 800 99272
rect 0 98744 800 98864
rect 0 98472 800 98592
rect 0 98200 800 98320
rect 0 97792 800 97912
rect 0 97520 800 97640
rect 0 97248 800 97368
rect 0 96976 800 97096
rect 0 96568 800 96688
rect 0 96296 800 96416
rect 0 96024 800 96144
rect 0 95616 800 95736
rect 0 95344 800 95464
rect 0 95072 800 95192
rect 0 94664 800 94784
rect 0 94392 800 94512
rect 0 94120 800 94240
rect 0 93848 800 93968
rect 0 93440 800 93560
rect 0 93168 800 93288
rect 0 92896 800 93016
rect 0 92488 800 92608
rect 0 92216 800 92336
rect 0 91944 800 92064
rect 0 91536 800 91656
rect 0 91264 800 91384
rect 0 90992 800 91112
rect 0 90720 800 90840
rect 0 90312 800 90432
rect 0 90040 800 90160
rect 0 89768 800 89888
rect 0 89360 800 89480
rect 0 89088 800 89208
rect 0 88816 800 88936
rect 0 88544 800 88664
rect 0 88136 800 88256
rect 0 87864 800 87984
rect 0 87592 800 87712
rect 0 87184 800 87304
rect 0 86912 800 87032
rect 0 86640 800 86760
rect 0 86232 800 86352
rect 0 85960 800 86080
rect 0 85688 800 85808
rect 0 85416 800 85536
rect 0 85008 800 85128
rect 0 84736 800 84856
rect 0 84464 800 84584
rect 0 84056 800 84176
rect 0 83784 800 83904
rect 0 83512 800 83632
rect 0 83104 800 83224
rect 0 82832 800 82952
rect 0 82560 800 82680
rect 0 82288 800 82408
rect 0 81880 800 82000
rect 0 81608 800 81728
rect 0 81336 800 81456
rect 0 80928 800 81048
rect 0 80656 800 80776
rect 0 80384 800 80504
rect 0 80112 800 80232
rect 0 79704 800 79824
rect 0 79432 800 79552
rect 0 79160 800 79280
rect 0 78752 800 78872
rect 0 78480 800 78600
rect 0 78208 800 78328
rect 0 77800 800 77920
rect 0 77528 800 77648
rect 0 77256 800 77376
rect 0 76984 800 77104
rect 0 76576 800 76696
rect 0 76304 800 76424
rect 0 76032 800 76152
rect 0 75624 800 75744
rect 0 75352 800 75472
rect 0 75080 800 75200
rect 0 74672 800 74792
rect 0 74400 800 74520
rect 0 74128 800 74248
rect 0 73856 800 73976
rect 0 73448 800 73568
rect 0 73176 800 73296
rect 0 72904 800 73024
rect 0 72496 800 72616
rect 0 72224 800 72344
rect 0 71952 800 72072
rect 0 71544 800 71664
rect 0 71272 800 71392
rect 0 71000 800 71120
rect 0 70728 800 70848
rect 0 70320 800 70440
rect 0 70048 800 70168
rect 0 69776 800 69896
rect 0 69368 800 69488
rect 0 69096 800 69216
rect 0 68824 800 68944
rect 0 68552 800 68672
rect 0 68144 800 68264
rect 0 67872 800 67992
rect 0 67600 800 67720
rect 0 67192 800 67312
rect 0 66920 800 67040
rect 0 66648 800 66768
rect 0 66240 800 66360
rect 0 65968 800 66088
rect 0 65696 800 65816
rect 0 65424 800 65544
rect 0 65016 800 65136
rect 0 64744 800 64864
rect 0 64472 800 64592
rect 0 64064 800 64184
rect 0 63792 800 63912
rect 0 63520 800 63640
rect 0 63112 800 63232
rect 0 62840 800 62960
rect 0 62568 800 62688
rect 0 62296 800 62416
rect 0 61888 800 62008
rect 0 61616 800 61736
rect 0 61344 800 61464
rect 0 60936 800 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 179200 59984 180000 60104
rect 0 59712 800 59832
rect 0 59440 800 59560
rect 0 59168 800 59288
rect 0 58760 800 58880
rect 0 58488 800 58608
rect 0 58216 800 58336
rect 0 57808 800 57928
rect 0 57536 800 57656
rect 0 57264 800 57384
rect 0 56992 800 57112
rect 0 56584 800 56704
rect 0 56312 800 56432
rect 0 56040 800 56160
rect 0 55632 800 55752
rect 0 55360 800 55480
rect 0 55088 800 55208
rect 0 54680 800 54800
rect 0 54408 800 54528
rect 0 54136 800 54256
rect 0 53864 800 53984
rect 0 53456 800 53576
rect 0 53184 800 53304
rect 0 52912 800 53032
rect 0 52504 800 52624
rect 0 52232 800 52352
rect 0 51960 800 52080
rect 0 51552 800 51672
rect 0 51280 800 51400
rect 0 51008 800 51128
rect 0 50736 800 50856
rect 0 50328 800 50448
rect 0 50056 800 50176
rect 0 49784 800 49904
rect 0 49376 800 49496
rect 0 49104 800 49224
rect 0 48832 800 48952
rect 0 48560 800 48680
rect 0 48152 800 48272
rect 0 47880 800 48000
rect 0 47608 800 47728
rect 0 47200 800 47320
rect 0 46928 800 47048
rect 0 46656 800 46776
rect 0 46248 800 46368
rect 0 45976 800 46096
rect 0 45704 800 45824
rect 0 45432 800 45552
rect 0 45024 800 45144
rect 0 44752 800 44872
rect 0 44480 800 44600
rect 0 44072 800 44192
rect 0 43800 800 43920
rect 0 43528 800 43648
rect 0 43120 800 43240
rect 0 42848 800 42968
rect 0 42576 800 42696
rect 0 42304 800 42424
rect 0 41896 800 42016
rect 0 41624 800 41744
rect 0 41352 800 41472
rect 0 40944 800 41064
rect 0 40672 800 40792
rect 0 40400 800 40520
rect 0 40128 800 40248
rect 0 39720 800 39840
rect 0 39448 800 39568
rect 0 39176 800 39296
rect 0 38768 800 38888
rect 0 38496 800 38616
rect 0 38224 800 38344
rect 0 37816 800 37936
rect 0 37544 800 37664
rect 0 37272 800 37392
rect 0 37000 800 37120
rect 0 36592 800 36712
rect 0 36320 800 36440
rect 0 36048 800 36168
rect 0 35640 800 35760
rect 0 35368 800 35488
rect 0 35096 800 35216
rect 0 34688 800 34808
rect 0 34416 800 34536
rect 0 34144 800 34264
rect 0 33872 800 33992
rect 0 33464 800 33584
rect 0 33192 800 33312
rect 0 32920 800 33040
rect 0 32512 800 32632
rect 0 32240 800 32360
rect 0 31968 800 32088
rect 0 31560 800 31680
rect 0 31288 800 31408
rect 0 31016 800 31136
rect 0 30744 800 30864
rect 0 30336 800 30456
rect 0 30064 800 30184
rect 0 29792 800 29912
rect 0 29384 800 29504
rect 0 29112 800 29232
rect 0 28840 800 28960
rect 0 28568 800 28688
rect 0 28160 800 28280
rect 0 27888 800 28008
rect 0 27616 800 27736
rect 0 27208 800 27328
rect 0 26936 800 27056
rect 0 26664 800 26784
rect 0 26256 800 26376
rect 0 25984 800 26104
rect 0 25712 800 25832
rect 0 25440 800 25560
rect 0 25032 800 25152
rect 0 24760 800 24880
rect 0 24488 800 24608
rect 0 24080 800 24200
rect 0 23808 800 23928
rect 0 23536 800 23656
rect 0 23128 800 23248
rect 0 22856 800 22976
rect 0 22584 800 22704
rect 0 22312 800 22432
rect 0 21904 800 22024
rect 0 21632 800 21752
rect 0 21360 800 21480
rect 0 20952 800 21072
rect 0 20680 800 20800
rect 0 20408 800 20528
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19456 800 19576
rect 0 19184 800 19304
rect 0 18776 800 18896
rect 0 18504 800 18624
rect 0 18232 800 18352
rect 0 17824 800 17944
rect 0 17552 800 17672
rect 0 17280 800 17400
rect 0 17008 800 17128
rect 0 16600 800 16720
rect 0 16328 800 16448
rect 0 16056 800 16176
rect 0 15648 800 15768
rect 0 15376 800 15496
rect 0 15104 800 15224
rect 0 14696 800 14816
rect 0 14424 800 14544
rect 0 14152 800 14272
rect 0 13880 800 14000
rect 0 13472 800 13592
rect 0 13200 800 13320
rect 0 12928 800 13048
rect 0 12520 800 12640
rect 0 12248 800 12368
rect 0 11976 800 12096
rect 0 11568 800 11688
rect 0 11296 800 11416
rect 0 11024 800 11144
rect 0 10752 800 10872
rect 0 10344 800 10464
rect 0 10072 800 10192
rect 0 9800 800 9920
rect 0 9392 800 9512
rect 0 9120 800 9240
rect 0 8848 800 8968
rect 0 8576 800 8696
rect 0 8168 800 8288
rect 0 7896 800 8016
rect 0 7624 800 7744
rect 0 7216 800 7336
rect 0 6944 800 7064
rect 0 6672 800 6792
rect 0 6264 800 6384
rect 0 5992 800 6112
rect 0 5720 800 5840
rect 0 5448 800 5568
rect 0 5040 800 5160
rect 0 4768 800 4888
rect 0 4496 800 4616
rect 0 4088 800 4208
rect 0 3816 800 3936
rect 0 3544 800 3664
rect 0 3136 800 3256
rect 0 2864 800 2984
rect 0 2592 800 2712
rect 0 2320 800 2440
rect 0 1912 800 2032
rect 0 1640 800 1760
rect 0 1368 800 1488
rect 0 960 800 1080
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
<< obsm3 >>
rect 880 119064 179200 119781
rect 800 118936 179200 119064
rect 880 118112 179200 118936
rect 800 117984 179200 118112
rect 880 116888 179200 117984
rect 800 116760 179200 116888
rect 880 115936 179200 116760
rect 800 115808 179200 115936
rect 880 114984 179200 115808
rect 800 114856 179200 114984
rect 880 113760 179200 114856
rect 800 113632 179200 113760
rect 880 112808 179200 113632
rect 800 112680 179200 112808
rect 880 111856 179200 112680
rect 800 111728 179200 111856
rect 880 110632 179200 111728
rect 800 110504 179200 110632
rect 880 109680 179200 110504
rect 800 109552 179200 109680
rect 880 108456 179200 109552
rect 800 108328 179200 108456
rect 880 107504 179200 108328
rect 800 107376 179200 107504
rect 880 106552 179200 107376
rect 800 106424 179200 106552
rect 880 105328 179200 106424
rect 800 105200 179200 105328
rect 880 104376 179200 105200
rect 800 104248 179200 104376
rect 880 103424 179200 104248
rect 800 103296 179200 103424
rect 880 102200 179200 103296
rect 800 102072 179200 102200
rect 880 101248 179200 102072
rect 800 101120 179200 101248
rect 880 100024 179200 101120
rect 800 99896 179200 100024
rect 880 99072 179200 99896
rect 800 98944 179200 99072
rect 880 98120 179200 98944
rect 800 97992 179200 98120
rect 880 96896 179200 97992
rect 800 96768 179200 96896
rect 880 95944 179200 96768
rect 800 95816 179200 95944
rect 880 94992 179200 95816
rect 800 94864 179200 94992
rect 880 93768 179200 94864
rect 800 93640 179200 93768
rect 880 92816 179200 93640
rect 800 92688 179200 92816
rect 880 91864 179200 92688
rect 800 91736 179200 91864
rect 880 90640 179200 91736
rect 800 90512 179200 90640
rect 880 89688 179200 90512
rect 800 89560 179200 89688
rect 880 88464 179200 89560
rect 800 88336 179200 88464
rect 880 87512 179200 88336
rect 800 87384 179200 87512
rect 880 86560 179200 87384
rect 800 86432 179200 86560
rect 880 85336 179200 86432
rect 800 85208 179200 85336
rect 880 84384 179200 85208
rect 800 84256 179200 84384
rect 880 83432 179200 84256
rect 800 83304 179200 83432
rect 880 82208 179200 83304
rect 800 82080 179200 82208
rect 880 81256 179200 82080
rect 800 81128 179200 81256
rect 880 80032 179200 81128
rect 800 79904 179200 80032
rect 880 79080 179200 79904
rect 800 78952 179200 79080
rect 880 78128 179200 78952
rect 800 78000 179200 78128
rect 880 76904 179200 78000
rect 800 76776 179200 76904
rect 880 75952 179200 76776
rect 800 75824 179200 75952
rect 880 75000 179200 75824
rect 800 74872 179200 75000
rect 880 73776 179200 74872
rect 800 73648 179200 73776
rect 880 72824 179200 73648
rect 800 72696 179200 72824
rect 880 71872 179200 72696
rect 800 71744 179200 71872
rect 880 70648 179200 71744
rect 800 70520 179200 70648
rect 880 69696 179200 70520
rect 800 69568 179200 69696
rect 880 68472 179200 69568
rect 800 68344 179200 68472
rect 880 67520 179200 68344
rect 800 67392 179200 67520
rect 880 66568 179200 67392
rect 800 66440 179200 66568
rect 880 65344 179200 66440
rect 800 65216 179200 65344
rect 880 64392 179200 65216
rect 800 64264 179200 64392
rect 880 63440 179200 64264
rect 800 63312 179200 63440
rect 880 62216 179200 63312
rect 800 62088 179200 62216
rect 880 61264 179200 62088
rect 800 61136 179200 61264
rect 880 60184 179200 61136
rect 880 60040 179120 60184
rect 800 59912 179120 60040
rect 880 59904 179120 59912
rect 880 59088 179200 59904
rect 800 58960 179200 59088
rect 880 58136 179200 58960
rect 800 58008 179200 58136
rect 880 56912 179200 58008
rect 800 56784 179200 56912
rect 880 55960 179200 56784
rect 800 55832 179200 55960
rect 880 55008 179200 55832
rect 800 54880 179200 55008
rect 880 53784 179200 54880
rect 800 53656 179200 53784
rect 880 52832 179200 53656
rect 800 52704 179200 52832
rect 880 51880 179200 52704
rect 800 51752 179200 51880
rect 880 50656 179200 51752
rect 800 50528 179200 50656
rect 880 49704 179200 50528
rect 800 49576 179200 49704
rect 880 48480 179200 49576
rect 800 48352 179200 48480
rect 880 47528 179200 48352
rect 800 47400 179200 47528
rect 880 46576 179200 47400
rect 800 46448 179200 46576
rect 880 45352 179200 46448
rect 800 45224 179200 45352
rect 880 44400 179200 45224
rect 800 44272 179200 44400
rect 880 43448 179200 44272
rect 800 43320 179200 43448
rect 880 42224 179200 43320
rect 800 42096 179200 42224
rect 880 41272 179200 42096
rect 800 41144 179200 41272
rect 880 40048 179200 41144
rect 800 39920 179200 40048
rect 880 39096 179200 39920
rect 800 38968 179200 39096
rect 880 38144 179200 38968
rect 800 38016 179200 38144
rect 880 36920 179200 38016
rect 800 36792 179200 36920
rect 880 35968 179200 36792
rect 800 35840 179200 35968
rect 880 35016 179200 35840
rect 800 34888 179200 35016
rect 880 33792 179200 34888
rect 800 33664 179200 33792
rect 880 32840 179200 33664
rect 800 32712 179200 32840
rect 880 31888 179200 32712
rect 800 31760 179200 31888
rect 880 30664 179200 31760
rect 800 30536 179200 30664
rect 880 29712 179200 30536
rect 800 29584 179200 29712
rect 880 28488 179200 29584
rect 800 28360 179200 28488
rect 880 27536 179200 28360
rect 800 27408 179200 27536
rect 880 26584 179200 27408
rect 800 26456 179200 26584
rect 880 25360 179200 26456
rect 800 25232 179200 25360
rect 880 24408 179200 25232
rect 800 24280 179200 24408
rect 880 23456 179200 24280
rect 800 23328 179200 23456
rect 880 22232 179200 23328
rect 800 22104 179200 22232
rect 880 21280 179200 22104
rect 800 21152 179200 21280
rect 880 20056 179200 21152
rect 800 19928 179200 20056
rect 880 19104 179200 19928
rect 800 18976 179200 19104
rect 880 18152 179200 18976
rect 800 18024 179200 18152
rect 880 16928 179200 18024
rect 800 16800 179200 16928
rect 880 15976 179200 16800
rect 800 15848 179200 15976
rect 880 15024 179200 15848
rect 800 14896 179200 15024
rect 880 13800 179200 14896
rect 800 13672 179200 13800
rect 880 12848 179200 13672
rect 800 12720 179200 12848
rect 880 11896 179200 12720
rect 800 11768 179200 11896
rect 880 10672 179200 11768
rect 800 10544 179200 10672
rect 880 9720 179200 10544
rect 800 9592 179200 9720
rect 880 8496 179200 9592
rect 800 8368 179200 8496
rect 880 7544 179200 8368
rect 800 7416 179200 7544
rect 880 6592 179200 7416
rect 800 6464 179200 6592
rect 880 5368 179200 6464
rect 800 5240 179200 5368
rect 880 4416 179200 5240
rect 800 4288 179200 4416
rect 880 3464 179200 4288
rect 800 3336 179200 3464
rect 880 2240 179200 3336
rect 800 2112 179200 2240
rect 880 1288 179200 2112
rect 800 1160 179200 1288
rect 880 171 179200 1160
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< obsm4 >>
rect 106227 15539 106293 16149
<< labels >>
rlabel metal2 s 662 119200 718 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 43166 119200 43222 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 47398 119200 47454 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 51630 119200 51686 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 55862 119200 55918 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 60186 119200 60242 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 64418 119200 64474 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 68650 119200 68706 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 72882 119200 72938 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 77206 119200 77262 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 81438 119200 81494 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4894 119200 4950 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 85670 119200 85726 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 89902 119200 89958 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 94226 119200 94282 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 98458 119200 98514 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 102690 119200 102746 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 106922 119200 106978 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 111154 119200 111210 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 115478 119200 115534 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 119710 119200 119766 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 123942 119200 123998 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9126 119200 9182 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 128174 119200 128230 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 132498 119200 132554 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 136730 119200 136786 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 140962 119200 141018 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 145194 119200 145250 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 149426 119200 149482 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 153750 119200 153806 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 157982 119200 158038 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13358 119200 13414 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17590 119200 17646 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 21914 119200 21970 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 26146 119200 26202 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 30378 119200 30434 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 34610 119200 34666 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 38934 119200 38990 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2042 119200 2098 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 44546 119200 44602 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 48778 119200 48834 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 53102 119200 53158 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 57334 119200 57390 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 61566 119200 61622 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 65798 119200 65854 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 70122 119200 70178 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 74354 119200 74410 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 78586 119200 78642 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 82818 119200 82874 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6274 119200 6330 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 87050 119200 87106 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 91374 119200 91430 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 95606 119200 95662 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 99838 119200 99894 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 104070 119200 104126 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 108394 119200 108450 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 112626 119200 112682 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 116858 119200 116914 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 121090 119200 121146 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 125414 119200 125470 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 10506 119200 10562 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 129646 119200 129702 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 133878 119200 133934 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 138110 119200 138166 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 142342 119200 142398 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 146666 119200 146722 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 150898 119200 150954 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 155130 119200 155186 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 159362 119200 159418 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 14830 119200 14886 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 19062 119200 19118 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 23294 119200 23350 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 27526 119200 27582 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 31850 119200 31906 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 36082 119200 36138 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 40314 119200 40370 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3422 119200 3478 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 46018 119200 46074 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 50250 119200 50306 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 54482 119200 54538 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 58714 119200 58770 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 63038 119200 63094 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 67270 119200 67326 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 71502 119200 71558 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 75734 119200 75790 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 79966 119200 80022 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 84290 119200 84346 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7746 119200 7802 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 88522 119200 88578 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 92754 119200 92810 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 96986 119200 97042 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 101310 119200 101366 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 105542 119200 105598 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 109774 119200 109830 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 114006 119200 114062 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 118238 119200 118294 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 122562 119200 122618 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 126794 119200 126850 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 11978 119200 12034 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 131026 119200 131082 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 135258 119200 135314 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 139582 119200 139638 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 143814 119200 143870 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 148046 119200 148102 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 152278 119200 152334 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 156602 119200 156658 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 160834 119200 160890 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16210 119200 16266 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20442 119200 20498 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 24674 119200 24730 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 28998 119200 29054 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 33230 119200 33286 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 37462 119200 37518 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 41694 119200 41750 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 177854 119200 177910 120000 6 irq[0]
port 115 nsew signal output
rlabel metal3 s 179200 59984 180000 60104 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 179234 119200 179290 120000 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 0 144 800 264 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 la_data_in[100]
port 119 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 la_data_in[101]
port 120 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 la_data_in[106]
port 125 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 la_data_in[108]
port 127 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 la_data_in[10]
port 129 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 0 105952 800 106072 6 la_data_in[113]
port 133 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 la_data_in[114]
port 134 nsew signal input
rlabel metal3 s 0 107856 800 107976 6 la_data_in[115]
port 135 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 la_data_in[116]
port 136 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 la_data_in[117]
port 137 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 la_data_in[11]
port 140 nsew signal input
rlabel metal3 s 0 112480 800 112600 6 la_data_in[120]
port 141 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 la_data_in[121]
port 142 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 la_data_in[122]
port 143 nsew signal input
rlabel metal3 s 0 115336 800 115456 6 la_data_in[123]
port 144 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 la_data_in[125]
port 146 nsew signal input
rlabel metal3 s 0 118192 800 118312 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 la_data_in[12]
port 149 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 la_data_in[18]
port 155 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 la_data_in[19]
port 156 nsew signal input
rlabel metal3 s 0 960 800 1080 6 la_data_in[1]
port 157 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 la_data_in[21]
port 159 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 la_data_in[28]
port 166 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 la_data_in[29]
port 167 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 la_data_in[2]
port 168 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 la_data_in[30]
port 169 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 la_data_in[31]
port 170 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 la_data_in[32]
port 171 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 la_data_in[33]
port 172 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 la_data_in[35]
port 174 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 la_data_in[36]
port 175 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 la_data_in[38]
port 177 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 la_data_in[3]
port 179 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 la_data_in[40]
port 180 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 la_data_in[43]
port 183 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 la_data_in[46]
port 186 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 la_data_in[47]
port 187 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 la_data_in[48]
port 188 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 la_data_in[49]
port 189 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 la_data_in[50]
port 191 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 la_data_in[51]
port 192 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 la_data_in[53]
port 194 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 la_data_in[54]
port 195 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 la_data_in[55]
port 196 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 la_data_in[56]
port 197 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 la_data_in[57]
port 198 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_data_in[58]
port 199 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_data_in[5]
port 201 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 la_data_in[60]
port 202 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 la_data_in[64]
port 206 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 la_data_in[66]
port 208 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 la_data_in[71]
port 214 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 la_data_in[72]
port 215 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 la_data_in[73]
port 216 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 la_data_in[74]
port 217 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 la_data_in[75]
port 218 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 la_data_in[7]
port 223 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 la_data_in[82]
port 226 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 la_data_in[84]
port 228 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 0 80656 800 80776 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 la_data_in[88]
port 232 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 la_data_in[89]
port 233 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 la_data_in[8]
port 234 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 la_data_in[90]
port 235 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 la_data_in[92]
port 237 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 la_data_in[93]
port 238 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 0 90992 800 91112 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 la_data_in[99]
port 244 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 416 800 536 6 la_data_out[0]
port 246 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 0 95072 800 95192 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 0 96976 800 97096 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 la_data_out[105]
port 252 nsew signal output
rlabel metal3 s 0 99696 800 99816 6 la_data_out[106]
port 253 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 la_data_out[108]
port 255 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 la_data_out[109]
port 256 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 la_data_out[10]
port 257 nsew signal output
rlabel metal3 s 0 103504 800 103624 6 la_data_out[110]
port 258 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 la_data_out[111]
port 259 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 106224 800 106344 6 la_data_out[113]
port 261 nsew signal output
rlabel metal3 s 0 107176 800 107296 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 110032 800 110152 6 la_data_out[117]
port 265 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 111936 800 112056 6 la_data_out[119]
port 267 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 la_data_out[120]
port 269 nsew signal output
rlabel metal3 s 0 113840 800 113960 6 la_data_out[121]
port 270 nsew signal output
rlabel metal3 s 0 114656 800 114776 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 116560 800 116680 6 la_data_out[124]
port 273 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 la_data_out[125]
port 274 nsew signal output
rlabel metal3 s 0 118464 800 118584 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 119416 800 119536 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 la_data_out[15]
port 280 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 la_data_out[16]
port 281 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 la_data_out[19]
port 284 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 la_data_out[21]
port 287 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 la_data_out[23]
port 289 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 la_data_out[24]
port 290 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 la_data_out[27]
port 293 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 la_data_out[2]
port 296 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 la_data_out[31]
port 298 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 la_data_out[32]
port 299 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 la_data_out[33]
port 300 nsew signal output
rlabel metal3 s 0 32240 800 32360 6 la_data_out[34]
port 301 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 la_data_out[37]
port 304 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 la_data_out[39]
port 306 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 la_data_out[40]
port 308 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 la_data_out[41]
port 309 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 la_data_out[42]
port 310 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 la_data_out[43]
port 311 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 la_data_out[45]
port 313 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 la_data_out[46]
port 314 nsew signal output
rlabel metal3 s 0 44480 800 44600 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 la_data_out[48]
port 316 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 la_data_out[50]
port 319 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 49104 800 49224 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 la_data_out[56]
port 325 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 la_data_out[57]
port 326 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 la_data_out[59]
port 328 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 la_data_out[5]
port 329 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 la_data_out[60]
port 330 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 la_data_out[65]
port 335 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 la_data_out[66]
port 336 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 la_data_out[67]
port 337 nsew signal output
rlabel metal3 s 0 64064 800 64184 6 la_data_out[68]
port 338 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 la_data_out[69]
port 339 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 la_data_out[6]
port 340 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 0 66920 800 67040 6 la_data_out[71]
port 342 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 la_data_out[72]
port 343 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 la_data_out[73]
port 344 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 la_data_out[75]
port 346 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 0 72496 800 72616 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 la_data_out[78]
port 349 nsew signal output
rlabel metal3 s 0 74400 800 74520 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 la_data_out[80]
port 352 nsew signal output
rlabel metal3 s 0 76304 800 76424 6 la_data_out[81]
port 353 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 la_data_out[82]
port 354 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 79160 800 79280 6 la_data_out[84]
port 356 nsew signal output
rlabel metal3 s 0 80112 800 80232 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 la_data_out[86]
port 358 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 la_data_out[87]
port 359 nsew signal output
rlabel metal3 s 0 82832 800 82952 6 la_data_out[88]
port 360 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 la_data_out[89]
port 361 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 la_data_out[8]
port 362 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 la_data_out[90]
port 363 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 la_data_out[91]
port 364 nsew signal output
rlabel metal3 s 0 86640 800 86760 6 la_data_out[92]
port 365 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 la_data_out[93]
port 366 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 la_data_out[94]
port 367 nsew signal output
rlabel metal3 s 0 89360 800 89480 6 la_data_out[95]
port 368 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 91264 800 91384 6 la_data_out[97]
port 370 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 la_data_out[98]
port 371 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 la_data_out[99]
port 372 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 la_data_out[9]
port 373 nsew signal output
rlabel metal3 s 0 688 800 808 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 0 95344 800 95464 6 la_oenb[101]
port 376 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 la_oenb[102]
port 377 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 la_oenb[104]
port 379 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 la_oenb[105]
port 380 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 la_oenb[107]
port 382 nsew signal input
rlabel metal3 s 0 101872 800 101992 6 la_oenb[108]
port 383 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 la_oenb[109]
port 384 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 0 103776 800 103896 6 la_oenb[110]
port 386 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 la_oenb[113]
port 389 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 la_oenb[114]
port 390 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 la_oenb[115]
port 391 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 0 110304 800 110424 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 la_oenb[11]
port 396 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 la_oenb[120]
port 397 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 0 116016 800 116136 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 la_oenb[125]
port 402 nsew signal input
rlabel metal3 s 0 118736 800 118856 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 la_oenb[14]
port 407 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 la_oenb[15]
port 408 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 la_oenb[17]
port 410 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 la_oenb[18]
port 411 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_oenb[21]
port 415 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 la_oenb[23]
port 417 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_oenb[24]
port 418 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 la_oenb[25]
port 419 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 la_oenb[27]
port 421 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 la_oenb[28]
port 422 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 la_oenb[30]
port 425 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 la_oenb[31]
port 426 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 la_oenb[32]
port 427 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 la_oenb[36]
port 431 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 la_oenb[39]
port 434 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 la_oenb[40]
port 436 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 la_oenb[41]
port 437 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 la_oenb[44]
port 440 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_oenb[45]
port 441 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 la_oenb[46]
port 442 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 la_oenb[4]
port 446 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 la_oenb[50]
port 447 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 51280 800 51400 6 la_oenb[54]
port 451 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 la_oenb[57]
port 454 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 la_oenb[59]
port 456 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 la_oenb[5]
port 457 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 la_oenb[60]
port 458 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 la_oenb[61]
port 459 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 la_oenb[62]
port 460 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 la_oenb[63]
port 461 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 la_oenb[64]
port 462 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 la_oenb[65]
port 463 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 63520 800 63640 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 65424 800 65544 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 la_oenb[73]
port 472 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 la_oenb[74]
port 473 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 la_oenb[75]
port 474 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 la_oenb[82]
port 482 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 la_oenb[84]
port 484 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 la_oenb[87]
port 487 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 la_oenb[8]
port 490 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 la_oenb[91]
port 492 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 la_oenb[93]
port 494 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 la_oenb[95]
port 496 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 la_oenb[96]
port 497 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 0 93440 800 93560 6 la_oenb[99]
port 500 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 162214 119200 162270 120000 6 phase_in[0]
port 502 nsew signal input
rlabel metal2 s 176382 119200 176438 120000 6 phase_in[10]
port 503 nsew signal input
rlabel metal2 s 163686 119200 163742 120000 6 phase_in[1]
port 504 nsew signal input
rlabel metal2 s 165066 119200 165122 120000 6 phase_in[2]
port 505 nsew signal input
rlabel metal2 s 166446 119200 166502 120000 6 phase_in[3]
port 506 nsew signal input
rlabel metal2 s 167918 119200 167974 120000 6 phase_in[4]
port 507 nsew signal input
rlabel metal2 s 169298 119200 169354 120000 6 phase_in[5]
port 508 nsew signal input
rlabel metal2 s 170770 119200 170826 120000 6 phase_in[6]
port 509 nsew signal input
rlabel metal2 s 172150 119200 172206 120000 6 phase_in[7]
port 510 nsew signal input
rlabel metal2 s 173530 119200 173586 120000 6 phase_in[8]
port 511 nsew signal input
rlabel metal2 s 175002 119200 175058 120000 6 phase_in[9]
port 512 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_clk_i
port 513 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wb_rst_i
port 514 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_ack_o
port 515 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 wbs_adr_i[0]
port 516 nsew signal input
rlabel metal2 s 68742 0 68798 800 6 wbs_adr_i[10]
port 517 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 wbs_adr_i[11]
port 518 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 wbs_adr_i[12]
port 519 nsew signal input
rlabel metal2 s 84014 0 84070 800 6 wbs_adr_i[13]
port 520 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_adr_i[14]
port 521 nsew signal input
rlabel metal2 s 94226 0 94282 800 6 wbs_adr_i[15]
port 522 nsew signal input
rlabel metal2 s 99286 0 99342 800 6 wbs_adr_i[16]
port 523 nsew signal input
rlabel metal2 s 104438 0 104494 800 6 wbs_adr_i[17]
port 524 nsew signal input
rlabel metal2 s 109498 0 109554 800 6 wbs_adr_i[18]
port 525 nsew signal input
rlabel metal2 s 114558 0 114614 800 6 wbs_adr_i[19]
port 526 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_adr_i[1]
port 527 nsew signal input
rlabel metal2 s 119710 0 119766 800 6 wbs_adr_i[20]
port 528 nsew signal input
rlabel metal2 s 124770 0 124826 800 6 wbs_adr_i[21]
port 529 nsew signal input
rlabel metal2 s 129922 0 129978 800 6 wbs_adr_i[22]
port 530 nsew signal input
rlabel metal2 s 134982 0 135038 800 6 wbs_adr_i[23]
port 531 nsew signal input
rlabel metal2 s 140042 0 140098 800 6 wbs_adr_i[24]
port 532 nsew signal input
rlabel metal2 s 145194 0 145250 800 6 wbs_adr_i[25]
port 533 nsew signal input
rlabel metal2 s 150254 0 150310 800 6 wbs_adr_i[26]
port 534 nsew signal input
rlabel metal2 s 155406 0 155462 800 6 wbs_adr_i[27]
port 535 nsew signal input
rlabel metal2 s 160466 0 160522 800 6 wbs_adr_i[28]
port 536 nsew signal input
rlabel metal2 s 165526 0 165582 800 6 wbs_adr_i[29]
port 537 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 wbs_adr_i[2]
port 538 nsew signal input
rlabel metal2 s 170678 0 170734 800 6 wbs_adr_i[30]
port 539 nsew signal input
rlabel metal2 s 175738 0 175794 800 6 wbs_adr_i[31]
port 540 nsew signal input
rlabel metal2 s 31390 0 31446 800 6 wbs_adr_i[3]
port 541 nsew signal input
rlabel metal2 s 38198 0 38254 800 6 wbs_adr_i[4]
port 542 nsew signal input
rlabel metal2 s 43258 0 43314 800 6 wbs_adr_i[5]
port 543 nsew signal input
rlabel metal2 s 48318 0 48374 800 6 wbs_adr_i[6]
port 544 nsew signal input
rlabel metal2 s 53470 0 53526 800 6 wbs_adr_i[7]
port 545 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 wbs_adr_i[8]
port 546 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 wbs_adr_i[9]
port 547 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 wbs_cyc_i
port 548 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_dat_i[0]
port 549 nsew signal input
rlabel metal2 s 70398 0 70454 800 6 wbs_dat_i[10]
port 550 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 wbs_dat_i[11]
port 551 nsew signal input
rlabel metal2 s 80610 0 80666 800 6 wbs_dat_i[12]
port 552 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 wbs_dat_i[13]
port 553 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_i[14]
port 554 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 wbs_dat_i[15]
port 555 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 wbs_dat_i[16]
port 556 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 wbs_dat_i[17]
port 557 nsew signal input
rlabel metal2 s 111246 0 111302 800 6 wbs_dat_i[18]
port 558 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 wbs_dat_i[19]
port 559 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[1]
port 560 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 wbs_dat_i[20]
port 561 nsew signal input
rlabel metal2 s 126518 0 126574 800 6 wbs_dat_i[21]
port 562 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 wbs_dat_i[22]
port 563 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 wbs_dat_i[23]
port 564 nsew signal input
rlabel metal2 s 141790 0 141846 800 6 wbs_dat_i[24]
port 565 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 wbs_dat_i[25]
port 566 nsew signal input
rlabel metal2 s 152002 0 152058 800 6 wbs_dat_i[26]
port 567 nsew signal input
rlabel metal2 s 157062 0 157118 800 6 wbs_dat_i[27]
port 568 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 wbs_dat_i[28]
port 569 nsew signal input
rlabel metal2 s 167274 0 167330 800 6 wbs_dat_i[29]
port 570 nsew signal input
rlabel metal2 s 26238 0 26294 800 6 wbs_dat_i[2]
port 571 nsew signal input
rlabel metal2 s 172334 0 172390 800 6 wbs_dat_i[30]
port 572 nsew signal input
rlabel metal2 s 177486 0 177542 800 6 wbs_dat_i[31]
port 573 nsew signal input
rlabel metal2 s 33046 0 33102 800 6 wbs_dat_i[3]
port 574 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 wbs_dat_i[4]
port 575 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 wbs_dat_i[5]
port 576 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 wbs_dat_i[6]
port 577 nsew signal input
rlabel metal2 s 55126 0 55182 800 6 wbs_dat_i[7]
port 578 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 wbs_dat_i[8]
port 579 nsew signal input
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_i[9]
port 580 nsew signal input
rlabel metal2 s 14370 0 14426 800 6 wbs_dat_o[0]
port 581 nsew signal output
rlabel metal2 s 72146 0 72202 800 6 wbs_dat_o[10]
port 582 nsew signal output
rlabel metal2 s 77206 0 77262 800 6 wbs_dat_o[11]
port 583 nsew signal output
rlabel metal2 s 82358 0 82414 800 6 wbs_dat_o[12]
port 584 nsew signal output
rlabel metal2 s 87418 0 87474 800 6 wbs_dat_o[13]
port 585 nsew signal output
rlabel metal2 s 92478 0 92534 800 6 wbs_dat_o[14]
port 586 nsew signal output
rlabel metal2 s 97630 0 97686 800 6 wbs_dat_o[15]
port 587 nsew signal output
rlabel metal2 s 102690 0 102746 800 6 wbs_dat_o[16]
port 588 nsew signal output
rlabel metal2 s 107842 0 107898 800 6 wbs_dat_o[17]
port 589 nsew signal output
rlabel metal2 s 112902 0 112958 800 6 wbs_dat_o[18]
port 590 nsew signal output
rlabel metal2 s 117962 0 118018 800 6 wbs_dat_o[19]
port 591 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 wbs_dat_o[1]
port 592 nsew signal output
rlabel metal2 s 123114 0 123170 800 6 wbs_dat_o[20]
port 593 nsew signal output
rlabel metal2 s 128174 0 128230 800 6 wbs_dat_o[21]
port 594 nsew signal output
rlabel metal2 s 133326 0 133382 800 6 wbs_dat_o[22]
port 595 nsew signal output
rlabel metal2 s 138386 0 138442 800 6 wbs_dat_o[23]
port 596 nsew signal output
rlabel metal2 s 143446 0 143502 800 6 wbs_dat_o[24]
port 597 nsew signal output
rlabel metal2 s 148598 0 148654 800 6 wbs_dat_o[25]
port 598 nsew signal output
rlabel metal2 s 153658 0 153714 800 6 wbs_dat_o[26]
port 599 nsew signal output
rlabel metal2 s 158718 0 158774 800 6 wbs_dat_o[27]
port 600 nsew signal output
rlabel metal2 s 163870 0 163926 800 6 wbs_dat_o[28]
port 601 nsew signal output
rlabel metal2 s 168930 0 168986 800 6 wbs_dat_o[29]
port 602 nsew signal output
rlabel metal2 s 27986 0 28042 800 6 wbs_dat_o[2]
port 603 nsew signal output
rlabel metal2 s 174082 0 174138 800 6 wbs_dat_o[30]
port 604 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 wbs_dat_o[31]
port 605 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 wbs_dat_o[3]
port 606 nsew signal output
rlabel metal2 s 41602 0 41658 800 6 wbs_dat_o[4]
port 607 nsew signal output
rlabel metal2 s 46662 0 46718 800 6 wbs_dat_o[5]
port 608 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 wbs_dat_o[6]
port 609 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[7]
port 610 nsew signal output
rlabel metal2 s 61934 0 61990 800 6 wbs_dat_o[8]
port 611 nsew signal output
rlabel metal2 s 67086 0 67142 800 6 wbs_dat_o[9]
port 612 nsew signal output
rlabel metal2 s 16118 0 16174 800 6 wbs_sel_i[0]
port 613 nsew signal input
rlabel metal2 s 22926 0 22982 800 6 wbs_sel_i[1]
port 614 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 wbs_sel_i[2]
port 615 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 wbs_sel_i[3]
port 616 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_stb_i
port 617 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_we_i
port 618 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 619 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 620 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 621 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 622 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 624 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 625 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 626 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 627 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 628 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 629 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 630 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 634 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 635 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 636 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 637 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 642 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 643 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 644 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 645 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 646 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 649 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 650 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 651 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 652 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 653 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 654 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 655 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 656 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 657 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 658 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 659 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 660 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 661 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 662 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 663 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 664 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 665 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 666 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 17864168
string GDS_START 1001754
<< end >>

