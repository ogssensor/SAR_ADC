VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vco_adc_wrapper
  CLASS BLOCK ;
  FOREIGN vco_adc_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 900.000 BY 700.000 ;
  PIN adc0_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 2.760 900.000 3.360 ;
    END
  END adc0_dat_i[0]
  PIN adc0_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 214.240 900.000 214.840 ;
    END
  END adc0_dat_i[10]
  PIN adc0_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 233.280 900.000 233.880 ;
    END
  END adc0_dat_i[11]
  PIN adc0_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 253.000 900.000 253.600 ;
    END
  END adc0_dat_i[12]
  PIN adc0_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 272.040 900.000 272.640 ;
    END
  END adc0_dat_i[13]
  PIN adc0_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 291.080 900.000 291.680 ;
    END
  END adc0_dat_i[14]
  PIN adc0_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 310.800 900.000 311.400 ;
    END
  END adc0_dat_i[15]
  PIN adc0_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 329.840 900.000 330.440 ;
    END
  END adc0_dat_i[16]
  PIN adc0_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 348.880 900.000 349.480 ;
    END
  END adc0_dat_i[17]
  PIN adc0_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 368.600 900.000 369.200 ;
    END
  END adc0_dat_i[18]
  PIN adc0_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 387.640 900.000 388.240 ;
    END
  END adc0_dat_i[19]
  PIN adc0_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 27.920 900.000 28.520 ;
    END
  END adc0_dat_i[1]
  PIN adc0_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 406.680 900.000 407.280 ;
    END
  END adc0_dat_i[20]
  PIN adc0_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 426.400 900.000 427.000 ;
    END
  END adc0_dat_i[21]
  PIN adc0_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 445.440 900.000 446.040 ;
    END
  END adc0_dat_i[22]
  PIN adc0_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 464.480 900.000 465.080 ;
    END
  END adc0_dat_i[23]
  PIN adc0_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 484.200 900.000 484.800 ;
    END
  END adc0_dat_i[24]
  PIN adc0_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 503.240 900.000 503.840 ;
    END
  END adc0_dat_i[25]
  PIN adc0_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 522.280 900.000 522.880 ;
    END
  END adc0_dat_i[26]
  PIN adc0_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 541.320 900.000 541.920 ;
    END
  END adc0_dat_i[27]
  PIN adc0_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 561.040 900.000 561.640 ;
    END
  END adc0_dat_i[28]
  PIN adc0_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 580.080 900.000 580.680 ;
    END
  END adc0_dat_i[29]
  PIN adc0_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 53.760 900.000 54.360 ;
    END
  END adc0_dat_i[2]
  PIN adc0_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 599.120 900.000 599.720 ;
    END
  END adc0_dat_i[30]
  PIN adc0_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 618.840 900.000 619.440 ;
    END
  END adc0_dat_i[31]
  PIN adc0_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 79.600 900.000 80.200 ;
    END
  END adc0_dat_i[3]
  PIN adc0_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 98.640 900.000 99.240 ;
    END
  END adc0_dat_i[4]
  PIN adc0_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 117.680 900.000 118.280 ;
    END
  END adc0_dat_i[5]
  PIN adc0_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 137.400 900.000 138.000 ;
    END
  END adc0_dat_i[6]
  PIN adc0_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 156.440 900.000 157.040 ;
    END
  END adc0_dat_i[7]
  PIN adc0_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 175.480 900.000 176.080 ;
    END
  END adc0_dat_i[8]
  PIN adc0_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 195.200 900.000 195.800 ;
    END
  END adc0_dat_i[9]
  PIN adc1_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 8.880 900.000 9.480 ;
    END
  END adc1_dat_i[0]
  PIN adc1_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 220.360 900.000 220.960 ;
    END
  END adc1_dat_i[10]
  PIN adc1_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 240.080 900.000 240.680 ;
    END
  END adc1_dat_i[11]
  PIN adc1_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 259.120 900.000 259.720 ;
    END
  END adc1_dat_i[12]
  PIN adc1_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 278.160 900.000 278.760 ;
    END
  END adc1_dat_i[13]
  PIN adc1_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 297.880 900.000 298.480 ;
    END
  END adc1_dat_i[14]
  PIN adc1_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 316.920 900.000 317.520 ;
    END
  END adc1_dat_i[15]
  PIN adc1_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 335.960 900.000 336.560 ;
    END
  END adc1_dat_i[16]
  PIN adc1_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 355.680 900.000 356.280 ;
    END
  END adc1_dat_i[17]
  PIN adc1_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 374.720 900.000 375.320 ;
    END
  END adc1_dat_i[18]
  PIN adc1_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 393.760 900.000 394.360 ;
    END
  END adc1_dat_i[19]
  PIN adc1_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 34.720 900.000 35.320 ;
    END
  END adc1_dat_i[1]
  PIN adc1_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 413.480 900.000 414.080 ;
    END
  END adc1_dat_i[20]
  PIN adc1_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 432.520 900.000 433.120 ;
    END
  END adc1_dat_i[21]
  PIN adc1_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 451.560 900.000 452.160 ;
    END
  END adc1_dat_i[22]
  PIN adc1_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 471.280 900.000 471.880 ;
    END
  END adc1_dat_i[23]
  PIN adc1_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 490.320 900.000 490.920 ;
    END
  END adc1_dat_i[24]
  PIN adc1_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 509.360 900.000 509.960 ;
    END
  END adc1_dat_i[25]
  PIN adc1_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 529.080 900.000 529.680 ;
    END
  END adc1_dat_i[26]
  PIN adc1_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 548.120 900.000 548.720 ;
    END
  END adc1_dat_i[27]
  PIN adc1_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 567.160 900.000 567.760 ;
    END
  END adc1_dat_i[28]
  PIN adc1_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 586.880 900.000 587.480 ;
    END
  END adc1_dat_i[29]
  PIN adc1_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 59.880 900.000 60.480 ;
    END
  END adc1_dat_i[2]
  PIN adc1_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 605.920 900.000 606.520 ;
    END
  END adc1_dat_i[30]
  PIN adc1_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 624.960 900.000 625.560 ;
    END
  END adc1_dat_i[31]
  PIN adc1_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 85.720 900.000 86.320 ;
    END
  END adc1_dat_i[3]
  PIN adc1_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 105.440 900.000 106.040 ;
    END
  END adc1_dat_i[4]
  PIN adc1_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 124.480 900.000 125.080 ;
    END
  END adc1_dat_i[5]
  PIN adc1_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 143.520 900.000 144.120 ;
    END
  END adc1_dat_i[6]
  PIN adc1_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 163.240 900.000 163.840 ;
    END
  END adc1_dat_i[7]
  PIN adc1_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 182.280 900.000 182.880 ;
    END
  END adc1_dat_i[8]
  PIN adc1_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 201.320 900.000 201.920 ;
    END
  END adc1_dat_i[9]
  PIN adc2_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 15.000 900.000 15.600 ;
    END
  END adc2_dat_i[0]
  PIN adc2_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 227.160 900.000 227.760 ;
    END
  END adc2_dat_i[10]
  PIN adc2_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 246.200 900.000 246.800 ;
    END
  END adc2_dat_i[11]
  PIN adc2_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 265.920 900.000 266.520 ;
    END
  END adc2_dat_i[12]
  PIN adc2_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 284.960 900.000 285.560 ;
    END
  END adc2_dat_i[13]
  PIN adc2_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 304.000 900.000 304.600 ;
    END
  END adc2_dat_i[14]
  PIN adc2_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 323.720 900.000 324.320 ;
    END
  END adc2_dat_i[15]
  PIN adc2_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 342.760 900.000 343.360 ;
    END
  END adc2_dat_i[16]
  PIN adc2_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 361.800 900.000 362.400 ;
    END
  END adc2_dat_i[17]
  PIN adc2_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 380.840 900.000 381.440 ;
    END
  END adc2_dat_i[18]
  PIN adc2_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 400.560 900.000 401.160 ;
    END
  END adc2_dat_i[19]
  PIN adc2_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 40.840 900.000 41.440 ;
    END
  END adc2_dat_i[1]
  PIN adc2_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 419.600 900.000 420.200 ;
    END
  END adc2_dat_i[20]
  PIN adc2_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 438.640 900.000 439.240 ;
    END
  END adc2_dat_i[21]
  PIN adc2_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 458.360 900.000 458.960 ;
    END
  END adc2_dat_i[22]
  PIN adc2_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 477.400 900.000 478.000 ;
    END
  END adc2_dat_i[23]
  PIN adc2_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 496.440 900.000 497.040 ;
    END
  END adc2_dat_i[24]
  PIN adc2_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 516.160 900.000 516.760 ;
    END
  END adc2_dat_i[25]
  PIN adc2_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 535.200 900.000 535.800 ;
    END
  END adc2_dat_i[26]
  PIN adc2_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 554.240 900.000 554.840 ;
    END
  END adc2_dat_i[27]
  PIN adc2_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 573.960 900.000 574.560 ;
    END
  END adc2_dat_i[28]
  PIN adc2_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 593.000 900.000 593.600 ;
    END
  END adc2_dat_i[29]
  PIN adc2_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 66.680 900.000 67.280 ;
    END
  END adc2_dat_i[2]
  PIN adc2_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 612.040 900.000 612.640 ;
    END
  END adc2_dat_i[30]
  PIN adc2_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 631.760 900.000 632.360 ;
    END
  END adc2_dat_i[31]
  PIN adc2_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 92.520 900.000 93.120 ;
    END
  END adc2_dat_i[3]
  PIN adc2_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 111.560 900.000 112.160 ;
    END
  END adc2_dat_i[4]
  PIN adc2_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 130.600 900.000 131.200 ;
    END
  END adc2_dat_i[5]
  PIN adc2_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 150.320 900.000 150.920 ;
    END
  END adc2_dat_i[6]
  PIN adc2_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 169.360 900.000 169.960 ;
    END
  END adc2_dat_i[7]
  PIN adc2_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 188.400 900.000 189.000 ;
    END
  END adc2_dat_i[8]
  PIN adc2_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 208.120 900.000 208.720 ;
    END
  END adc2_dat_i[9]
  PIN adc_dvalid_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 21.800 900.000 22.400 ;
    END
  END adc_dvalid_i[0]
  PIN adc_dvalid_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 47.640 900.000 48.240 ;
    END
  END adc_dvalid_i[1]
  PIN adc_dvalid_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 72.800 900.000 73.400 ;
    END
  END adc_dvalid_i[2]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 696.000 5.430 700.000 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 696.000 224.850 700.000 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 696.000 246.930 700.000 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.270 696.000 268.550 700.000 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 696.000 290.630 700.000 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 696.000 312.710 700.000 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.050 696.000 334.330 700.000 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 696.000 356.410 700.000 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 378.210 696.000 378.490 700.000 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 400.290 696.000 400.570 700.000 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 696.000 422.190 700.000 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 696.000 27.050 700.000 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.990 696.000 444.270 700.000 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 696.000 466.350 700.000 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 696.000 488.430 700.000 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.770 696.000 510.050 700.000 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 696.000 532.130 700.000 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.930 696.000 554.210 700.000 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.010 696.000 576.290 700.000 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.630 696.000 597.910 700.000 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.710 696.000 619.990 700.000 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 641.790 696.000 642.070 700.000 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 696.000 49.130 700.000 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 663.410 696.000 663.690 700.000 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 685.490 696.000 685.770 700.000 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 707.570 696.000 707.850 700.000 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.650 696.000 729.930 700.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 696.000 751.550 700.000 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 773.350 696.000 773.630 700.000 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 795.430 696.000 795.710 700.000 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 817.510 696.000 817.790 700.000 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 696.000 71.210 700.000 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 696.000 92.830 700.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 696.000 114.910 700.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.710 696.000 136.990 700.000 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.790 696.000 159.070 700.000 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 696.000 180.690 700.000 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.490 696.000 202.770 700.000 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 15.730 696.000 16.010 700.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.610 696.000 235.890 700.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.230 696.000 257.510 700.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.310 696.000 279.590 700.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 696.000 301.670 700.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.470 696.000 323.750 700.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.090 696.000 345.370 700.000 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 696.000 367.450 700.000 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.250 696.000 389.530 700.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.330 696.000 411.610 700.000 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 696.000 433.230 700.000 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 696.000 38.090 700.000 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 455.030 696.000 455.310 700.000 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 477.110 696.000 477.390 700.000 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 696.000 499.010 700.000 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.810 696.000 521.090 700.000 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 696.000 543.170 700.000 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 696.000 565.250 700.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.590 696.000 586.870 700.000 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.670 696.000 608.950 700.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 630.750 696.000 631.030 700.000 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 696.000 653.110 700.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.890 696.000 60.170 700.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.450 696.000 674.730 700.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.530 696.000 696.810 700.000 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 718.610 696.000 718.890 700.000 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 740.690 696.000 740.970 700.000 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.310 696.000 762.590 700.000 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 784.390 696.000 784.670 700.000 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.470 696.000 806.750 700.000 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 828.090 696.000 828.370 700.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.970 696.000 82.250 700.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.590 696.000 103.870 700.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 696.000 125.950 700.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 696.000 148.030 700.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.370 696.000 169.650 700.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 696.000 191.730 700.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 213.530 696.000 213.810 700.000 ;
    END
  END io_out[9]
  PIN mem1_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END mem1_data_i[0]
  PIN mem1_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 323.720 4.000 324.320 ;
    END
  END mem1_data_i[10]
  PIN mem1_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END mem1_data_i[11]
  PIN mem1_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.720 4.000 358.320 ;
    END
  END mem1_data_i[12]
  PIN mem1_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END mem1_data_i[13]
  PIN mem1_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 392.400 4.000 393.000 ;
    END
  END mem1_data_i[14]
  PIN mem1_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 409.400 4.000 410.000 ;
    END
  END mem1_data_i[15]
  PIN mem1_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.080 4.000 427.680 ;
    END
  END mem1_data_i[16]
  PIN mem1_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END mem1_data_i[17]
  PIN mem1_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.080 4.000 461.680 ;
    END
  END mem1_data_i[18]
  PIN mem1_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.760 4.000 479.360 ;
    END
  END mem1_data_i[19]
  PIN mem1_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 65.320 4.000 65.920 ;
    END
  END mem1_data_i[1]
  PIN mem1_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.760 4.000 496.360 ;
    END
  END mem1_data_i[20]
  PIN mem1_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 512.760 4.000 513.360 ;
    END
  END mem1_data_i[21]
  PIN mem1_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 529.760 4.000 530.360 ;
    END
  END mem1_data_i[22]
  PIN mem1_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END mem1_data_i[23]
  PIN mem1_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END mem1_data_i[24]
  PIN mem1_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END mem1_data_i[25]
  PIN mem1_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 599.120 4.000 599.720 ;
    END
  END mem1_data_i[26]
  PIN mem1_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END mem1_data_i[27]
  PIN mem1_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 633.120 4.000 633.720 ;
    END
  END mem1_data_i[28]
  PIN mem1_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 650.800 4.000 651.400 ;
    END
  END mem1_data_i[29]
  PIN mem1_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END mem1_data_i[2]
  PIN mem1_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 667.800 4.000 668.400 ;
    END
  END mem1_data_i[30]
  PIN mem1_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 684.800 4.000 685.400 ;
    END
  END mem1_data_i[31]
  PIN mem1_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 134.000 4.000 134.600 ;
    END
  END mem1_data_i[3]
  PIN mem1_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END mem1_data_i[4]
  PIN mem1_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END mem1_data_i[5]
  PIN mem1_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 220.360 4.000 220.960 ;
    END
  END mem1_data_i[6]
  PIN mem1_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END mem1_data_i[7]
  PIN mem1_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 277.480 4.000 278.080 ;
    END
  END mem1_data_i[8]
  PIN mem1_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END mem1_data_i[9]
  PIN mem_data_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 31.320 4.000 31.920 ;
    END
  END mem_data_i[0]
  PIN mem_data_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 329.160 4.000 329.760 ;
    END
  END mem_data_i[10]
  PIN mem_data_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END mem_data_i[11]
  PIN mem_data_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END mem_data_i[12]
  PIN mem_data_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END mem_data_i[13]
  PIN mem_data_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END mem_data_i[14]
  PIN mem_data_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END mem_data_i[15]
  PIN mem_data_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 432.520 4.000 433.120 ;
    END
  END mem_data_i[16]
  PIN mem_data_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END mem_data_i[17]
  PIN mem_data_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.200 4.000 467.800 ;
    END
  END mem_data_i[18]
  PIN mem_data_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.200 4.000 484.800 ;
    END
  END mem_data_i[19]
  PIN mem_data_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END mem_data_i[1]
  PIN mem_data_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END mem_data_i[20]
  PIN mem_data_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END mem_data_i[21]
  PIN mem_data_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 535.880 4.000 536.480 ;
    END
  END mem_data_i[22]
  PIN mem_data_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END mem_data_i[23]
  PIN mem_data_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 570.560 4.000 571.160 ;
    END
  END mem_data_i[24]
  PIN mem_data_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 587.560 4.000 588.160 ;
    END
  END mem_data_i[25]
  PIN mem_data_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 604.560 4.000 605.160 ;
    END
  END mem_data_i[26]
  PIN mem_data_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 621.560 4.000 622.160 ;
    END
  END mem_data_i[27]
  PIN mem_data_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 639.240 4.000 639.840 ;
    END
  END mem_data_i[28]
  PIN mem_data_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 656.240 4.000 656.840 ;
    END
  END mem_data_i[29]
  PIN mem_data_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 111.560 4.000 112.160 ;
    END
  END mem_data_i[2]
  PIN mem_data_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.240 4.000 673.840 ;
    END
  END mem_data_i[30]
  PIN mem_data_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END mem_data_i[31]
  PIN mem_data_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 140.120 4.000 140.720 ;
    END
  END mem_data_i[3]
  PIN mem_data_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 168.680 4.000 169.280 ;
    END
  END mem_data_i[4]
  PIN mem_data_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END mem_data_i[5]
  PIN mem_data_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 225.800 4.000 226.400 ;
    END
  END mem_data_i[6]
  PIN mem_data_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END mem_data_i[7]
  PIN mem_data_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 283.600 4.000 284.200 ;
    END
  END mem_data_i[8]
  PIN mem_data_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END mem_data_i[9]
  PIN mem_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END mem_data_o[0]
  PIN mem_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 335.280 4.000 335.880 ;
    END
  END mem_data_o[10]
  PIN mem_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 352.280 4.000 352.880 ;
    END
  END mem_data_o[11]
  PIN mem_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END mem_data_o[12]
  PIN mem_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.960 4.000 387.560 ;
    END
  END mem_data_o[13]
  PIN mem_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.960 4.000 404.560 ;
    END
  END mem_data_o[14]
  PIN mem_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.960 4.000 421.560 ;
    END
  END mem_data_o[15]
  PIN mem_data_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END mem_data_o[16]
  PIN mem_data_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 455.640 4.000 456.240 ;
    END
  END mem_data_o[17]
  PIN mem_data_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END mem_data_o[18]
  PIN mem_data_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 489.640 4.000 490.240 ;
    END
  END mem_data_o[19]
  PIN mem_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 76.880 4.000 77.480 ;
    END
  END mem_data_o[1]
  PIN mem_data_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END mem_data_o[20]
  PIN mem_data_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 524.320 4.000 524.920 ;
    END
  END mem_data_o[21]
  PIN mem_data_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END mem_data_o[22]
  PIN mem_data_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 559.000 4.000 559.600 ;
    END
  END mem_data_o[23]
  PIN mem_data_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 576.000 4.000 576.600 ;
    END
  END mem_data_o[24]
  PIN mem_data_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.000 4.000 593.600 ;
    END
  END mem_data_o[25]
  PIN mem_data_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 610.680 4.000 611.280 ;
    END
  END mem_data_o[26]
  PIN mem_data_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 627.680 4.000 628.280 ;
    END
  END mem_data_o[27]
  PIN mem_data_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.680 4.000 645.280 ;
    END
  END mem_data_o[28]
  PIN mem_data_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.680 4.000 662.280 ;
    END
  END mem_data_o[29]
  PIN mem_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END mem_data_o[2]
  PIN mem_data_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 679.360 4.000 679.960 ;
    END
  END mem_data_o[30]
  PIN mem_data_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 696.360 4.000 696.960 ;
    END
  END mem_data_o[31]
  PIN mem_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END mem_data_o[3]
  PIN mem_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END mem_data_o[4]
  PIN mem_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 203.360 4.000 203.960 ;
    END
  END mem_data_o[5]
  PIN mem_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.920 4.000 232.520 ;
    END
  END mem_data_o[6]
  PIN mem_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 260.480 4.000 261.080 ;
    END
  END mem_data_o[7]
  PIN mem_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END mem_data_o[8]
  PIN mem_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END mem_data_o[9]
  PIN mem_raddr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 42.880 4.000 43.480 ;
    END
  END mem_raddr_o[0]
  PIN mem_raddr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END mem_raddr_o[1]
  PIN mem_raddr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 123.120 4.000 123.720 ;
    END
  END mem_raddr_o[2]
  PIN mem_raddr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.680 4.000 152.280 ;
    END
  END mem_raddr_o[3]
  PIN mem_raddr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.240 4.000 180.840 ;
    END
  END mem_raddr_o[4]
  PIN mem_raddr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.800 4.000 209.400 ;
    END
  END mem_raddr_o[5]
  PIN mem_raddr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 237.360 4.000 237.960 ;
    END
  END mem_raddr_o[6]
  PIN mem_raddr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.920 4.000 266.520 ;
    END
  END mem_raddr_o[7]
  PIN mem_raddr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END mem_raddr_o[8]
  PIN mem_renb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 48.320 4.000 48.920 ;
    END
  END mem_renb_o[0]
  PIN mem_renb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END mem_renb_o[1]
  PIN mem_waddr_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 53.760 4.000 54.360 ;
    END
  END mem_waddr_o[0]
  PIN mem_waddr_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 93.880 4.000 94.480 ;
    END
  END mem_waddr_o[1]
  PIN mem_waddr_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END mem_waddr_o[2]
  PIN mem_waddr_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 157.120 4.000 157.720 ;
    END
  END mem_waddr_o[3]
  PIN mem_waddr_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END mem_waddr_o[4]
  PIN mem_waddr_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.920 4.000 215.520 ;
    END
  END mem_waddr_o[5]
  PIN mem_waddr_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END mem_waddr_o[6]
  PIN mem_waddr_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END mem_waddr_o[7]
  PIN mem_waddr_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END mem_waddr_o[8]
  PIN mem_wenb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END mem_wenb_o[0]
  PIN mem_wenb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END mem_wenb_o[1]
  PIN oversample_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 637.880 900.000 638.480 ;
    END
  END oversample_o[0]
  PIN oversample_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 644.680 900.000 645.280 ;
    END
  END oversample_o[1]
  PIN oversample_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 650.800 900.000 651.400 ;
    END
  END oversample_o[2]
  PIN oversample_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 656.920 900.000 657.520 ;
    END
  END oversample_o[3]
  PIN oversample_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 663.720 900.000 664.320 ;
    END
  END oversample_o[4]
  PIN oversample_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 669.840 900.000 670.440 ;
    END
  END oversample_o[5]
  PIN oversample_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 676.640 900.000 677.240 ;
    END
  END oversample_o[6]
  PIN oversample_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 682.760 900.000 683.360 ;
    END
  END oversample_o[7]
  PIN oversample_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 689.560 900.000 690.160 ;
    END
  END oversample_o[8]
  PIN oversample_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 896.000 695.680 900.000 696.280 ;
    END
  END oversample_o[9]
  PIN sinc3_en_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 872.250 696.000 872.530 700.000 ;
    END
  END sinc3_en_o[0]
  PIN sinc3_en_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.290 696.000 883.570 700.000 ;
    END
  END sinc3_en_o[1]
  PIN sinc3_en_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 894.330 696.000 894.610 700.000 ;
    END
  END sinc3_en_o[2]
  PIN vco_enb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 839.130 696.000 839.410 700.000 ;
    END
  END vco_enb_o[0]
  PIN vco_enb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 850.170 696.000 850.450 700.000 ;
    END
  END vco_enb_o[1]
  PIN vco_enb_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.210 696.000 861.490 700.000 ;
    END
  END vco_enb_o[2]
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.510 0.000 12.790 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 343.710 0.000 343.990 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.010 0.000 369.290 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 420.070 0.000 420.350 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.830 0.000 446.110 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.430 0.000 496.710 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 0.000 522.470 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 572.790 0.000 573.070 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.870 0.000 89.150 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.550 0.000 598.830 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.850 0.000 624.130 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 649.610 0.000 649.890 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.210 0.000 700.490 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 0.000 726.250 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.330 0.000 802.610 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.390 0.000 853.670 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 878.690 0.000 878.970 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 0.000 157.230 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.290 0.000 216.570 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 0.000 292.930 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.410 0.000 318.690 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.530 0.000 29.810 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 0.000 352.270 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.050 0.000 403.330 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.810 0.000 429.090 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.170 0.000 505.450 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 530.470 0.000 530.750 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.230 0.000 556.510 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.530 0.000 581.810 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.610 0.000 97.890 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.830 0.000 607.110 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 632.590 0.000 632.870 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.890 0.000 658.170 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 0.000 683.470 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.950 0.000 709.230 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.010 0.000 760.290 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.310 0.000 785.590 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 836.370 0.000 836.650 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.430 0.000 887.710 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.230 0.000 165.510 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.270 0.000 199.550 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.030 0.000 225.310 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.630 0.000 275.910 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 326.690 0.000 326.970 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.030 0.000 386.310 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 411.790 0.000 412.070 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.390 0.000 462.670 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.450 0.000 513.730 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.210 0.000 539.490 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.810 0.000 590.090 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 105.890 0.000 106.170 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 615.570 0.000 615.850 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.630 0.000 666.910 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.930 0.000 692.210 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.230 0.000 717.510 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 742.990 0.000 743.270 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 0.000 768.570 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.590 0.000 793.870 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 819.350 0.000 819.630 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.650 0.000 844.930 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 870.410 0.000 870.690 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.710 0.000 895.990 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.310 0.000 233.590 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 0.000 309.950 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.430 0.000 335.710 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 0.000 46.830 4.000 ;
    END
  END wbs_we_i
  PIN wmask_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END wmask_o[0]
  PIN wmask_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 8.200 4.000 8.800 ;
    END
  END wmask_o[1]
  PIN wmask_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END wmask_o[2]
  PIN wmask_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.760 4.000 20.360 ;
    END
  END wmask_o[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 688.400 ;
    END
  END vccd1
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 688.400 ;
    END
  END vssd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 688.400 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 792.340 10.880 793.940 688.160 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 638.740 10.880 640.340 688.160 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 485.140 10.880 486.740 688.160 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 331.540 10.880 333.140 688.160 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 177.940 10.880 179.540 688.160 ;
    END
  END vccd2
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.880 25.940 688.160 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 869.140 10.880 870.740 688.160 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 715.540 10.880 717.140 688.160 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 561.940 10.880 563.540 688.160 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 408.340 10.880 409.940 688.160 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 254.740 10.880 256.340 688.160 ;
    END
  END vssd2
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 101.140 10.880 102.740 688.160 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 795.640 10.880 797.240 688.160 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 642.040 10.880 643.640 688.160 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 488.440 10.880 490.040 688.160 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 334.840 10.880 336.440 688.160 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 181.240 10.880 182.840 688.160 ;
    END
  END vdda1
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 27.640 10.880 29.240 688.160 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 872.440 10.880 874.040 688.160 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 718.840 10.880 720.440 688.160 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 565.240 10.880 566.840 688.160 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 411.640 10.880 413.240 688.160 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 258.040 10.880 259.640 688.160 ;
    END
  END vssa1
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 104.440 10.880 106.040 688.160 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 798.940 10.880 800.540 688.160 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 645.340 10.880 646.940 688.160 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 491.740 10.880 493.340 688.160 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 338.140 10.880 339.740 688.160 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 184.540 10.880 186.140 688.160 ;
    END
  END vdda2
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 30.940 10.880 32.540 688.160 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 875.740 10.880 877.340 688.160 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 722.140 10.880 723.740 688.160 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 568.540 10.880 570.140 688.160 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 414.940 10.880 416.540 688.160 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 261.340 10.880 262.940 688.160 ;
    END
  END vssa2
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 107.740 10.880 109.340 688.160 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 5.520 8.925 895.015 688.245 ;
      LAYER met1 ;
        RECT 4.210 7.860 896.010 688.400 ;
      LAYER met2 ;
        RECT 4.240 695.720 4.870 696.845 ;
        RECT 5.710 695.720 15.450 696.845 ;
        RECT 16.290 695.720 26.490 696.845 ;
        RECT 27.330 695.720 37.530 696.845 ;
        RECT 38.370 695.720 48.570 696.845 ;
        RECT 49.410 695.720 59.610 696.845 ;
        RECT 60.450 695.720 70.650 696.845 ;
        RECT 71.490 695.720 81.690 696.845 ;
        RECT 82.530 695.720 92.270 696.845 ;
        RECT 93.110 695.720 103.310 696.845 ;
        RECT 104.150 695.720 114.350 696.845 ;
        RECT 115.190 695.720 125.390 696.845 ;
        RECT 126.230 695.720 136.430 696.845 ;
        RECT 137.270 695.720 147.470 696.845 ;
        RECT 148.310 695.720 158.510 696.845 ;
        RECT 159.350 695.720 169.090 696.845 ;
        RECT 169.930 695.720 180.130 696.845 ;
        RECT 180.970 695.720 191.170 696.845 ;
        RECT 192.010 695.720 202.210 696.845 ;
        RECT 203.050 695.720 213.250 696.845 ;
        RECT 214.090 695.720 224.290 696.845 ;
        RECT 225.130 695.720 235.330 696.845 ;
        RECT 236.170 695.720 246.370 696.845 ;
        RECT 247.210 695.720 256.950 696.845 ;
        RECT 257.790 695.720 267.990 696.845 ;
        RECT 268.830 695.720 279.030 696.845 ;
        RECT 279.870 695.720 290.070 696.845 ;
        RECT 290.910 695.720 301.110 696.845 ;
        RECT 301.950 695.720 312.150 696.845 ;
        RECT 312.990 695.720 323.190 696.845 ;
        RECT 324.030 695.720 333.770 696.845 ;
        RECT 334.610 695.720 344.810 696.845 ;
        RECT 345.650 695.720 355.850 696.845 ;
        RECT 356.690 695.720 366.890 696.845 ;
        RECT 367.730 695.720 377.930 696.845 ;
        RECT 378.770 695.720 388.970 696.845 ;
        RECT 389.810 695.720 400.010 696.845 ;
        RECT 400.850 695.720 411.050 696.845 ;
        RECT 411.890 695.720 421.630 696.845 ;
        RECT 422.470 695.720 432.670 696.845 ;
        RECT 433.510 695.720 443.710 696.845 ;
        RECT 444.550 695.720 454.750 696.845 ;
        RECT 455.590 695.720 465.790 696.845 ;
        RECT 466.630 695.720 476.830 696.845 ;
        RECT 477.670 695.720 487.870 696.845 ;
        RECT 488.710 695.720 498.450 696.845 ;
        RECT 499.290 695.720 509.490 696.845 ;
        RECT 510.330 695.720 520.530 696.845 ;
        RECT 521.370 695.720 531.570 696.845 ;
        RECT 532.410 695.720 542.610 696.845 ;
        RECT 543.450 695.720 553.650 696.845 ;
        RECT 554.490 695.720 564.690 696.845 ;
        RECT 565.530 695.720 575.730 696.845 ;
        RECT 576.570 695.720 586.310 696.845 ;
        RECT 587.150 695.720 597.350 696.845 ;
        RECT 598.190 695.720 608.390 696.845 ;
        RECT 609.230 695.720 619.430 696.845 ;
        RECT 620.270 695.720 630.470 696.845 ;
        RECT 631.310 695.720 641.510 696.845 ;
        RECT 642.350 695.720 652.550 696.845 ;
        RECT 653.390 695.720 663.130 696.845 ;
        RECT 663.970 695.720 674.170 696.845 ;
        RECT 675.010 695.720 685.210 696.845 ;
        RECT 686.050 695.720 696.250 696.845 ;
        RECT 697.090 695.720 707.290 696.845 ;
        RECT 708.130 695.720 718.330 696.845 ;
        RECT 719.170 695.720 729.370 696.845 ;
        RECT 730.210 695.720 740.410 696.845 ;
        RECT 741.250 695.720 750.990 696.845 ;
        RECT 751.830 695.720 762.030 696.845 ;
        RECT 762.870 695.720 773.070 696.845 ;
        RECT 773.910 695.720 784.110 696.845 ;
        RECT 784.950 695.720 795.150 696.845 ;
        RECT 795.990 695.720 806.190 696.845 ;
        RECT 807.030 695.720 817.230 696.845 ;
        RECT 818.070 695.720 827.810 696.845 ;
        RECT 828.650 695.720 838.850 696.845 ;
        RECT 839.690 695.720 849.890 696.845 ;
        RECT 850.730 695.720 860.930 696.845 ;
        RECT 861.770 695.720 871.970 696.845 ;
        RECT 872.810 695.720 883.010 696.845 ;
        RECT 883.850 695.720 894.050 696.845 ;
        RECT 894.890 695.720 895.980 696.845 ;
        RECT 4.240 4.280 895.980 695.720 ;
        RECT 4.790 2.875 12.230 4.280 ;
        RECT 13.070 2.875 20.510 4.280 ;
        RECT 21.350 2.875 29.250 4.280 ;
        RECT 30.090 2.875 37.530 4.280 ;
        RECT 38.370 2.875 46.270 4.280 ;
        RECT 47.110 2.875 54.550 4.280 ;
        RECT 55.390 2.875 63.290 4.280 ;
        RECT 64.130 2.875 71.570 4.280 ;
        RECT 72.410 2.875 80.310 4.280 ;
        RECT 81.150 2.875 88.590 4.280 ;
        RECT 89.430 2.875 97.330 4.280 ;
        RECT 98.170 2.875 105.610 4.280 ;
        RECT 106.450 2.875 114.350 4.280 ;
        RECT 115.190 2.875 122.630 4.280 ;
        RECT 123.470 2.875 130.910 4.280 ;
        RECT 131.750 2.875 139.650 4.280 ;
        RECT 140.490 2.875 147.930 4.280 ;
        RECT 148.770 2.875 156.670 4.280 ;
        RECT 157.510 2.875 164.950 4.280 ;
        RECT 165.790 2.875 173.690 4.280 ;
        RECT 174.530 2.875 181.970 4.280 ;
        RECT 182.810 2.875 190.710 4.280 ;
        RECT 191.550 2.875 198.990 4.280 ;
        RECT 199.830 2.875 207.730 4.280 ;
        RECT 208.570 2.875 216.010 4.280 ;
        RECT 216.850 2.875 224.750 4.280 ;
        RECT 225.590 2.875 233.030 4.280 ;
        RECT 233.870 2.875 241.310 4.280 ;
        RECT 242.150 2.875 250.050 4.280 ;
        RECT 250.890 2.875 258.330 4.280 ;
        RECT 259.170 2.875 267.070 4.280 ;
        RECT 267.910 2.875 275.350 4.280 ;
        RECT 276.190 2.875 284.090 4.280 ;
        RECT 284.930 2.875 292.370 4.280 ;
        RECT 293.210 2.875 301.110 4.280 ;
        RECT 301.950 2.875 309.390 4.280 ;
        RECT 310.230 2.875 318.130 4.280 ;
        RECT 318.970 2.875 326.410 4.280 ;
        RECT 327.250 2.875 335.150 4.280 ;
        RECT 335.990 2.875 343.430 4.280 ;
        RECT 344.270 2.875 351.710 4.280 ;
        RECT 352.550 2.875 360.450 4.280 ;
        RECT 361.290 2.875 368.730 4.280 ;
        RECT 369.570 2.875 377.470 4.280 ;
        RECT 378.310 2.875 385.750 4.280 ;
        RECT 386.590 2.875 394.490 4.280 ;
        RECT 395.330 2.875 402.770 4.280 ;
        RECT 403.610 2.875 411.510 4.280 ;
        RECT 412.350 2.875 419.790 4.280 ;
        RECT 420.630 2.875 428.530 4.280 ;
        RECT 429.370 2.875 436.810 4.280 ;
        RECT 437.650 2.875 445.550 4.280 ;
        RECT 446.390 2.875 453.830 4.280 ;
        RECT 454.670 2.875 462.110 4.280 ;
        RECT 462.950 2.875 470.850 4.280 ;
        RECT 471.690 2.875 479.130 4.280 ;
        RECT 479.970 2.875 487.870 4.280 ;
        RECT 488.710 2.875 496.150 4.280 ;
        RECT 496.990 2.875 504.890 4.280 ;
        RECT 505.730 2.875 513.170 4.280 ;
        RECT 514.010 2.875 521.910 4.280 ;
        RECT 522.750 2.875 530.190 4.280 ;
        RECT 531.030 2.875 538.930 4.280 ;
        RECT 539.770 2.875 547.210 4.280 ;
        RECT 548.050 2.875 555.950 4.280 ;
        RECT 556.790 2.875 564.230 4.280 ;
        RECT 565.070 2.875 572.510 4.280 ;
        RECT 573.350 2.875 581.250 4.280 ;
        RECT 582.090 2.875 589.530 4.280 ;
        RECT 590.370 2.875 598.270 4.280 ;
        RECT 599.110 2.875 606.550 4.280 ;
        RECT 607.390 2.875 615.290 4.280 ;
        RECT 616.130 2.875 623.570 4.280 ;
        RECT 624.410 2.875 632.310 4.280 ;
        RECT 633.150 2.875 640.590 4.280 ;
        RECT 641.430 2.875 649.330 4.280 ;
        RECT 650.170 2.875 657.610 4.280 ;
        RECT 658.450 2.875 666.350 4.280 ;
        RECT 667.190 2.875 674.630 4.280 ;
        RECT 675.470 2.875 682.910 4.280 ;
        RECT 683.750 2.875 691.650 4.280 ;
        RECT 692.490 2.875 699.930 4.280 ;
        RECT 700.770 2.875 708.670 4.280 ;
        RECT 709.510 2.875 716.950 4.280 ;
        RECT 717.790 2.875 725.690 4.280 ;
        RECT 726.530 2.875 733.970 4.280 ;
        RECT 734.810 2.875 742.710 4.280 ;
        RECT 743.550 2.875 750.990 4.280 ;
        RECT 751.830 2.875 759.730 4.280 ;
        RECT 760.570 2.875 768.010 4.280 ;
        RECT 768.850 2.875 776.750 4.280 ;
        RECT 777.590 2.875 785.030 4.280 ;
        RECT 785.870 2.875 793.310 4.280 ;
        RECT 794.150 2.875 802.050 4.280 ;
        RECT 802.890 2.875 810.330 4.280 ;
        RECT 811.170 2.875 819.070 4.280 ;
        RECT 819.910 2.875 827.350 4.280 ;
        RECT 828.190 2.875 836.090 4.280 ;
        RECT 836.930 2.875 844.370 4.280 ;
        RECT 845.210 2.875 853.110 4.280 ;
        RECT 853.950 2.875 861.390 4.280 ;
        RECT 862.230 2.875 870.130 4.280 ;
        RECT 870.970 2.875 878.410 4.280 ;
        RECT 879.250 2.875 887.150 4.280 ;
        RECT 887.990 2.875 895.430 4.280 ;
      LAYER met3 ;
        RECT 4.400 696.680 896.000 696.825 ;
        RECT 4.400 695.960 895.600 696.680 ;
        RECT 4.000 695.280 895.600 695.960 ;
        RECT 4.000 691.920 896.000 695.280 ;
        RECT 4.400 690.560 896.000 691.920 ;
        RECT 4.400 690.520 895.600 690.560 ;
        RECT 4.000 689.160 895.600 690.520 ;
        RECT 4.000 685.800 896.000 689.160 ;
        RECT 4.400 684.400 896.000 685.800 ;
        RECT 4.000 683.760 896.000 684.400 ;
        RECT 4.000 682.360 895.600 683.760 ;
        RECT 4.000 680.360 896.000 682.360 ;
        RECT 4.400 678.960 896.000 680.360 ;
        RECT 4.000 677.640 896.000 678.960 ;
        RECT 4.000 676.240 895.600 677.640 ;
        RECT 4.000 674.240 896.000 676.240 ;
        RECT 4.400 672.840 896.000 674.240 ;
        RECT 4.000 670.840 896.000 672.840 ;
        RECT 4.000 669.440 895.600 670.840 ;
        RECT 4.000 668.800 896.000 669.440 ;
        RECT 4.400 667.400 896.000 668.800 ;
        RECT 4.000 664.720 896.000 667.400 ;
        RECT 4.000 663.320 895.600 664.720 ;
        RECT 4.000 662.680 896.000 663.320 ;
        RECT 4.400 661.280 896.000 662.680 ;
        RECT 4.000 657.920 896.000 661.280 ;
        RECT 4.000 657.240 895.600 657.920 ;
        RECT 4.400 656.520 895.600 657.240 ;
        RECT 4.400 655.840 896.000 656.520 ;
        RECT 4.000 651.800 896.000 655.840 ;
        RECT 4.400 650.400 895.600 651.800 ;
        RECT 4.000 645.680 896.000 650.400 ;
        RECT 4.400 644.280 895.600 645.680 ;
        RECT 4.000 640.240 896.000 644.280 ;
        RECT 4.400 638.880 896.000 640.240 ;
        RECT 4.400 638.840 895.600 638.880 ;
        RECT 4.000 637.480 895.600 638.840 ;
        RECT 4.000 634.120 896.000 637.480 ;
        RECT 4.400 632.760 896.000 634.120 ;
        RECT 4.400 632.720 895.600 632.760 ;
        RECT 4.000 631.360 895.600 632.720 ;
        RECT 4.000 628.680 896.000 631.360 ;
        RECT 4.400 627.280 896.000 628.680 ;
        RECT 4.000 625.960 896.000 627.280 ;
        RECT 4.000 624.560 895.600 625.960 ;
        RECT 4.000 622.560 896.000 624.560 ;
        RECT 4.400 621.160 896.000 622.560 ;
        RECT 4.000 619.840 896.000 621.160 ;
        RECT 4.000 618.440 895.600 619.840 ;
        RECT 4.000 617.120 896.000 618.440 ;
        RECT 4.400 615.720 896.000 617.120 ;
        RECT 4.000 613.040 896.000 615.720 ;
        RECT 4.000 611.680 895.600 613.040 ;
        RECT 4.400 611.640 895.600 611.680 ;
        RECT 4.400 610.280 896.000 611.640 ;
        RECT 4.000 606.920 896.000 610.280 ;
        RECT 4.000 605.560 895.600 606.920 ;
        RECT 4.400 605.520 895.600 605.560 ;
        RECT 4.400 604.160 896.000 605.520 ;
        RECT 4.000 600.120 896.000 604.160 ;
        RECT 4.400 598.720 895.600 600.120 ;
        RECT 4.000 594.000 896.000 598.720 ;
        RECT 4.400 592.600 895.600 594.000 ;
        RECT 4.000 588.560 896.000 592.600 ;
        RECT 4.400 587.880 896.000 588.560 ;
        RECT 4.400 587.160 895.600 587.880 ;
        RECT 4.000 586.480 895.600 587.160 ;
        RECT 4.000 582.440 896.000 586.480 ;
        RECT 4.400 581.080 896.000 582.440 ;
        RECT 4.400 581.040 895.600 581.080 ;
        RECT 4.000 579.680 895.600 581.040 ;
        RECT 4.000 577.000 896.000 579.680 ;
        RECT 4.400 575.600 896.000 577.000 ;
        RECT 4.000 574.960 896.000 575.600 ;
        RECT 4.000 573.560 895.600 574.960 ;
        RECT 4.000 571.560 896.000 573.560 ;
        RECT 4.400 570.160 896.000 571.560 ;
        RECT 4.000 568.160 896.000 570.160 ;
        RECT 4.000 566.760 895.600 568.160 ;
        RECT 4.000 565.440 896.000 566.760 ;
        RECT 4.400 564.040 896.000 565.440 ;
        RECT 4.000 562.040 896.000 564.040 ;
        RECT 4.000 560.640 895.600 562.040 ;
        RECT 4.000 560.000 896.000 560.640 ;
        RECT 4.400 558.600 896.000 560.000 ;
        RECT 4.000 555.240 896.000 558.600 ;
        RECT 4.000 553.880 895.600 555.240 ;
        RECT 4.400 553.840 895.600 553.880 ;
        RECT 4.400 552.480 896.000 553.840 ;
        RECT 4.000 549.120 896.000 552.480 ;
        RECT 4.000 548.440 895.600 549.120 ;
        RECT 4.400 547.720 895.600 548.440 ;
        RECT 4.400 547.040 896.000 547.720 ;
        RECT 4.000 542.320 896.000 547.040 ;
        RECT 4.400 540.920 895.600 542.320 ;
        RECT 4.000 536.880 896.000 540.920 ;
        RECT 4.400 536.200 896.000 536.880 ;
        RECT 4.400 535.480 895.600 536.200 ;
        RECT 4.000 534.800 895.600 535.480 ;
        RECT 4.000 530.760 896.000 534.800 ;
        RECT 4.400 530.080 896.000 530.760 ;
        RECT 4.400 529.360 895.600 530.080 ;
        RECT 4.000 528.680 895.600 529.360 ;
        RECT 4.000 525.320 896.000 528.680 ;
        RECT 4.400 523.920 896.000 525.320 ;
        RECT 4.000 523.280 896.000 523.920 ;
        RECT 4.000 521.880 895.600 523.280 ;
        RECT 4.000 519.880 896.000 521.880 ;
        RECT 4.400 518.480 896.000 519.880 ;
        RECT 4.000 517.160 896.000 518.480 ;
        RECT 4.000 515.760 895.600 517.160 ;
        RECT 4.000 513.760 896.000 515.760 ;
        RECT 4.400 512.360 896.000 513.760 ;
        RECT 4.000 510.360 896.000 512.360 ;
        RECT 4.000 508.960 895.600 510.360 ;
        RECT 4.000 508.320 896.000 508.960 ;
        RECT 4.400 506.920 896.000 508.320 ;
        RECT 4.000 504.240 896.000 506.920 ;
        RECT 4.000 502.840 895.600 504.240 ;
        RECT 4.000 502.200 896.000 502.840 ;
        RECT 4.400 500.800 896.000 502.200 ;
        RECT 4.000 497.440 896.000 500.800 ;
        RECT 4.000 496.760 895.600 497.440 ;
        RECT 4.400 496.040 895.600 496.760 ;
        RECT 4.400 495.360 896.000 496.040 ;
        RECT 4.000 491.320 896.000 495.360 ;
        RECT 4.000 490.640 895.600 491.320 ;
        RECT 4.400 489.920 895.600 490.640 ;
        RECT 4.400 489.240 896.000 489.920 ;
        RECT 4.000 485.200 896.000 489.240 ;
        RECT 4.400 483.800 895.600 485.200 ;
        RECT 4.000 479.760 896.000 483.800 ;
        RECT 4.400 478.400 896.000 479.760 ;
        RECT 4.400 478.360 895.600 478.400 ;
        RECT 4.000 477.000 895.600 478.360 ;
        RECT 4.000 473.640 896.000 477.000 ;
        RECT 4.400 472.280 896.000 473.640 ;
        RECT 4.400 472.240 895.600 472.280 ;
        RECT 4.000 470.880 895.600 472.240 ;
        RECT 4.000 468.200 896.000 470.880 ;
        RECT 4.400 466.800 896.000 468.200 ;
        RECT 4.000 465.480 896.000 466.800 ;
        RECT 4.000 464.080 895.600 465.480 ;
        RECT 4.000 462.080 896.000 464.080 ;
        RECT 4.400 460.680 896.000 462.080 ;
        RECT 4.000 459.360 896.000 460.680 ;
        RECT 4.000 457.960 895.600 459.360 ;
        RECT 4.000 456.640 896.000 457.960 ;
        RECT 4.400 455.240 896.000 456.640 ;
        RECT 4.000 452.560 896.000 455.240 ;
        RECT 4.000 451.160 895.600 452.560 ;
        RECT 4.000 450.520 896.000 451.160 ;
        RECT 4.400 449.120 896.000 450.520 ;
        RECT 4.000 446.440 896.000 449.120 ;
        RECT 4.000 445.080 895.600 446.440 ;
        RECT 4.400 445.040 895.600 445.080 ;
        RECT 4.400 443.680 896.000 445.040 ;
        RECT 4.000 439.640 896.000 443.680 ;
        RECT 4.400 438.240 895.600 439.640 ;
        RECT 4.000 433.520 896.000 438.240 ;
        RECT 4.400 432.120 895.600 433.520 ;
        RECT 4.000 428.080 896.000 432.120 ;
        RECT 4.400 427.400 896.000 428.080 ;
        RECT 4.400 426.680 895.600 427.400 ;
        RECT 4.000 426.000 895.600 426.680 ;
        RECT 4.000 421.960 896.000 426.000 ;
        RECT 4.400 420.600 896.000 421.960 ;
        RECT 4.400 420.560 895.600 420.600 ;
        RECT 4.000 419.200 895.600 420.560 ;
        RECT 4.000 416.520 896.000 419.200 ;
        RECT 4.400 415.120 896.000 416.520 ;
        RECT 4.000 414.480 896.000 415.120 ;
        RECT 4.000 413.080 895.600 414.480 ;
        RECT 4.000 410.400 896.000 413.080 ;
        RECT 4.400 409.000 896.000 410.400 ;
        RECT 4.000 407.680 896.000 409.000 ;
        RECT 4.000 406.280 895.600 407.680 ;
        RECT 4.000 404.960 896.000 406.280 ;
        RECT 4.400 403.560 896.000 404.960 ;
        RECT 4.000 401.560 896.000 403.560 ;
        RECT 4.000 400.160 895.600 401.560 ;
        RECT 4.000 398.840 896.000 400.160 ;
        RECT 4.400 397.440 896.000 398.840 ;
        RECT 4.000 394.760 896.000 397.440 ;
        RECT 4.000 393.400 895.600 394.760 ;
        RECT 4.400 393.360 895.600 393.400 ;
        RECT 4.400 392.000 896.000 393.360 ;
        RECT 4.000 388.640 896.000 392.000 ;
        RECT 4.000 387.960 895.600 388.640 ;
        RECT 4.400 387.240 895.600 387.960 ;
        RECT 4.400 386.560 896.000 387.240 ;
        RECT 4.000 381.840 896.000 386.560 ;
        RECT 4.400 380.440 895.600 381.840 ;
        RECT 4.000 376.400 896.000 380.440 ;
        RECT 4.400 375.720 896.000 376.400 ;
        RECT 4.400 375.000 895.600 375.720 ;
        RECT 4.000 374.320 895.600 375.000 ;
        RECT 4.000 370.280 896.000 374.320 ;
        RECT 4.400 369.600 896.000 370.280 ;
        RECT 4.400 368.880 895.600 369.600 ;
        RECT 4.000 368.200 895.600 368.880 ;
        RECT 4.000 364.840 896.000 368.200 ;
        RECT 4.400 363.440 896.000 364.840 ;
        RECT 4.000 362.800 896.000 363.440 ;
        RECT 4.000 361.400 895.600 362.800 ;
        RECT 4.000 358.720 896.000 361.400 ;
        RECT 4.400 357.320 896.000 358.720 ;
        RECT 4.000 356.680 896.000 357.320 ;
        RECT 4.000 355.280 895.600 356.680 ;
        RECT 4.000 353.280 896.000 355.280 ;
        RECT 4.400 351.880 896.000 353.280 ;
        RECT 4.000 349.880 896.000 351.880 ;
        RECT 4.000 348.480 895.600 349.880 ;
        RECT 4.000 347.840 896.000 348.480 ;
        RECT 4.400 346.440 896.000 347.840 ;
        RECT 4.000 343.760 896.000 346.440 ;
        RECT 4.000 342.360 895.600 343.760 ;
        RECT 4.000 341.720 896.000 342.360 ;
        RECT 4.400 340.320 896.000 341.720 ;
        RECT 4.000 336.960 896.000 340.320 ;
        RECT 4.000 336.280 895.600 336.960 ;
        RECT 4.400 335.560 895.600 336.280 ;
        RECT 4.400 334.880 896.000 335.560 ;
        RECT 4.000 330.840 896.000 334.880 ;
        RECT 4.000 330.160 895.600 330.840 ;
        RECT 4.400 329.440 895.600 330.160 ;
        RECT 4.400 328.760 896.000 329.440 ;
        RECT 4.000 324.720 896.000 328.760 ;
        RECT 4.400 323.320 895.600 324.720 ;
        RECT 4.000 318.600 896.000 323.320 ;
        RECT 4.400 317.920 896.000 318.600 ;
        RECT 4.400 317.200 895.600 317.920 ;
        RECT 4.000 316.520 895.600 317.200 ;
        RECT 4.000 313.160 896.000 316.520 ;
        RECT 4.400 311.800 896.000 313.160 ;
        RECT 4.400 311.760 895.600 311.800 ;
        RECT 4.000 310.400 895.600 311.760 ;
        RECT 4.000 307.720 896.000 310.400 ;
        RECT 4.400 306.320 896.000 307.720 ;
        RECT 4.000 305.000 896.000 306.320 ;
        RECT 4.000 303.600 895.600 305.000 ;
        RECT 4.000 301.600 896.000 303.600 ;
        RECT 4.400 300.200 896.000 301.600 ;
        RECT 4.000 298.880 896.000 300.200 ;
        RECT 4.000 297.480 895.600 298.880 ;
        RECT 4.000 296.160 896.000 297.480 ;
        RECT 4.400 294.760 896.000 296.160 ;
        RECT 4.000 292.080 896.000 294.760 ;
        RECT 4.000 290.680 895.600 292.080 ;
        RECT 4.000 290.040 896.000 290.680 ;
        RECT 4.400 288.640 896.000 290.040 ;
        RECT 4.000 285.960 896.000 288.640 ;
        RECT 4.000 284.600 895.600 285.960 ;
        RECT 4.400 284.560 895.600 284.600 ;
        RECT 4.400 283.200 896.000 284.560 ;
        RECT 4.000 279.160 896.000 283.200 ;
        RECT 4.000 278.480 895.600 279.160 ;
        RECT 4.400 277.760 895.600 278.480 ;
        RECT 4.400 277.080 896.000 277.760 ;
        RECT 4.000 273.040 896.000 277.080 ;
        RECT 4.400 271.640 895.600 273.040 ;
        RECT 4.000 266.920 896.000 271.640 ;
        RECT 4.400 265.520 895.600 266.920 ;
        RECT 4.000 261.480 896.000 265.520 ;
        RECT 4.400 260.120 896.000 261.480 ;
        RECT 4.400 260.080 895.600 260.120 ;
        RECT 4.000 258.720 895.600 260.080 ;
        RECT 4.000 256.040 896.000 258.720 ;
        RECT 4.400 254.640 896.000 256.040 ;
        RECT 4.000 254.000 896.000 254.640 ;
        RECT 4.000 252.600 895.600 254.000 ;
        RECT 4.000 249.920 896.000 252.600 ;
        RECT 4.400 248.520 896.000 249.920 ;
        RECT 4.000 247.200 896.000 248.520 ;
        RECT 4.000 245.800 895.600 247.200 ;
        RECT 4.000 244.480 896.000 245.800 ;
        RECT 4.400 243.080 896.000 244.480 ;
        RECT 4.000 241.080 896.000 243.080 ;
        RECT 4.000 239.680 895.600 241.080 ;
        RECT 4.000 238.360 896.000 239.680 ;
        RECT 4.400 236.960 896.000 238.360 ;
        RECT 4.000 234.280 896.000 236.960 ;
        RECT 4.000 232.920 895.600 234.280 ;
        RECT 4.400 232.880 895.600 232.920 ;
        RECT 4.400 231.520 896.000 232.880 ;
        RECT 4.000 228.160 896.000 231.520 ;
        RECT 4.000 226.800 895.600 228.160 ;
        RECT 4.400 226.760 895.600 226.800 ;
        RECT 4.400 225.400 896.000 226.760 ;
        RECT 4.000 221.360 896.000 225.400 ;
        RECT 4.400 219.960 895.600 221.360 ;
        RECT 4.000 215.920 896.000 219.960 ;
        RECT 4.400 215.240 896.000 215.920 ;
        RECT 4.400 214.520 895.600 215.240 ;
        RECT 4.000 213.840 895.600 214.520 ;
        RECT 4.000 209.800 896.000 213.840 ;
        RECT 4.400 209.120 896.000 209.800 ;
        RECT 4.400 208.400 895.600 209.120 ;
        RECT 4.000 207.720 895.600 208.400 ;
        RECT 4.000 204.360 896.000 207.720 ;
        RECT 4.400 202.960 896.000 204.360 ;
        RECT 4.000 202.320 896.000 202.960 ;
        RECT 4.000 200.920 895.600 202.320 ;
        RECT 4.000 198.240 896.000 200.920 ;
        RECT 4.400 196.840 896.000 198.240 ;
        RECT 4.000 196.200 896.000 196.840 ;
        RECT 4.000 194.800 895.600 196.200 ;
        RECT 4.000 192.800 896.000 194.800 ;
        RECT 4.400 191.400 896.000 192.800 ;
        RECT 4.000 189.400 896.000 191.400 ;
        RECT 4.000 188.000 895.600 189.400 ;
        RECT 4.000 186.680 896.000 188.000 ;
        RECT 4.400 185.280 896.000 186.680 ;
        RECT 4.000 183.280 896.000 185.280 ;
        RECT 4.000 181.880 895.600 183.280 ;
        RECT 4.000 181.240 896.000 181.880 ;
        RECT 4.400 179.840 896.000 181.240 ;
        RECT 4.000 176.480 896.000 179.840 ;
        RECT 4.000 175.800 895.600 176.480 ;
        RECT 4.400 175.080 895.600 175.800 ;
        RECT 4.400 174.400 896.000 175.080 ;
        RECT 4.000 170.360 896.000 174.400 ;
        RECT 4.000 169.680 895.600 170.360 ;
        RECT 4.400 168.960 895.600 169.680 ;
        RECT 4.400 168.280 896.000 168.960 ;
        RECT 4.000 164.240 896.000 168.280 ;
        RECT 4.400 162.840 895.600 164.240 ;
        RECT 4.000 158.120 896.000 162.840 ;
        RECT 4.400 157.440 896.000 158.120 ;
        RECT 4.400 156.720 895.600 157.440 ;
        RECT 4.000 156.040 895.600 156.720 ;
        RECT 4.000 152.680 896.000 156.040 ;
        RECT 4.400 151.320 896.000 152.680 ;
        RECT 4.400 151.280 895.600 151.320 ;
        RECT 4.000 149.920 895.600 151.280 ;
        RECT 4.000 146.560 896.000 149.920 ;
        RECT 4.400 145.160 896.000 146.560 ;
        RECT 4.000 144.520 896.000 145.160 ;
        RECT 4.000 143.120 895.600 144.520 ;
        RECT 4.000 141.120 896.000 143.120 ;
        RECT 4.400 139.720 896.000 141.120 ;
        RECT 4.000 138.400 896.000 139.720 ;
        RECT 4.000 137.000 895.600 138.400 ;
        RECT 4.000 135.000 896.000 137.000 ;
        RECT 4.400 133.600 896.000 135.000 ;
        RECT 4.000 131.600 896.000 133.600 ;
        RECT 4.000 130.200 895.600 131.600 ;
        RECT 4.000 129.560 896.000 130.200 ;
        RECT 4.400 128.160 896.000 129.560 ;
        RECT 4.000 125.480 896.000 128.160 ;
        RECT 4.000 124.120 895.600 125.480 ;
        RECT 4.400 124.080 895.600 124.120 ;
        RECT 4.400 122.720 896.000 124.080 ;
        RECT 4.000 118.680 896.000 122.720 ;
        RECT 4.000 118.000 895.600 118.680 ;
        RECT 4.400 117.280 895.600 118.000 ;
        RECT 4.400 116.600 896.000 117.280 ;
        RECT 4.000 112.560 896.000 116.600 ;
        RECT 4.400 111.160 895.600 112.560 ;
        RECT 4.000 106.440 896.000 111.160 ;
        RECT 4.400 105.040 895.600 106.440 ;
        RECT 4.000 101.000 896.000 105.040 ;
        RECT 4.400 99.640 896.000 101.000 ;
        RECT 4.400 99.600 895.600 99.640 ;
        RECT 4.000 98.240 895.600 99.600 ;
        RECT 4.000 94.880 896.000 98.240 ;
        RECT 4.400 93.520 896.000 94.880 ;
        RECT 4.400 93.480 895.600 93.520 ;
        RECT 4.000 92.120 895.600 93.480 ;
        RECT 4.000 89.440 896.000 92.120 ;
        RECT 4.400 88.040 896.000 89.440 ;
        RECT 4.000 86.720 896.000 88.040 ;
        RECT 4.000 85.320 895.600 86.720 ;
        RECT 4.000 84.000 896.000 85.320 ;
        RECT 4.400 82.600 896.000 84.000 ;
        RECT 4.000 80.600 896.000 82.600 ;
        RECT 4.000 79.200 895.600 80.600 ;
        RECT 4.000 77.880 896.000 79.200 ;
        RECT 4.400 76.480 896.000 77.880 ;
        RECT 4.000 73.800 896.000 76.480 ;
        RECT 4.000 72.440 895.600 73.800 ;
        RECT 4.400 72.400 895.600 72.440 ;
        RECT 4.400 71.040 896.000 72.400 ;
        RECT 4.000 67.680 896.000 71.040 ;
        RECT 4.000 66.320 895.600 67.680 ;
        RECT 4.400 66.280 895.600 66.320 ;
        RECT 4.400 64.920 896.000 66.280 ;
        RECT 4.000 60.880 896.000 64.920 ;
        RECT 4.400 59.480 895.600 60.880 ;
        RECT 4.000 54.760 896.000 59.480 ;
        RECT 4.400 53.360 895.600 54.760 ;
        RECT 4.000 49.320 896.000 53.360 ;
        RECT 4.400 48.640 896.000 49.320 ;
        RECT 4.400 47.920 895.600 48.640 ;
        RECT 4.000 47.240 895.600 47.920 ;
        RECT 4.000 43.880 896.000 47.240 ;
        RECT 4.400 42.480 896.000 43.880 ;
        RECT 4.000 41.840 896.000 42.480 ;
        RECT 4.000 40.440 895.600 41.840 ;
        RECT 4.000 37.760 896.000 40.440 ;
        RECT 4.400 36.360 896.000 37.760 ;
        RECT 4.000 35.720 896.000 36.360 ;
        RECT 4.000 34.320 895.600 35.720 ;
        RECT 4.000 32.320 896.000 34.320 ;
        RECT 4.400 30.920 896.000 32.320 ;
        RECT 4.000 28.920 896.000 30.920 ;
        RECT 4.000 27.520 895.600 28.920 ;
        RECT 4.000 26.200 896.000 27.520 ;
        RECT 4.400 24.800 896.000 26.200 ;
        RECT 4.000 22.800 896.000 24.800 ;
        RECT 4.000 21.400 895.600 22.800 ;
        RECT 4.000 20.760 896.000 21.400 ;
        RECT 4.400 19.360 896.000 20.760 ;
        RECT 4.000 16.000 896.000 19.360 ;
        RECT 4.000 14.640 895.600 16.000 ;
        RECT 4.400 14.600 895.600 14.640 ;
        RECT 4.400 13.240 896.000 14.600 ;
        RECT 4.000 9.880 896.000 13.240 ;
        RECT 4.000 9.200 895.600 9.880 ;
        RECT 4.400 8.480 895.600 9.200 ;
        RECT 4.400 7.800 896.000 8.480 ;
        RECT 4.000 3.760 896.000 7.800 ;
        RECT 4.400 2.895 895.600 3.760 ;
      LAYER met4 ;
        RECT 400.035 14.455 404.640 685.945 ;
        RECT 407.040 14.455 407.940 685.945 ;
        RECT 410.340 14.455 411.240 685.945 ;
        RECT 413.640 14.455 414.540 685.945 ;
        RECT 416.940 14.455 481.440 685.945 ;
        RECT 483.840 14.455 484.740 685.945 ;
        RECT 487.140 14.455 488.040 685.945 ;
        RECT 490.440 14.455 491.340 685.945 ;
        RECT 493.740 14.455 558.240 685.945 ;
        RECT 560.640 14.455 561.540 685.945 ;
        RECT 563.940 14.455 564.840 685.945 ;
        RECT 567.240 14.455 568.140 685.945 ;
        RECT 570.540 14.455 635.040 685.945 ;
        RECT 637.440 14.455 638.340 685.945 ;
        RECT 640.740 14.455 641.640 685.945 ;
        RECT 644.040 14.455 644.940 685.945 ;
        RECT 647.340 14.455 711.840 685.945 ;
        RECT 714.240 14.455 715.140 685.945 ;
        RECT 717.540 14.455 718.440 685.945 ;
        RECT 720.840 14.455 721.740 685.945 ;
        RECT 724.140 14.455 788.640 685.945 ;
        RECT 791.040 14.455 791.940 685.945 ;
        RECT 794.340 14.455 795.240 685.945 ;
        RECT 797.640 14.455 798.540 685.945 ;
        RECT 800.940 14.455 865.440 685.945 ;
        RECT 867.840 14.455 868.740 685.945 ;
        RECT 871.140 14.455 872.040 685.945 ;
        RECT 874.440 14.455 875.340 685.945 ;
        RECT 877.740 14.455 889.345 685.945 ;
  END
END vco_adc_wrapper
END LIBRARY

