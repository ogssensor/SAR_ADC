magic
tech sky130A
magscale 1 2
timestamp 1621791239
<< obsli1 >>
rect 1104 2159 178848 117521
<< obsm1 >>
rect 658 1028 179294 118108
<< metal2 >>
rect 662 119200 718 120000
rect 2042 119200 2098 120000
rect 3514 119200 3570 120000
rect 4894 119200 4950 120000
rect 6366 119200 6422 120000
rect 7838 119200 7894 120000
rect 9218 119200 9274 120000
rect 10690 119200 10746 120000
rect 12162 119200 12218 120000
rect 13542 119200 13598 120000
rect 15014 119200 15070 120000
rect 16486 119200 16542 120000
rect 17866 119200 17922 120000
rect 19338 119200 19394 120000
rect 20810 119200 20866 120000
rect 22190 119200 22246 120000
rect 23662 119200 23718 120000
rect 25134 119200 25190 120000
rect 26514 119200 26570 120000
rect 27986 119200 28042 120000
rect 29458 119200 29514 120000
rect 30838 119200 30894 120000
rect 32310 119200 32366 120000
rect 33782 119200 33838 120000
rect 35162 119200 35218 120000
rect 36634 119200 36690 120000
rect 38106 119200 38162 120000
rect 39486 119200 39542 120000
rect 40958 119200 41014 120000
rect 42430 119200 42486 120000
rect 43810 119200 43866 120000
rect 45282 119200 45338 120000
rect 46662 119200 46718 120000
rect 48134 119200 48190 120000
rect 49606 119200 49662 120000
rect 50986 119200 51042 120000
rect 52458 119200 52514 120000
rect 53930 119200 53986 120000
rect 55310 119200 55366 120000
rect 56782 119200 56838 120000
rect 58254 119200 58310 120000
rect 59634 119200 59690 120000
rect 61106 119200 61162 120000
rect 62578 119200 62634 120000
rect 63958 119200 64014 120000
rect 65430 119200 65486 120000
rect 66902 119200 66958 120000
rect 68282 119200 68338 120000
rect 69754 119200 69810 120000
rect 71226 119200 71282 120000
rect 72606 119200 72662 120000
rect 74078 119200 74134 120000
rect 75550 119200 75606 120000
rect 76930 119200 76986 120000
rect 78402 119200 78458 120000
rect 79874 119200 79930 120000
rect 81254 119200 81310 120000
rect 82726 119200 82782 120000
rect 84198 119200 84254 120000
rect 85578 119200 85634 120000
rect 87050 119200 87106 120000
rect 88522 119200 88578 120000
rect 89902 119200 89958 120000
rect 91374 119200 91430 120000
rect 92754 119200 92810 120000
rect 94226 119200 94282 120000
rect 95698 119200 95754 120000
rect 97078 119200 97134 120000
rect 98550 119200 98606 120000
rect 100022 119200 100078 120000
rect 101402 119200 101458 120000
rect 102874 119200 102930 120000
rect 104346 119200 104402 120000
rect 105726 119200 105782 120000
rect 107198 119200 107254 120000
rect 108670 119200 108726 120000
rect 110050 119200 110106 120000
rect 111522 119200 111578 120000
rect 112994 119200 113050 120000
rect 114374 119200 114430 120000
rect 115846 119200 115902 120000
rect 117318 119200 117374 120000
rect 118698 119200 118754 120000
rect 120170 119200 120226 120000
rect 121642 119200 121698 120000
rect 123022 119200 123078 120000
rect 124494 119200 124550 120000
rect 125966 119200 126022 120000
rect 127346 119200 127402 120000
rect 128818 119200 128874 120000
rect 130290 119200 130346 120000
rect 131670 119200 131726 120000
rect 133142 119200 133198 120000
rect 134614 119200 134670 120000
rect 135994 119200 136050 120000
rect 137466 119200 137522 120000
rect 138846 119200 138902 120000
rect 140318 119200 140374 120000
rect 141790 119200 141846 120000
rect 143170 119200 143226 120000
rect 144642 119200 144698 120000
rect 146114 119200 146170 120000
rect 147494 119200 147550 120000
rect 148966 119200 149022 120000
rect 150438 119200 150494 120000
rect 151818 119200 151874 120000
rect 153290 119200 153346 120000
rect 154762 119200 154818 120000
rect 156142 119200 156198 120000
rect 157614 119200 157670 120000
rect 159086 119200 159142 120000
rect 160466 119200 160522 120000
rect 161938 119200 161994 120000
rect 163410 119200 163466 120000
rect 164790 119200 164846 120000
rect 166262 119200 166318 120000
rect 167734 119200 167790 120000
rect 169114 119200 169170 120000
rect 170586 119200 170642 120000
rect 172058 119200 172114 120000
rect 173438 119200 173494 120000
rect 174910 119200 174966 120000
rect 176382 119200 176438 120000
rect 177762 119200 177818 120000
rect 179234 119200 179290 120000
rect 846 0 902 800
rect 2502 0 2558 800
rect 4158 0 4214 800
rect 5814 0 5870 800
rect 7470 0 7526 800
rect 9126 0 9182 800
rect 10782 0 10838 800
rect 12438 0 12494 800
rect 14094 0 14150 800
rect 15842 0 15898 800
rect 17498 0 17554 800
rect 19154 0 19210 800
rect 20810 0 20866 800
rect 22466 0 22522 800
rect 24122 0 24178 800
rect 25778 0 25834 800
rect 27434 0 27490 800
rect 29182 0 29238 800
rect 30838 0 30894 800
rect 32494 0 32550 800
rect 34150 0 34206 800
rect 35806 0 35862 800
rect 37462 0 37518 800
rect 39118 0 39174 800
rect 40774 0 40830 800
rect 42522 0 42578 800
rect 44178 0 44234 800
rect 45834 0 45890 800
rect 47490 0 47546 800
rect 49146 0 49202 800
rect 50802 0 50858 800
rect 52458 0 52514 800
rect 54114 0 54170 800
rect 55770 0 55826 800
rect 57518 0 57574 800
rect 59174 0 59230 800
rect 60830 0 60886 800
rect 62486 0 62542 800
rect 64142 0 64198 800
rect 65798 0 65854 800
rect 67454 0 67510 800
rect 69110 0 69166 800
rect 70858 0 70914 800
rect 72514 0 72570 800
rect 74170 0 74226 800
rect 75826 0 75882 800
rect 77482 0 77538 800
rect 79138 0 79194 800
rect 80794 0 80850 800
rect 82450 0 82506 800
rect 84198 0 84254 800
rect 85854 0 85910 800
rect 87510 0 87566 800
rect 89166 0 89222 800
rect 90822 0 90878 800
rect 92478 0 92534 800
rect 94134 0 94190 800
rect 95790 0 95846 800
rect 97446 0 97502 800
rect 99194 0 99250 800
rect 100850 0 100906 800
rect 102506 0 102562 800
rect 104162 0 104218 800
rect 105818 0 105874 800
rect 107474 0 107530 800
rect 109130 0 109186 800
rect 110786 0 110842 800
rect 112534 0 112590 800
rect 114190 0 114246 800
rect 115846 0 115902 800
rect 117502 0 117558 800
rect 119158 0 119214 800
rect 120814 0 120870 800
rect 122470 0 122526 800
rect 124126 0 124182 800
rect 125874 0 125930 800
rect 127530 0 127586 800
rect 129186 0 129242 800
rect 130842 0 130898 800
rect 132498 0 132554 800
rect 134154 0 134210 800
rect 135810 0 135866 800
rect 137466 0 137522 800
rect 139122 0 139178 800
rect 140870 0 140926 800
rect 142526 0 142582 800
rect 144182 0 144238 800
rect 145838 0 145894 800
rect 147494 0 147550 800
rect 149150 0 149206 800
rect 150806 0 150862 800
rect 152462 0 152518 800
rect 154210 0 154266 800
rect 155866 0 155922 800
rect 157522 0 157578 800
rect 159178 0 159234 800
rect 160834 0 160890 800
rect 162490 0 162546 800
rect 164146 0 164202 800
rect 165802 0 165858 800
rect 167550 0 167606 800
rect 169206 0 169262 800
rect 170862 0 170918 800
rect 172518 0 172574 800
rect 174174 0 174230 800
rect 175830 0 175886 800
rect 177486 0 177542 800
rect 179142 0 179198 800
<< obsm2 >>
rect 774 119144 1986 119785
rect 2154 119144 3458 119785
rect 3626 119144 4838 119785
rect 5006 119144 6310 119785
rect 6478 119144 7782 119785
rect 7950 119144 9162 119785
rect 9330 119144 10634 119785
rect 10802 119144 12106 119785
rect 12274 119144 13486 119785
rect 13654 119144 14958 119785
rect 15126 119144 16430 119785
rect 16598 119144 17810 119785
rect 17978 119144 19282 119785
rect 19450 119144 20754 119785
rect 20922 119144 22134 119785
rect 22302 119144 23606 119785
rect 23774 119144 25078 119785
rect 25246 119144 26458 119785
rect 26626 119144 27930 119785
rect 28098 119144 29402 119785
rect 29570 119144 30782 119785
rect 30950 119144 32254 119785
rect 32422 119144 33726 119785
rect 33894 119144 35106 119785
rect 35274 119144 36578 119785
rect 36746 119144 38050 119785
rect 38218 119144 39430 119785
rect 39598 119144 40902 119785
rect 41070 119144 42374 119785
rect 42542 119144 43754 119785
rect 43922 119144 45226 119785
rect 45394 119144 46606 119785
rect 46774 119144 48078 119785
rect 48246 119144 49550 119785
rect 49718 119144 50930 119785
rect 51098 119144 52402 119785
rect 52570 119144 53874 119785
rect 54042 119144 55254 119785
rect 55422 119144 56726 119785
rect 56894 119144 58198 119785
rect 58366 119144 59578 119785
rect 59746 119144 61050 119785
rect 61218 119144 62522 119785
rect 62690 119144 63902 119785
rect 64070 119144 65374 119785
rect 65542 119144 66846 119785
rect 67014 119144 68226 119785
rect 68394 119144 69698 119785
rect 69866 119144 71170 119785
rect 71338 119144 72550 119785
rect 72718 119144 74022 119785
rect 74190 119144 75494 119785
rect 75662 119144 76874 119785
rect 77042 119144 78346 119785
rect 78514 119144 79818 119785
rect 79986 119144 81198 119785
rect 81366 119144 82670 119785
rect 82838 119144 84142 119785
rect 84310 119144 85522 119785
rect 85690 119144 86994 119785
rect 87162 119144 88466 119785
rect 88634 119144 89846 119785
rect 90014 119144 91318 119785
rect 91486 119144 92698 119785
rect 92866 119144 94170 119785
rect 94338 119144 95642 119785
rect 95810 119144 97022 119785
rect 97190 119144 98494 119785
rect 98662 119144 99966 119785
rect 100134 119144 101346 119785
rect 101514 119144 102818 119785
rect 102986 119144 104290 119785
rect 104458 119144 105670 119785
rect 105838 119144 107142 119785
rect 107310 119144 108614 119785
rect 108782 119144 109994 119785
rect 110162 119144 111466 119785
rect 111634 119144 112938 119785
rect 113106 119144 114318 119785
rect 114486 119144 115790 119785
rect 115958 119144 117262 119785
rect 117430 119144 118642 119785
rect 118810 119144 120114 119785
rect 120282 119144 121586 119785
rect 121754 119144 122966 119785
rect 123134 119144 124438 119785
rect 124606 119144 125910 119785
rect 126078 119144 127290 119785
rect 127458 119144 128762 119785
rect 128930 119144 130234 119785
rect 130402 119144 131614 119785
rect 131782 119144 133086 119785
rect 133254 119144 134558 119785
rect 134726 119144 135938 119785
rect 136106 119144 137410 119785
rect 137578 119144 138790 119785
rect 138958 119144 140262 119785
rect 140430 119144 141734 119785
rect 141902 119144 143114 119785
rect 143282 119144 144586 119785
rect 144754 119144 146058 119785
rect 146226 119144 147438 119785
rect 147606 119144 148910 119785
rect 149078 119144 150382 119785
rect 150550 119144 151762 119785
rect 151930 119144 153234 119785
rect 153402 119144 154706 119785
rect 154874 119144 156086 119785
rect 156254 119144 157558 119785
rect 157726 119144 159030 119785
rect 159198 119144 160410 119785
rect 160578 119144 161882 119785
rect 162050 119144 163354 119785
rect 163522 119144 164734 119785
rect 164902 119144 166206 119785
rect 166374 119144 167678 119785
rect 167846 119144 169058 119785
rect 169226 119144 170530 119785
rect 170698 119144 172002 119785
rect 172170 119144 173382 119785
rect 173550 119144 174854 119785
rect 175022 119144 176326 119785
rect 176494 119144 177706 119785
rect 177874 119144 179178 119785
rect 664 856 179288 119144
rect 664 167 790 856
rect 958 167 2446 856
rect 2614 167 4102 856
rect 4270 167 5758 856
rect 5926 167 7414 856
rect 7582 167 9070 856
rect 9238 167 10726 856
rect 10894 167 12382 856
rect 12550 167 14038 856
rect 14206 167 15786 856
rect 15954 167 17442 856
rect 17610 167 19098 856
rect 19266 167 20754 856
rect 20922 167 22410 856
rect 22578 167 24066 856
rect 24234 167 25722 856
rect 25890 167 27378 856
rect 27546 167 29126 856
rect 29294 167 30782 856
rect 30950 167 32438 856
rect 32606 167 34094 856
rect 34262 167 35750 856
rect 35918 167 37406 856
rect 37574 167 39062 856
rect 39230 167 40718 856
rect 40886 167 42466 856
rect 42634 167 44122 856
rect 44290 167 45778 856
rect 45946 167 47434 856
rect 47602 167 49090 856
rect 49258 167 50746 856
rect 50914 167 52402 856
rect 52570 167 54058 856
rect 54226 167 55714 856
rect 55882 167 57462 856
rect 57630 167 59118 856
rect 59286 167 60774 856
rect 60942 167 62430 856
rect 62598 167 64086 856
rect 64254 167 65742 856
rect 65910 167 67398 856
rect 67566 167 69054 856
rect 69222 167 70802 856
rect 70970 167 72458 856
rect 72626 167 74114 856
rect 74282 167 75770 856
rect 75938 167 77426 856
rect 77594 167 79082 856
rect 79250 167 80738 856
rect 80906 167 82394 856
rect 82562 167 84142 856
rect 84310 167 85798 856
rect 85966 167 87454 856
rect 87622 167 89110 856
rect 89278 167 90766 856
rect 90934 167 92422 856
rect 92590 167 94078 856
rect 94246 167 95734 856
rect 95902 167 97390 856
rect 97558 167 99138 856
rect 99306 167 100794 856
rect 100962 167 102450 856
rect 102618 167 104106 856
rect 104274 167 105762 856
rect 105930 167 107418 856
rect 107586 167 109074 856
rect 109242 167 110730 856
rect 110898 167 112478 856
rect 112646 167 114134 856
rect 114302 167 115790 856
rect 115958 167 117446 856
rect 117614 167 119102 856
rect 119270 167 120758 856
rect 120926 167 122414 856
rect 122582 167 124070 856
rect 124238 167 125818 856
rect 125986 167 127474 856
rect 127642 167 129130 856
rect 129298 167 130786 856
rect 130954 167 132442 856
rect 132610 167 134098 856
rect 134266 167 135754 856
rect 135922 167 137410 856
rect 137578 167 139066 856
rect 139234 167 140814 856
rect 140982 167 142470 856
rect 142638 167 144126 856
rect 144294 167 145782 856
rect 145950 167 147438 856
rect 147606 167 149094 856
rect 149262 167 150750 856
rect 150918 167 152406 856
rect 152574 167 154154 856
rect 154322 167 155810 856
rect 155978 167 157466 856
rect 157634 167 159122 856
rect 159290 167 160778 856
rect 160946 167 162434 856
rect 162602 167 164090 856
rect 164258 167 165746 856
rect 165914 167 167494 856
rect 167662 167 169150 856
rect 169318 167 170806 856
rect 170974 167 172462 856
rect 172630 167 174118 856
rect 174286 167 175774 856
rect 175942 167 177430 856
rect 177598 167 179086 856
rect 179254 167 179288 856
<< metal3 >>
rect 0 119688 800 119808
rect 0 119416 800 119536
rect 0 119144 800 119264
rect 0 118736 800 118856
rect 0 118464 800 118584
rect 0 118192 800 118312
rect 0 117784 800 117904
rect 0 117512 800 117632
rect 0 117240 800 117360
rect 0 116968 800 117088
rect 0 116560 800 116680
rect 0 116288 800 116408
rect 0 116016 800 116136
rect 0 115608 800 115728
rect 0 115336 800 115456
rect 0 115064 800 115184
rect 0 114656 800 114776
rect 0 114384 800 114504
rect 0 114112 800 114232
rect 0 113840 800 113960
rect 0 113432 800 113552
rect 0 113160 800 113280
rect 0 112888 800 113008
rect 0 112480 800 112600
rect 0 112208 800 112328
rect 0 111936 800 112056
rect 0 111528 800 111648
rect 0 111256 800 111376
rect 0 110984 800 111104
rect 0 110712 800 110832
rect 0 110304 800 110424
rect 0 110032 800 110152
rect 0 109760 800 109880
rect 0 109352 800 109472
rect 0 109080 800 109200
rect 0 108808 800 108928
rect 0 108536 800 108656
rect 0 108128 800 108248
rect 0 107856 800 107976
rect 0 107584 800 107704
rect 0 107176 800 107296
rect 0 106904 800 107024
rect 0 106632 800 106752
rect 0 106224 800 106344
rect 0 105952 800 106072
rect 0 105680 800 105800
rect 0 105408 800 105528
rect 0 105000 800 105120
rect 0 104728 800 104848
rect 0 104456 800 104576
rect 0 104048 800 104168
rect 0 103776 800 103896
rect 0 103504 800 103624
rect 0 103096 800 103216
rect 0 102824 800 102944
rect 0 102552 800 102672
rect 0 102280 800 102400
rect 0 101872 800 101992
rect 0 101600 800 101720
rect 0 101328 800 101448
rect 0 100920 800 101040
rect 0 100648 800 100768
rect 0 100376 800 100496
rect 0 100104 800 100224
rect 0 99696 800 99816
rect 0 99424 800 99544
rect 0 99152 800 99272
rect 0 98744 800 98864
rect 0 98472 800 98592
rect 0 98200 800 98320
rect 0 97792 800 97912
rect 0 97520 800 97640
rect 0 97248 800 97368
rect 0 96976 800 97096
rect 0 96568 800 96688
rect 0 96296 800 96416
rect 0 96024 800 96144
rect 0 95616 800 95736
rect 0 95344 800 95464
rect 0 95072 800 95192
rect 0 94664 800 94784
rect 0 94392 800 94512
rect 0 94120 800 94240
rect 0 93848 800 93968
rect 0 93440 800 93560
rect 0 93168 800 93288
rect 0 92896 800 93016
rect 0 92488 800 92608
rect 0 92216 800 92336
rect 0 91944 800 92064
rect 0 91536 800 91656
rect 0 91264 800 91384
rect 0 90992 800 91112
rect 0 90720 800 90840
rect 0 90312 800 90432
rect 0 90040 800 90160
rect 0 89768 800 89888
rect 0 89360 800 89480
rect 0 89088 800 89208
rect 0 88816 800 88936
rect 0 88544 800 88664
rect 0 88136 800 88256
rect 0 87864 800 87984
rect 0 87592 800 87712
rect 0 87184 800 87304
rect 0 86912 800 87032
rect 0 86640 800 86760
rect 0 86232 800 86352
rect 0 85960 800 86080
rect 0 85688 800 85808
rect 0 85416 800 85536
rect 0 85008 800 85128
rect 0 84736 800 84856
rect 0 84464 800 84584
rect 0 84056 800 84176
rect 0 83784 800 83904
rect 0 83512 800 83632
rect 0 83104 800 83224
rect 0 82832 800 82952
rect 0 82560 800 82680
rect 0 82288 800 82408
rect 0 81880 800 82000
rect 0 81608 800 81728
rect 0 81336 800 81456
rect 0 80928 800 81048
rect 0 80656 800 80776
rect 0 80384 800 80504
rect 0 80112 800 80232
rect 0 79704 800 79824
rect 0 79432 800 79552
rect 0 79160 800 79280
rect 0 78752 800 78872
rect 0 78480 800 78600
rect 0 78208 800 78328
rect 0 77800 800 77920
rect 0 77528 800 77648
rect 0 77256 800 77376
rect 0 76984 800 77104
rect 0 76576 800 76696
rect 0 76304 800 76424
rect 0 76032 800 76152
rect 0 75624 800 75744
rect 0 75352 800 75472
rect 0 75080 800 75200
rect 0 74672 800 74792
rect 0 74400 800 74520
rect 0 74128 800 74248
rect 0 73856 800 73976
rect 0 73448 800 73568
rect 0 73176 800 73296
rect 0 72904 800 73024
rect 0 72496 800 72616
rect 0 72224 800 72344
rect 0 71952 800 72072
rect 0 71544 800 71664
rect 0 71272 800 71392
rect 0 71000 800 71120
rect 0 70728 800 70848
rect 0 70320 800 70440
rect 0 70048 800 70168
rect 0 69776 800 69896
rect 0 69368 800 69488
rect 0 69096 800 69216
rect 0 68824 800 68944
rect 0 68552 800 68672
rect 0 68144 800 68264
rect 0 67872 800 67992
rect 0 67600 800 67720
rect 0 67192 800 67312
rect 0 66920 800 67040
rect 0 66648 800 66768
rect 0 66240 800 66360
rect 0 65968 800 66088
rect 0 65696 800 65816
rect 0 65424 800 65544
rect 0 65016 800 65136
rect 0 64744 800 64864
rect 0 64472 800 64592
rect 0 64064 800 64184
rect 0 63792 800 63912
rect 0 63520 800 63640
rect 0 63112 800 63232
rect 0 62840 800 62960
rect 0 62568 800 62688
rect 0 62296 800 62416
rect 0 61888 800 62008
rect 0 61616 800 61736
rect 0 61344 800 61464
rect 0 60936 800 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 179200 59984 180000 60104
rect 0 59712 800 59832
rect 0 59440 800 59560
rect 0 59168 800 59288
rect 0 58760 800 58880
rect 0 58488 800 58608
rect 0 58216 800 58336
rect 0 57808 800 57928
rect 0 57536 800 57656
rect 0 57264 800 57384
rect 0 56992 800 57112
rect 0 56584 800 56704
rect 0 56312 800 56432
rect 0 56040 800 56160
rect 0 55632 800 55752
rect 0 55360 800 55480
rect 0 55088 800 55208
rect 0 54680 800 54800
rect 0 54408 800 54528
rect 0 54136 800 54256
rect 0 53864 800 53984
rect 0 53456 800 53576
rect 0 53184 800 53304
rect 0 52912 800 53032
rect 0 52504 800 52624
rect 0 52232 800 52352
rect 0 51960 800 52080
rect 0 51552 800 51672
rect 0 51280 800 51400
rect 0 51008 800 51128
rect 0 50736 800 50856
rect 0 50328 800 50448
rect 0 50056 800 50176
rect 0 49784 800 49904
rect 0 49376 800 49496
rect 0 49104 800 49224
rect 0 48832 800 48952
rect 0 48560 800 48680
rect 0 48152 800 48272
rect 0 47880 800 48000
rect 0 47608 800 47728
rect 0 47200 800 47320
rect 0 46928 800 47048
rect 0 46656 800 46776
rect 0 46248 800 46368
rect 0 45976 800 46096
rect 0 45704 800 45824
rect 0 45432 800 45552
rect 0 45024 800 45144
rect 0 44752 800 44872
rect 0 44480 800 44600
rect 0 44072 800 44192
rect 0 43800 800 43920
rect 0 43528 800 43648
rect 0 43120 800 43240
rect 0 42848 800 42968
rect 0 42576 800 42696
rect 0 42304 800 42424
rect 0 41896 800 42016
rect 0 41624 800 41744
rect 0 41352 800 41472
rect 0 40944 800 41064
rect 0 40672 800 40792
rect 0 40400 800 40520
rect 0 40128 800 40248
rect 0 39720 800 39840
rect 0 39448 800 39568
rect 0 39176 800 39296
rect 0 38768 800 38888
rect 0 38496 800 38616
rect 0 38224 800 38344
rect 0 37816 800 37936
rect 0 37544 800 37664
rect 0 37272 800 37392
rect 0 37000 800 37120
rect 0 36592 800 36712
rect 0 36320 800 36440
rect 0 36048 800 36168
rect 0 35640 800 35760
rect 0 35368 800 35488
rect 0 35096 800 35216
rect 0 34688 800 34808
rect 0 34416 800 34536
rect 0 34144 800 34264
rect 0 33872 800 33992
rect 0 33464 800 33584
rect 0 33192 800 33312
rect 0 32920 800 33040
rect 0 32512 800 32632
rect 0 32240 800 32360
rect 0 31968 800 32088
rect 0 31560 800 31680
rect 0 31288 800 31408
rect 0 31016 800 31136
rect 0 30744 800 30864
rect 0 30336 800 30456
rect 0 30064 800 30184
rect 0 29792 800 29912
rect 0 29384 800 29504
rect 0 29112 800 29232
rect 0 28840 800 28960
rect 0 28568 800 28688
rect 0 28160 800 28280
rect 0 27888 800 28008
rect 0 27616 800 27736
rect 0 27208 800 27328
rect 0 26936 800 27056
rect 0 26664 800 26784
rect 0 26256 800 26376
rect 0 25984 800 26104
rect 0 25712 800 25832
rect 0 25440 800 25560
rect 0 25032 800 25152
rect 0 24760 800 24880
rect 0 24488 800 24608
rect 0 24080 800 24200
rect 0 23808 800 23928
rect 0 23536 800 23656
rect 0 23128 800 23248
rect 0 22856 800 22976
rect 0 22584 800 22704
rect 0 22312 800 22432
rect 0 21904 800 22024
rect 0 21632 800 21752
rect 0 21360 800 21480
rect 0 20952 800 21072
rect 0 20680 800 20800
rect 0 20408 800 20528
rect 0 20136 800 20256
rect 0 19728 800 19848
rect 0 19456 800 19576
rect 0 19184 800 19304
rect 0 18776 800 18896
rect 0 18504 800 18624
rect 0 18232 800 18352
rect 0 17824 800 17944
rect 0 17552 800 17672
rect 0 17280 800 17400
rect 0 17008 800 17128
rect 0 16600 800 16720
rect 0 16328 800 16448
rect 0 16056 800 16176
rect 0 15648 800 15768
rect 0 15376 800 15496
rect 0 15104 800 15224
rect 0 14696 800 14816
rect 0 14424 800 14544
rect 0 14152 800 14272
rect 0 13880 800 14000
rect 0 13472 800 13592
rect 0 13200 800 13320
rect 0 12928 800 13048
rect 0 12520 800 12640
rect 0 12248 800 12368
rect 0 11976 800 12096
rect 0 11568 800 11688
rect 0 11296 800 11416
rect 0 11024 800 11144
rect 0 10752 800 10872
rect 0 10344 800 10464
rect 0 10072 800 10192
rect 0 9800 800 9920
rect 0 9392 800 9512
rect 0 9120 800 9240
rect 0 8848 800 8968
rect 0 8576 800 8696
rect 0 8168 800 8288
rect 0 7896 800 8016
rect 0 7624 800 7744
rect 0 7216 800 7336
rect 0 6944 800 7064
rect 0 6672 800 6792
rect 0 6264 800 6384
rect 0 5992 800 6112
rect 0 5720 800 5840
rect 0 5448 800 5568
rect 0 5040 800 5160
rect 0 4768 800 4888
rect 0 4496 800 4616
rect 0 4088 800 4208
rect 0 3816 800 3936
rect 0 3544 800 3664
rect 0 3136 800 3256
rect 0 2864 800 2984
rect 0 2592 800 2712
rect 0 2320 800 2440
rect 0 1912 800 2032
rect 0 1640 800 1760
rect 0 1368 800 1488
rect 0 960 800 1080
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
<< obsm3 >>
rect 880 119064 179200 119781
rect 800 118936 179200 119064
rect 880 118112 179200 118936
rect 800 117984 179200 118112
rect 880 116888 179200 117984
rect 800 116760 179200 116888
rect 880 115936 179200 116760
rect 800 115808 179200 115936
rect 880 114984 179200 115808
rect 800 114856 179200 114984
rect 880 113760 179200 114856
rect 800 113632 179200 113760
rect 880 112808 179200 113632
rect 800 112680 179200 112808
rect 880 111856 179200 112680
rect 800 111728 179200 111856
rect 880 110632 179200 111728
rect 800 110504 179200 110632
rect 880 109680 179200 110504
rect 800 109552 179200 109680
rect 880 108456 179200 109552
rect 800 108328 179200 108456
rect 880 107504 179200 108328
rect 800 107376 179200 107504
rect 880 106552 179200 107376
rect 800 106424 179200 106552
rect 880 105328 179200 106424
rect 800 105200 179200 105328
rect 880 104376 179200 105200
rect 800 104248 179200 104376
rect 880 103424 179200 104248
rect 800 103296 179200 103424
rect 880 102200 179200 103296
rect 800 102072 179200 102200
rect 880 101248 179200 102072
rect 800 101120 179200 101248
rect 880 100024 179200 101120
rect 800 99896 179200 100024
rect 880 99072 179200 99896
rect 800 98944 179200 99072
rect 880 98120 179200 98944
rect 800 97992 179200 98120
rect 880 96896 179200 97992
rect 800 96768 179200 96896
rect 880 95944 179200 96768
rect 800 95816 179200 95944
rect 880 94992 179200 95816
rect 800 94864 179200 94992
rect 880 93768 179200 94864
rect 800 93640 179200 93768
rect 880 92816 179200 93640
rect 800 92688 179200 92816
rect 880 91864 179200 92688
rect 800 91736 179200 91864
rect 880 90640 179200 91736
rect 800 90512 179200 90640
rect 880 89688 179200 90512
rect 800 89560 179200 89688
rect 880 88464 179200 89560
rect 800 88336 179200 88464
rect 880 87512 179200 88336
rect 800 87384 179200 87512
rect 880 86560 179200 87384
rect 800 86432 179200 86560
rect 880 85336 179200 86432
rect 800 85208 179200 85336
rect 880 84384 179200 85208
rect 800 84256 179200 84384
rect 880 83432 179200 84256
rect 800 83304 179200 83432
rect 880 82208 179200 83304
rect 800 82080 179200 82208
rect 880 81256 179200 82080
rect 800 81128 179200 81256
rect 880 80032 179200 81128
rect 800 79904 179200 80032
rect 880 79080 179200 79904
rect 800 78952 179200 79080
rect 880 78128 179200 78952
rect 800 78000 179200 78128
rect 880 76904 179200 78000
rect 800 76776 179200 76904
rect 880 75952 179200 76776
rect 800 75824 179200 75952
rect 880 75000 179200 75824
rect 800 74872 179200 75000
rect 880 73776 179200 74872
rect 800 73648 179200 73776
rect 880 72824 179200 73648
rect 800 72696 179200 72824
rect 880 71872 179200 72696
rect 800 71744 179200 71872
rect 880 70648 179200 71744
rect 800 70520 179200 70648
rect 880 69696 179200 70520
rect 800 69568 179200 69696
rect 880 68472 179200 69568
rect 800 68344 179200 68472
rect 880 67520 179200 68344
rect 800 67392 179200 67520
rect 880 66568 179200 67392
rect 800 66440 179200 66568
rect 880 65344 179200 66440
rect 800 65216 179200 65344
rect 880 64392 179200 65216
rect 800 64264 179200 64392
rect 880 63440 179200 64264
rect 800 63312 179200 63440
rect 880 62216 179200 63312
rect 800 62088 179200 62216
rect 880 61264 179200 62088
rect 800 61136 179200 61264
rect 880 60184 179200 61136
rect 880 60040 179120 60184
rect 800 59912 179120 60040
rect 880 59904 179120 59912
rect 880 59088 179200 59904
rect 800 58960 179200 59088
rect 880 58136 179200 58960
rect 800 58008 179200 58136
rect 880 56912 179200 58008
rect 800 56784 179200 56912
rect 880 55960 179200 56784
rect 800 55832 179200 55960
rect 880 55008 179200 55832
rect 800 54880 179200 55008
rect 880 53784 179200 54880
rect 800 53656 179200 53784
rect 880 52832 179200 53656
rect 800 52704 179200 52832
rect 880 51880 179200 52704
rect 800 51752 179200 51880
rect 880 50656 179200 51752
rect 800 50528 179200 50656
rect 880 49704 179200 50528
rect 800 49576 179200 49704
rect 880 48480 179200 49576
rect 800 48352 179200 48480
rect 880 47528 179200 48352
rect 800 47400 179200 47528
rect 880 46576 179200 47400
rect 800 46448 179200 46576
rect 880 45352 179200 46448
rect 800 45224 179200 45352
rect 880 44400 179200 45224
rect 800 44272 179200 44400
rect 880 43448 179200 44272
rect 800 43320 179200 43448
rect 880 42224 179200 43320
rect 800 42096 179200 42224
rect 880 41272 179200 42096
rect 800 41144 179200 41272
rect 880 40048 179200 41144
rect 800 39920 179200 40048
rect 880 39096 179200 39920
rect 800 38968 179200 39096
rect 880 38144 179200 38968
rect 800 38016 179200 38144
rect 880 36920 179200 38016
rect 800 36792 179200 36920
rect 880 35968 179200 36792
rect 800 35840 179200 35968
rect 880 35016 179200 35840
rect 800 34888 179200 35016
rect 880 33792 179200 34888
rect 800 33664 179200 33792
rect 880 32840 179200 33664
rect 800 32712 179200 32840
rect 880 31888 179200 32712
rect 800 31760 179200 31888
rect 880 30664 179200 31760
rect 800 30536 179200 30664
rect 880 29712 179200 30536
rect 800 29584 179200 29712
rect 880 28488 179200 29584
rect 800 28360 179200 28488
rect 880 27536 179200 28360
rect 800 27408 179200 27536
rect 880 26584 179200 27408
rect 800 26456 179200 26584
rect 880 25360 179200 26456
rect 800 25232 179200 25360
rect 880 24408 179200 25232
rect 800 24280 179200 24408
rect 880 23456 179200 24280
rect 800 23328 179200 23456
rect 880 22232 179200 23328
rect 800 22104 179200 22232
rect 880 21280 179200 22104
rect 800 21152 179200 21280
rect 880 20056 179200 21152
rect 800 19928 179200 20056
rect 880 19104 179200 19928
rect 800 18976 179200 19104
rect 880 18152 179200 18976
rect 800 18024 179200 18152
rect 880 16928 179200 18024
rect 800 16800 179200 16928
rect 880 15976 179200 16800
rect 800 15848 179200 15976
rect 880 15024 179200 15848
rect 800 14896 179200 15024
rect 880 13800 179200 14896
rect 800 13672 179200 13800
rect 880 12848 179200 13672
rect 800 12720 179200 12848
rect 880 11896 179200 12720
rect 800 11768 179200 11896
rect 880 10672 179200 11768
rect 800 10544 179200 10672
rect 880 9720 179200 10544
rect 800 9592 179200 9720
rect 880 8496 179200 9592
rect 800 8368 179200 8496
rect 880 7544 179200 8368
rect 800 7416 179200 7544
rect 880 6592 179200 7416
rect 800 6464 179200 6592
rect 880 5368 179200 6464
rect 800 5240 179200 5368
rect 880 4416 179200 5240
rect 800 4288 179200 4416
rect 880 3464 179200 4288
rect 800 3336 179200 3464
rect 880 2240 179200 3336
rect 800 2112 179200 2240
rect 880 1288 179200 2112
rect 800 1160 179200 1288
rect 880 171 179200 1160
<< metal4 >>
rect 4208 2128 4528 117552
rect 4868 2176 5188 117504
rect 5528 2176 5848 117504
rect 6188 2176 6508 117504
rect 19568 2128 19888 117552
rect 20228 2176 20548 117504
rect 20888 2176 21208 117504
rect 21548 2176 21868 117504
rect 34928 2128 35248 117552
rect 35588 2176 35908 117504
rect 36248 2176 36568 117504
rect 36908 2176 37228 117504
rect 50288 2128 50608 117552
rect 50948 2176 51268 117504
rect 51608 2176 51928 117504
rect 52268 2176 52588 117504
rect 65648 2128 65968 117552
rect 66308 2176 66628 117504
rect 66968 2176 67288 117504
rect 67628 2176 67948 117504
rect 81008 2128 81328 117552
rect 81668 2176 81988 117504
rect 82328 2176 82648 117504
rect 82988 2176 83308 117504
rect 96368 2128 96688 117552
rect 97028 2176 97348 117504
rect 97688 2176 98008 117504
rect 98348 2176 98668 117504
rect 111728 2128 112048 117552
rect 112388 2176 112708 117504
rect 113048 2176 113368 117504
rect 113708 2176 114028 117504
rect 127088 2128 127408 117552
rect 127748 2176 128068 117504
rect 128408 2176 128728 117504
rect 129068 2176 129388 117504
rect 142448 2128 142768 117552
rect 143108 2176 143428 117504
rect 143768 2176 144088 117504
rect 144428 2176 144748 117504
rect 157808 2128 158128 117552
rect 158468 2176 158788 117504
rect 159128 2176 159448 117504
rect 159788 2176 160108 117504
rect 173168 2128 173488 117552
rect 173828 2176 174148 117504
rect 174488 2176 174808 117504
rect 175148 2176 175468 117504
<< labels >>
rlabel metal2 s 662 119200 718 120000 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 43810 119200 43866 120000 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 48134 119200 48190 120000 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 52458 119200 52514 120000 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 56782 119200 56838 120000 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 61106 119200 61162 120000 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 65430 119200 65486 120000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 69754 119200 69810 120000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 74078 119200 74134 120000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 78402 119200 78458 120000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 82726 119200 82782 120000 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 4894 119200 4950 120000 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 87050 119200 87106 120000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 91374 119200 91430 120000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 95698 119200 95754 120000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 100022 119200 100078 120000 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 104346 119200 104402 120000 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 108670 119200 108726 120000 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 112994 119200 113050 120000 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 117318 119200 117374 120000 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 121642 119200 121698 120000 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 125966 119200 126022 120000 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 9218 119200 9274 120000 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 130290 119200 130346 120000 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 134614 119200 134670 120000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 138846 119200 138902 120000 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 143170 119200 143226 120000 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 147494 119200 147550 120000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 151818 119200 151874 120000 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 156142 119200 156198 120000 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 160466 119200 160522 120000 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 13542 119200 13598 120000 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 17866 119200 17922 120000 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 22190 119200 22246 120000 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 26514 119200 26570 120000 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 30838 119200 30894 120000 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 35162 119200 35218 120000 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 39486 119200 39542 120000 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 2042 119200 2098 120000 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 45282 119200 45338 120000 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 49606 119200 49662 120000 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 53930 119200 53986 120000 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 58254 119200 58310 120000 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 62578 119200 62634 120000 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 66902 119200 66958 120000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 71226 119200 71282 120000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 75550 119200 75606 120000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 79874 119200 79930 120000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 84198 119200 84254 120000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 6366 119200 6422 120000 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 88522 119200 88578 120000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 92754 119200 92810 120000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 97078 119200 97134 120000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 101402 119200 101458 120000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 105726 119200 105782 120000 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 110050 119200 110106 120000 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 114374 119200 114430 120000 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 118698 119200 118754 120000 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 123022 119200 123078 120000 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 127346 119200 127402 120000 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 10690 119200 10746 120000 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 131670 119200 131726 120000 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 135994 119200 136050 120000 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 140318 119200 140374 120000 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 144642 119200 144698 120000 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 148966 119200 149022 120000 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 153290 119200 153346 120000 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 157614 119200 157670 120000 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 161938 119200 161994 120000 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 15014 119200 15070 120000 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 19338 119200 19394 120000 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 23662 119200 23718 120000 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 27986 119200 28042 120000 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 32310 119200 32366 120000 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 36634 119200 36690 120000 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 40958 119200 41014 120000 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 3514 119200 3570 120000 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 46662 119200 46718 120000 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 50986 119200 51042 120000 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 55310 119200 55366 120000 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 59634 119200 59690 120000 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 63958 119200 64014 120000 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 68282 119200 68338 120000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 72606 119200 72662 120000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 76930 119200 76986 120000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 81254 119200 81310 120000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 85578 119200 85634 120000 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 7838 119200 7894 120000 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 89902 119200 89958 120000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 94226 119200 94282 120000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 98550 119200 98606 120000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 102874 119200 102930 120000 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 107198 119200 107254 120000 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 111522 119200 111578 120000 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 115846 119200 115902 120000 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 120170 119200 120226 120000 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 124494 119200 124550 120000 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 128818 119200 128874 120000 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 12162 119200 12218 120000 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 133142 119200 133198 120000 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 137466 119200 137522 120000 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 141790 119200 141846 120000 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 146114 119200 146170 120000 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 150438 119200 150494 120000 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 154762 119200 154818 120000 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 159086 119200 159142 120000 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 163410 119200 163466 120000 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 16486 119200 16542 120000 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 20810 119200 20866 120000 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 25134 119200 25190 120000 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 29458 119200 29514 120000 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 33782 119200 33838 120000 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 38106 119200 38162 120000 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 42430 119200 42486 120000 6 io_out[9]
port 114 nsew signal output
rlabel metal3 s 179200 59984 180000 60104 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 177486 0 177542 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 179142 0 179198 800 6 irq[2]
port 117 nsew signal output
rlabel metal3 s 0 144 800 264 6 la_data_in[0]
port 118 nsew signal input
rlabel metal3 s 0 93848 800 93968 6 la_data_in[100]
port 119 nsew signal input
rlabel metal3 s 0 94664 800 94784 6 la_data_in[101]
port 120 nsew signal input
rlabel metal3 s 0 95616 800 95736 6 la_data_in[102]
port 121 nsew signal input
rlabel metal3 s 0 96568 800 96688 6 la_data_in[103]
port 122 nsew signal input
rlabel metal3 s 0 97520 800 97640 6 la_data_in[104]
port 123 nsew signal input
rlabel metal3 s 0 98472 800 98592 6 la_data_in[105]
port 124 nsew signal input
rlabel metal3 s 0 99424 800 99544 6 la_data_in[106]
port 125 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 la_data_in[107]
port 126 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 la_data_in[108]
port 127 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 la_data_in[109]
port 128 nsew signal input
rlabel metal3 s 0 9392 800 9512 6 la_data_in[10]
port 129 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 la_data_in[110]
port 130 nsew signal input
rlabel metal3 s 0 104048 800 104168 6 la_data_in[111]
port 131 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 la_data_in[112]
port 132 nsew signal input
rlabel metal3 s 0 105952 800 106072 6 la_data_in[113]
port 133 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 la_data_in[114]
port 134 nsew signal input
rlabel metal3 s 0 107856 800 107976 6 la_data_in[115]
port 135 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 la_data_in[116]
port 136 nsew signal input
rlabel metal3 s 0 109760 800 109880 6 la_data_in[117]
port 137 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 la_data_in[118]
port 138 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 la_data_in[119]
port 139 nsew signal input
rlabel metal3 s 0 10344 800 10464 6 la_data_in[11]
port 140 nsew signal input
rlabel metal3 s 0 112480 800 112600 6 la_data_in[120]
port 141 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 la_data_in[121]
port 142 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 la_data_in[122]
port 143 nsew signal input
rlabel metal3 s 0 115336 800 115456 6 la_data_in[123]
port 144 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 la_data_in[124]
port 145 nsew signal input
rlabel metal3 s 0 117240 800 117360 6 la_data_in[125]
port 146 nsew signal input
rlabel metal3 s 0 118192 800 118312 6 la_data_in[126]
port 147 nsew signal input
rlabel metal3 s 0 119144 800 119264 6 la_data_in[127]
port 148 nsew signal input
rlabel metal3 s 0 11296 800 11416 6 la_data_in[12]
port 149 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 la_data_in[13]
port 150 nsew signal input
rlabel metal3 s 0 13200 800 13320 6 la_data_in[14]
port 151 nsew signal input
rlabel metal3 s 0 14152 800 14272 6 la_data_in[15]
port 152 nsew signal input
rlabel metal3 s 0 15104 800 15224 6 la_data_in[16]
port 153 nsew signal input
rlabel metal3 s 0 16056 800 16176 6 la_data_in[17]
port 154 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 la_data_in[18]
port 155 nsew signal input
rlabel metal3 s 0 17824 800 17944 6 la_data_in[19]
port 156 nsew signal input
rlabel metal3 s 0 960 800 1080 6 la_data_in[1]
port 157 nsew signal input
rlabel metal3 s 0 18776 800 18896 6 la_data_in[20]
port 158 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 la_data_in[21]
port 159 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal3 s 0 21632 800 21752 6 la_data_in[23]
port 161 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 la_data_in[24]
port 162 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 la_data_in[25]
port 163 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 la_data_in[26]
port 164 nsew signal input
rlabel metal3 s 0 25440 800 25560 6 la_data_in[27]
port 165 nsew signal input
rlabel metal3 s 0 26256 800 26376 6 la_data_in[28]
port 166 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 la_data_in[29]
port 167 nsew signal input
rlabel metal3 s 0 1912 800 2032 6 la_data_in[2]
port 168 nsew signal input
rlabel metal3 s 0 28160 800 28280 6 la_data_in[30]
port 169 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 la_data_in[31]
port 170 nsew signal input
rlabel metal3 s 0 30064 800 30184 6 la_data_in[32]
port 171 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 la_data_in[33]
port 172 nsew signal input
rlabel metal3 s 0 31968 800 32088 6 la_data_in[34]
port 173 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 la_data_in[35]
port 174 nsew signal input
rlabel metal3 s 0 33872 800 33992 6 la_data_in[36]
port 175 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 la_data_in[37]
port 176 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 la_data_in[38]
port 177 nsew signal input
rlabel metal3 s 0 36592 800 36712 6 la_data_in[39]
port 178 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 la_data_in[3]
port 179 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 la_data_in[40]
port 180 nsew signal input
rlabel metal3 s 0 38496 800 38616 6 la_data_in[41]
port 181 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 la_data_in[42]
port 182 nsew signal input
rlabel metal3 s 0 40400 800 40520 6 la_data_in[43]
port 183 nsew signal input
rlabel metal3 s 0 41352 800 41472 6 la_data_in[44]
port 184 nsew signal input
rlabel metal3 s 0 42304 800 42424 6 la_data_in[45]
port 185 nsew signal input
rlabel metal3 s 0 43120 800 43240 6 la_data_in[46]
port 186 nsew signal input
rlabel metal3 s 0 44072 800 44192 6 la_data_in[47]
port 187 nsew signal input
rlabel metal3 s 0 45024 800 45144 6 la_data_in[48]
port 188 nsew signal input
rlabel metal3 s 0 45976 800 46096 6 la_data_in[49]
port 189 nsew signal input
rlabel metal3 s 0 3816 800 3936 6 la_data_in[4]
port 190 nsew signal input
rlabel metal3 s 0 46928 800 47048 6 la_data_in[50]
port 191 nsew signal input
rlabel metal3 s 0 47880 800 48000 6 la_data_in[51]
port 192 nsew signal input
rlabel metal3 s 0 48832 800 48952 6 la_data_in[52]
port 193 nsew signal input
rlabel metal3 s 0 49784 800 49904 6 la_data_in[53]
port 194 nsew signal input
rlabel metal3 s 0 50736 800 50856 6 la_data_in[54]
port 195 nsew signal input
rlabel metal3 s 0 51552 800 51672 6 la_data_in[55]
port 196 nsew signal input
rlabel metal3 s 0 52504 800 52624 6 la_data_in[56]
port 197 nsew signal input
rlabel metal3 s 0 53456 800 53576 6 la_data_in[57]
port 198 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 la_data_in[58]
port 199 nsew signal input
rlabel metal3 s 0 55360 800 55480 6 la_data_in[59]
port 200 nsew signal input
rlabel metal3 s 0 4768 800 4888 6 la_data_in[5]
port 201 nsew signal input
rlabel metal3 s 0 56312 800 56432 6 la_data_in[60]
port 202 nsew signal input
rlabel metal3 s 0 57264 800 57384 6 la_data_in[61]
port 203 nsew signal input
rlabel metal3 s 0 58216 800 58336 6 la_data_in[62]
port 204 nsew signal input
rlabel metal3 s 0 59168 800 59288 6 la_data_in[63]
port 205 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 la_data_in[64]
port 206 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 la_data_in[65]
port 207 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 la_data_in[66]
port 208 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 la_data_in[67]
port 209 nsew signal input
rlabel metal3 s 0 63792 800 63912 6 la_data_in[68]
port 210 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 la_data_in[69]
port 211 nsew signal input
rlabel metal3 s 0 5720 800 5840 6 la_data_in[6]
port 212 nsew signal input
rlabel metal3 s 0 65696 800 65816 6 la_data_in[70]
port 213 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 la_data_in[71]
port 214 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 la_data_in[72]
port 215 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 la_data_in[73]
port 216 nsew signal input
rlabel metal3 s 0 69368 800 69488 6 la_data_in[74]
port 217 nsew signal input
rlabel metal3 s 0 70320 800 70440 6 la_data_in[75]
port 218 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 la_data_in[76]
port 219 nsew signal input
rlabel metal3 s 0 72224 800 72344 6 la_data_in[77]
port 220 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 la_data_in[78]
port 221 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 la_data_in[79]
port 222 nsew signal input
rlabel metal3 s 0 6672 800 6792 6 la_data_in[7]
port 223 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 la_data_in[80]
port 224 nsew signal input
rlabel metal3 s 0 76032 800 76152 6 la_data_in[81]
port 225 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 la_data_in[82]
port 226 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 la_data_in[83]
port 227 nsew signal input
rlabel metal3 s 0 78752 800 78872 6 la_data_in[84]
port 228 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 la_data_in[85]
port 229 nsew signal input
rlabel metal3 s 0 80656 800 80776 6 la_data_in[86]
port 230 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 la_data_in[87]
port 231 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 la_data_in[88]
port 232 nsew signal input
rlabel metal3 s 0 83512 800 83632 6 la_data_in[89]
port 233 nsew signal input
rlabel metal3 s 0 7624 800 7744 6 la_data_in[8]
port 234 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 la_data_in[90]
port 235 nsew signal input
rlabel metal3 s 0 85416 800 85536 6 la_data_in[91]
port 236 nsew signal input
rlabel metal3 s 0 86232 800 86352 6 la_data_in[92]
port 237 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 la_data_in[93]
port 238 nsew signal input
rlabel metal3 s 0 88136 800 88256 6 la_data_in[94]
port 239 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 la_data_in[95]
port 240 nsew signal input
rlabel metal3 s 0 90040 800 90160 6 la_data_in[96]
port 241 nsew signal input
rlabel metal3 s 0 90992 800 91112 6 la_data_in[97]
port 242 nsew signal input
rlabel metal3 s 0 91944 800 92064 6 la_data_in[98]
port 243 nsew signal input
rlabel metal3 s 0 92896 800 93016 6 la_data_in[99]
port 244 nsew signal input
rlabel metal3 s 0 8576 800 8696 6 la_data_in[9]
port 245 nsew signal input
rlabel metal3 s 0 416 800 536 6 la_data_out[0]
port 246 nsew signal output
rlabel metal3 s 0 94120 800 94240 6 la_data_out[100]
port 247 nsew signal output
rlabel metal3 s 0 95072 800 95192 6 la_data_out[101]
port 248 nsew signal output
rlabel metal3 s 0 96024 800 96144 6 la_data_out[102]
port 249 nsew signal output
rlabel metal3 s 0 96976 800 97096 6 la_data_out[103]
port 250 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 la_data_out[104]
port 251 nsew signal output
rlabel metal3 s 0 98744 800 98864 6 la_data_out[105]
port 252 nsew signal output
rlabel metal3 s 0 99696 800 99816 6 la_data_out[106]
port 253 nsew signal output
rlabel metal3 s 0 100648 800 100768 6 la_data_out[107]
port 254 nsew signal output
rlabel metal3 s 0 101600 800 101720 6 la_data_out[108]
port 255 nsew signal output
rlabel metal3 s 0 102552 800 102672 6 la_data_out[109]
port 256 nsew signal output
rlabel metal3 s 0 9800 800 9920 6 la_data_out[10]
port 257 nsew signal output
rlabel metal3 s 0 103504 800 103624 6 la_data_out[110]
port 258 nsew signal output
rlabel metal3 s 0 104456 800 104576 6 la_data_out[111]
port 259 nsew signal output
rlabel metal3 s 0 105408 800 105528 6 la_data_out[112]
port 260 nsew signal output
rlabel metal3 s 0 106224 800 106344 6 la_data_out[113]
port 261 nsew signal output
rlabel metal3 s 0 107176 800 107296 6 la_data_out[114]
port 262 nsew signal output
rlabel metal3 s 0 108128 800 108248 6 la_data_out[115]
port 263 nsew signal output
rlabel metal3 s 0 109080 800 109200 6 la_data_out[116]
port 264 nsew signal output
rlabel metal3 s 0 110032 800 110152 6 la_data_out[117]
port 265 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 la_data_out[118]
port 266 nsew signal output
rlabel metal3 s 0 111936 800 112056 6 la_data_out[119]
port 267 nsew signal output
rlabel metal3 s 0 10752 800 10872 6 la_data_out[11]
port 268 nsew signal output
rlabel metal3 s 0 112888 800 113008 6 la_data_out[120]
port 269 nsew signal output
rlabel metal3 s 0 113840 800 113960 6 la_data_out[121]
port 270 nsew signal output
rlabel metal3 s 0 114656 800 114776 6 la_data_out[122]
port 271 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 la_data_out[123]
port 272 nsew signal output
rlabel metal3 s 0 116560 800 116680 6 la_data_out[124]
port 273 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 la_data_out[125]
port 274 nsew signal output
rlabel metal3 s 0 118464 800 118584 6 la_data_out[126]
port 275 nsew signal output
rlabel metal3 s 0 119416 800 119536 6 la_data_out[127]
port 276 nsew signal output
rlabel metal3 s 0 11568 800 11688 6 la_data_out[12]
port 277 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 la_data_out[13]
port 278 nsew signal output
rlabel metal3 s 0 13472 800 13592 6 la_data_out[14]
port 279 nsew signal output
rlabel metal3 s 0 14424 800 14544 6 la_data_out[15]
port 280 nsew signal output
rlabel metal3 s 0 15376 800 15496 6 la_data_out[16]
port 281 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 la_data_out[17]
port 282 nsew signal output
rlabel metal3 s 0 17280 800 17400 6 la_data_out[18]
port 283 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 la_data_out[19]
port 284 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 la_data_out[1]
port 285 nsew signal output
rlabel metal3 s 0 19184 800 19304 6 la_data_out[20]
port 286 nsew signal output
rlabel metal3 s 0 20136 800 20256 6 la_data_out[21]
port 287 nsew signal output
rlabel metal3 s 0 20952 800 21072 6 la_data_out[22]
port 288 nsew signal output
rlabel metal3 s 0 21904 800 22024 6 la_data_out[23]
port 289 nsew signal output
rlabel metal3 s 0 22856 800 22976 6 la_data_out[24]
port 290 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 la_data_out[25]
port 291 nsew signal output
rlabel metal3 s 0 24760 800 24880 6 la_data_out[26]
port 292 nsew signal output
rlabel metal3 s 0 25712 800 25832 6 la_data_out[27]
port 293 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 la_data_out[28]
port 294 nsew signal output
rlabel metal3 s 0 27616 800 27736 6 la_data_out[29]
port 295 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 la_data_out[2]
port 296 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 la_data_out[30]
port 297 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 la_data_out[31]
port 298 nsew signal output
rlabel metal3 s 0 30336 800 30456 6 la_data_out[32]
port 299 nsew signal output
rlabel metal3 s 0 31288 800 31408 6 la_data_out[33]
port 300 nsew signal output
rlabel metal3 s 0 32240 800 32360 6 la_data_out[34]
port 301 nsew signal output
rlabel metal3 s 0 33192 800 33312 6 la_data_out[35]
port 302 nsew signal output
rlabel metal3 s 0 34144 800 34264 6 la_data_out[36]
port 303 nsew signal output
rlabel metal3 s 0 35096 800 35216 6 la_data_out[37]
port 304 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 la_data_out[38]
port 305 nsew signal output
rlabel metal3 s 0 37000 800 37120 6 la_data_out[39]
port 306 nsew signal output
rlabel metal3 s 0 3136 800 3256 6 la_data_out[3]
port 307 nsew signal output
rlabel metal3 s 0 37816 800 37936 6 la_data_out[40]
port 308 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 la_data_out[41]
port 309 nsew signal output
rlabel metal3 s 0 39720 800 39840 6 la_data_out[42]
port 310 nsew signal output
rlabel metal3 s 0 40672 800 40792 6 la_data_out[43]
port 311 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 la_data_out[44]
port 312 nsew signal output
rlabel metal3 s 0 42576 800 42696 6 la_data_out[45]
port 313 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 la_data_out[46]
port 314 nsew signal output
rlabel metal3 s 0 44480 800 44600 6 la_data_out[47]
port 315 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 la_data_out[48]
port 316 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 la_data_out[49]
port 317 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 la_data_out[4]
port 318 nsew signal output
rlabel metal3 s 0 47200 800 47320 6 la_data_out[50]
port 319 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 la_data_out[51]
port 320 nsew signal output
rlabel metal3 s 0 49104 800 49224 6 la_data_out[52]
port 321 nsew signal output
rlabel metal3 s 0 50056 800 50176 6 la_data_out[53]
port 322 nsew signal output
rlabel metal3 s 0 51008 800 51128 6 la_data_out[54]
port 323 nsew signal output
rlabel metal3 s 0 51960 800 52080 6 la_data_out[55]
port 324 nsew signal output
rlabel metal3 s 0 52912 800 53032 6 la_data_out[56]
port 325 nsew signal output
rlabel metal3 s 0 53864 800 53984 6 la_data_out[57]
port 326 nsew signal output
rlabel metal3 s 0 54680 800 54800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal3 s 0 55632 800 55752 6 la_data_out[59]
port 328 nsew signal output
rlabel metal3 s 0 5040 800 5160 6 la_data_out[5]
port 329 nsew signal output
rlabel metal3 s 0 56584 800 56704 6 la_data_out[60]
port 330 nsew signal output
rlabel metal3 s 0 57536 800 57656 6 la_data_out[61]
port 331 nsew signal output
rlabel metal3 s 0 58488 800 58608 6 la_data_out[62]
port 332 nsew signal output
rlabel metal3 s 0 59440 800 59560 6 la_data_out[63]
port 333 nsew signal output
rlabel metal3 s 0 60392 800 60512 6 la_data_out[64]
port 334 nsew signal output
rlabel metal3 s 0 61344 800 61464 6 la_data_out[65]
port 335 nsew signal output
rlabel metal3 s 0 62296 800 62416 6 la_data_out[66]
port 336 nsew signal output
rlabel metal3 s 0 63112 800 63232 6 la_data_out[67]
port 337 nsew signal output
rlabel metal3 s 0 64064 800 64184 6 la_data_out[68]
port 338 nsew signal output
rlabel metal3 s 0 65016 800 65136 6 la_data_out[69]
port 339 nsew signal output
rlabel metal3 s 0 5992 800 6112 6 la_data_out[6]
port 340 nsew signal output
rlabel metal3 s 0 65968 800 66088 6 la_data_out[70]
port 341 nsew signal output
rlabel metal3 s 0 66920 800 67040 6 la_data_out[71]
port 342 nsew signal output
rlabel metal3 s 0 67872 800 67992 6 la_data_out[72]
port 343 nsew signal output
rlabel metal3 s 0 68824 800 68944 6 la_data_out[73]
port 344 nsew signal output
rlabel metal3 s 0 69776 800 69896 6 la_data_out[74]
port 345 nsew signal output
rlabel metal3 s 0 70728 800 70848 6 la_data_out[75]
port 346 nsew signal output
rlabel metal3 s 0 71544 800 71664 6 la_data_out[76]
port 347 nsew signal output
rlabel metal3 s 0 72496 800 72616 6 la_data_out[77]
port 348 nsew signal output
rlabel metal3 s 0 73448 800 73568 6 la_data_out[78]
port 349 nsew signal output
rlabel metal3 s 0 74400 800 74520 6 la_data_out[79]
port 350 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 la_data_out[7]
port 351 nsew signal output
rlabel metal3 s 0 75352 800 75472 6 la_data_out[80]
port 352 nsew signal output
rlabel metal3 s 0 76304 800 76424 6 la_data_out[81]
port 353 nsew signal output
rlabel metal3 s 0 77256 800 77376 6 la_data_out[82]
port 354 nsew signal output
rlabel metal3 s 0 78208 800 78328 6 la_data_out[83]
port 355 nsew signal output
rlabel metal3 s 0 79160 800 79280 6 la_data_out[84]
port 356 nsew signal output
rlabel metal3 s 0 80112 800 80232 6 la_data_out[85]
port 357 nsew signal output
rlabel metal3 s 0 80928 800 81048 6 la_data_out[86]
port 358 nsew signal output
rlabel metal3 s 0 81880 800 82000 6 la_data_out[87]
port 359 nsew signal output
rlabel metal3 s 0 82832 800 82952 6 la_data_out[88]
port 360 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 la_data_out[89]
port 361 nsew signal output
rlabel metal3 s 0 7896 800 8016 6 la_data_out[8]
port 362 nsew signal output
rlabel metal3 s 0 84736 800 84856 6 la_data_out[90]
port 363 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 la_data_out[91]
port 364 nsew signal output
rlabel metal3 s 0 86640 800 86760 6 la_data_out[92]
port 365 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 la_data_out[93]
port 366 nsew signal output
rlabel metal3 s 0 88544 800 88664 6 la_data_out[94]
port 367 nsew signal output
rlabel metal3 s 0 89360 800 89480 6 la_data_out[95]
port 368 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 la_data_out[96]
port 369 nsew signal output
rlabel metal3 s 0 91264 800 91384 6 la_data_out[97]
port 370 nsew signal output
rlabel metal3 s 0 92216 800 92336 6 la_data_out[98]
port 371 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 la_data_out[99]
port 372 nsew signal output
rlabel metal3 s 0 8848 800 8968 6 la_data_out[9]
port 373 nsew signal output
rlabel metal3 s 0 688 800 808 6 la_oenb[0]
port 374 nsew signal input
rlabel metal3 s 0 94392 800 94512 6 la_oenb[100]
port 375 nsew signal input
rlabel metal3 s 0 95344 800 95464 6 la_oenb[101]
port 376 nsew signal input
rlabel metal3 s 0 96296 800 96416 6 la_oenb[102]
port 377 nsew signal input
rlabel metal3 s 0 97248 800 97368 6 la_oenb[103]
port 378 nsew signal input
rlabel metal3 s 0 98200 800 98320 6 la_oenb[104]
port 379 nsew signal input
rlabel metal3 s 0 99152 800 99272 6 la_oenb[105]
port 380 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 la_oenb[106]
port 381 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 la_oenb[107]
port 382 nsew signal input
rlabel metal3 s 0 101872 800 101992 6 la_oenb[108]
port 383 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 la_oenb[109]
port 384 nsew signal input
rlabel metal3 s 0 10072 800 10192 6 la_oenb[10]
port 385 nsew signal input
rlabel metal3 s 0 103776 800 103896 6 la_oenb[110]
port 386 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 la_oenb[111]
port 387 nsew signal input
rlabel metal3 s 0 105680 800 105800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 la_oenb[113]
port 389 nsew signal input
rlabel metal3 s 0 107584 800 107704 6 la_oenb[114]
port 390 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 la_oenb[115]
port 391 nsew signal input
rlabel metal3 s 0 109352 800 109472 6 la_oenb[116]
port 392 nsew signal input
rlabel metal3 s 0 110304 800 110424 6 la_oenb[117]
port 393 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 la_oenb[118]
port 394 nsew signal input
rlabel metal3 s 0 112208 800 112328 6 la_oenb[119]
port 395 nsew signal input
rlabel metal3 s 0 11024 800 11144 6 la_oenb[11]
port 396 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 la_oenb[120]
port 397 nsew signal input
rlabel metal3 s 0 114112 800 114232 6 la_oenb[121]
port 398 nsew signal input
rlabel metal3 s 0 115064 800 115184 6 la_oenb[122]
port 399 nsew signal input
rlabel metal3 s 0 116016 800 116136 6 la_oenb[123]
port 400 nsew signal input
rlabel metal3 s 0 116968 800 117088 6 la_oenb[124]
port 401 nsew signal input
rlabel metal3 s 0 117784 800 117904 6 la_oenb[125]
port 402 nsew signal input
rlabel metal3 s 0 118736 800 118856 6 la_oenb[126]
port 403 nsew signal input
rlabel metal3 s 0 119688 800 119808 6 la_oenb[127]
port 404 nsew signal input
rlabel metal3 s 0 11976 800 12096 6 la_oenb[12]
port 405 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 la_oenb[13]
port 406 nsew signal input
rlabel metal3 s 0 13880 800 14000 6 la_oenb[14]
port 407 nsew signal input
rlabel metal3 s 0 14696 800 14816 6 la_oenb[15]
port 408 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 la_oenb[16]
port 409 nsew signal input
rlabel metal3 s 0 16600 800 16720 6 la_oenb[17]
port 410 nsew signal input
rlabel metal3 s 0 17552 800 17672 6 la_oenb[18]
port 411 nsew signal input
rlabel metal3 s 0 18504 800 18624 6 la_oenb[19]
port 412 nsew signal input
rlabel metal3 s 0 1640 800 1760 6 la_oenb[1]
port 413 nsew signal input
rlabel metal3 s 0 19456 800 19576 6 la_oenb[20]
port 414 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 la_oenb[21]
port 415 nsew signal input
rlabel metal3 s 0 21360 800 21480 6 la_oenb[22]
port 416 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 la_oenb[23]
port 417 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 la_oenb[24]
port 418 nsew signal input
rlabel metal3 s 0 24080 800 24200 6 la_oenb[25]
port 419 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 la_oenb[26]
port 420 nsew signal input
rlabel metal3 s 0 25984 800 26104 6 la_oenb[27]
port 421 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 la_oenb[28]
port 422 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 la_oenb[29]
port 423 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 la_oenb[2]
port 424 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 la_oenb[30]
port 425 nsew signal input
rlabel metal3 s 0 29792 800 29912 6 la_oenb[31]
port 426 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 la_oenb[32]
port 427 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 la_oenb[33]
port 428 nsew signal input
rlabel metal3 s 0 32512 800 32632 6 la_oenb[34]
port 429 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 la_oenb[35]
port 430 nsew signal input
rlabel metal3 s 0 34416 800 34536 6 la_oenb[36]
port 431 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 la_oenb[37]
port 432 nsew signal input
rlabel metal3 s 0 36320 800 36440 6 la_oenb[38]
port 433 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 la_oenb[39]
port 434 nsew signal input
rlabel metal3 s 0 3544 800 3664 6 la_oenb[3]
port 435 nsew signal input
rlabel metal3 s 0 38224 800 38344 6 la_oenb[40]
port 436 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 la_oenb[41]
port 437 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 la_oenb[42]
port 438 nsew signal input
rlabel metal3 s 0 40944 800 41064 6 la_oenb[43]
port 439 nsew signal input
rlabel metal3 s 0 41896 800 42016 6 la_oenb[44]
port 440 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 la_oenb[45]
port 441 nsew signal input
rlabel metal3 s 0 43800 800 43920 6 la_oenb[46]
port 442 nsew signal input
rlabel metal3 s 0 44752 800 44872 6 la_oenb[47]
port 443 nsew signal input
rlabel metal3 s 0 45704 800 45824 6 la_oenb[48]
port 444 nsew signal input
rlabel metal3 s 0 46656 800 46776 6 la_oenb[49]
port 445 nsew signal input
rlabel metal3 s 0 4496 800 4616 6 la_oenb[4]
port 446 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 la_oenb[50]
port 447 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 la_oenb[51]
port 448 nsew signal input
rlabel metal3 s 0 49376 800 49496 6 la_oenb[52]
port 449 nsew signal input
rlabel metal3 s 0 50328 800 50448 6 la_oenb[53]
port 450 nsew signal input
rlabel metal3 s 0 51280 800 51400 6 la_oenb[54]
port 451 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 la_oenb[55]
port 452 nsew signal input
rlabel metal3 s 0 53184 800 53304 6 la_oenb[56]
port 453 nsew signal input
rlabel metal3 s 0 54136 800 54256 6 la_oenb[57]
port 454 nsew signal input
rlabel metal3 s 0 55088 800 55208 6 la_oenb[58]
port 455 nsew signal input
rlabel metal3 s 0 56040 800 56160 6 la_oenb[59]
port 456 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 la_oenb[5]
port 457 nsew signal input
rlabel metal3 s 0 56992 800 57112 6 la_oenb[60]
port 458 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 la_oenb[61]
port 459 nsew signal input
rlabel metal3 s 0 58760 800 58880 6 la_oenb[62]
port 460 nsew signal input
rlabel metal3 s 0 59712 800 59832 6 la_oenb[63]
port 461 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 la_oenb[64]
port 462 nsew signal input
rlabel metal3 s 0 61616 800 61736 6 la_oenb[65]
port 463 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 la_oenb[66]
port 464 nsew signal input
rlabel metal3 s 0 63520 800 63640 6 la_oenb[67]
port 465 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 la_oenb[68]
port 466 nsew signal input
rlabel metal3 s 0 65424 800 65544 6 la_oenb[69]
port 467 nsew signal input
rlabel metal3 s 0 6264 800 6384 6 la_oenb[6]
port 468 nsew signal input
rlabel metal3 s 0 66240 800 66360 6 la_oenb[70]
port 469 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 la_oenb[71]
port 470 nsew signal input
rlabel metal3 s 0 68144 800 68264 6 la_oenb[72]
port 471 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 la_oenb[73]
port 472 nsew signal input
rlabel metal3 s 0 70048 800 70168 6 la_oenb[74]
port 473 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 la_oenb[75]
port 474 nsew signal input
rlabel metal3 s 0 71952 800 72072 6 la_oenb[76]
port 475 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 la_oenb[77]
port 476 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 la_oenb[78]
port 477 nsew signal input
rlabel metal3 s 0 74672 800 74792 6 la_oenb[79]
port 478 nsew signal input
rlabel metal3 s 0 7216 800 7336 6 la_oenb[7]
port 479 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 la_oenb[80]
port 480 nsew signal input
rlabel metal3 s 0 76576 800 76696 6 la_oenb[81]
port 481 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 la_oenb[82]
port 482 nsew signal input
rlabel metal3 s 0 78480 800 78600 6 la_oenb[83]
port 483 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 la_oenb[84]
port 484 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 la_oenb[85]
port 485 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 la_oenb[86]
port 486 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 la_oenb[87]
port 487 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 la_oenb[88]
port 488 nsew signal input
rlabel metal3 s 0 84056 800 84176 6 la_oenb[89]
port 489 nsew signal input
rlabel metal3 s 0 8168 800 8288 6 la_oenb[8]
port 490 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 la_oenb[90]
port 491 nsew signal input
rlabel metal3 s 0 85960 800 86080 6 la_oenb[91]
port 492 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 la_oenb[92]
port 493 nsew signal input
rlabel metal3 s 0 87864 800 87984 6 la_oenb[93]
port 494 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 la_oenb[94]
port 495 nsew signal input
rlabel metal3 s 0 89768 800 89888 6 la_oenb[95]
port 496 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 la_oenb[96]
port 497 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 la_oenb[97]
port 498 nsew signal input
rlabel metal3 s 0 92488 800 92608 6 la_oenb[98]
port 499 nsew signal input
rlabel metal3 s 0 93440 800 93560 6 la_oenb[99]
port 500 nsew signal input
rlabel metal3 s 0 9120 800 9240 6 la_oenb[9]
port 501 nsew signal input
rlabel metal2 s 164790 119200 164846 120000 6 phase_in[0]
port 502 nsew signal input
rlabel metal2 s 179234 119200 179290 120000 6 phase_in[10]
port 503 nsew signal input
rlabel metal2 s 166262 119200 166318 120000 6 phase_in[1]
port 504 nsew signal input
rlabel metal2 s 167734 119200 167790 120000 6 phase_in[2]
port 505 nsew signal input
rlabel metal2 s 169114 119200 169170 120000 6 phase_in[3]
port 506 nsew signal input
rlabel metal2 s 170586 119200 170642 120000 6 phase_in[4]
port 507 nsew signal input
rlabel metal2 s 172058 119200 172114 120000 6 phase_in[5]
port 508 nsew signal input
rlabel metal2 s 173438 119200 173494 120000 6 phase_in[6]
port 509 nsew signal input
rlabel metal2 s 174910 119200 174966 120000 6 phase_in[7]
port 510 nsew signal input
rlabel metal2 s 176382 119200 176438 120000 6 phase_in[8]
port 511 nsew signal input
rlabel metal2 s 177762 119200 177818 120000 6 phase_in[9]
port 512 nsew signal input
rlabel metal2 s 846 0 902 800 6 wb_clk_i
port 513 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wb_rst_i
port 514 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_ack_o
port 515 nsew signal output
rlabel metal2 s 10782 0 10838 800 6 wbs_adr_i[0]
port 516 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 wbs_adr_i[10]
port 517 nsew signal input
rlabel metal2 s 72514 0 72570 800 6 wbs_adr_i[11]
port 518 nsew signal input
rlabel metal2 s 77482 0 77538 800 6 wbs_adr_i[12]
port 519 nsew signal input
rlabel metal2 s 82450 0 82506 800 6 wbs_adr_i[13]
port 520 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 wbs_adr_i[14]
port 521 nsew signal input
rlabel metal2 s 92478 0 92534 800 6 wbs_adr_i[15]
port 522 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 wbs_adr_i[16]
port 523 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 wbs_adr_i[17]
port 524 nsew signal input
rlabel metal2 s 107474 0 107530 800 6 wbs_adr_i[18]
port 525 nsew signal input
rlabel metal2 s 112534 0 112590 800 6 wbs_adr_i[19]
port 526 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 wbs_adr_i[1]
port 527 nsew signal input
rlabel metal2 s 117502 0 117558 800 6 wbs_adr_i[20]
port 528 nsew signal input
rlabel metal2 s 122470 0 122526 800 6 wbs_adr_i[21]
port 529 nsew signal input
rlabel metal2 s 127530 0 127586 800 6 wbs_adr_i[22]
port 530 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 wbs_adr_i[23]
port 531 nsew signal input
rlabel metal2 s 137466 0 137522 800 6 wbs_adr_i[24]
port 532 nsew signal input
rlabel metal2 s 142526 0 142582 800 6 wbs_adr_i[25]
port 533 nsew signal input
rlabel metal2 s 147494 0 147550 800 6 wbs_adr_i[26]
port 534 nsew signal input
rlabel metal2 s 152462 0 152518 800 6 wbs_adr_i[27]
port 535 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 wbs_adr_i[28]
port 536 nsew signal input
rlabel metal2 s 162490 0 162546 800 6 wbs_adr_i[29]
port 537 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 wbs_adr_i[2]
port 538 nsew signal input
rlabel metal2 s 167550 0 167606 800 6 wbs_adr_i[30]
port 539 nsew signal input
rlabel metal2 s 172518 0 172574 800 6 wbs_adr_i[31]
port 540 nsew signal input
rlabel metal2 s 30838 0 30894 800 6 wbs_adr_i[3]
port 541 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 wbs_adr_i[4]
port 542 nsew signal input
rlabel metal2 s 42522 0 42578 800 6 wbs_adr_i[5]
port 543 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_adr_i[6]
port 544 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 wbs_adr_i[7]
port 545 nsew signal input
rlabel metal2 s 57518 0 57574 800 6 wbs_adr_i[8]
port 546 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 wbs_adr_i[9]
port 547 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 wbs_cyc_i
port 548 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_i[0]
port 549 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 wbs_dat_i[10]
port 550 nsew signal input
rlabel metal2 s 74170 0 74226 800 6 wbs_dat_i[11]
port 551 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 wbs_dat_i[12]
port 552 nsew signal input
rlabel metal2 s 84198 0 84254 800 6 wbs_dat_i[13]
port 553 nsew signal input
rlabel metal2 s 89166 0 89222 800 6 wbs_dat_i[14]
port 554 nsew signal input
rlabel metal2 s 94134 0 94190 800 6 wbs_dat_i[15]
port 555 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 wbs_dat_i[16]
port 556 nsew signal input
rlabel metal2 s 104162 0 104218 800 6 wbs_dat_i[17]
port 557 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 wbs_dat_i[18]
port 558 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 wbs_dat_i[19]
port 559 nsew signal input
rlabel metal2 s 19154 0 19210 800 6 wbs_dat_i[1]
port 560 nsew signal input
rlabel metal2 s 119158 0 119214 800 6 wbs_dat_i[20]
port 561 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 wbs_dat_i[21]
port 562 nsew signal input
rlabel metal2 s 129186 0 129242 800 6 wbs_dat_i[22]
port 563 nsew signal input
rlabel metal2 s 134154 0 134210 800 6 wbs_dat_i[23]
port 564 nsew signal input
rlabel metal2 s 139122 0 139178 800 6 wbs_dat_i[24]
port 565 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 wbs_dat_i[25]
port 566 nsew signal input
rlabel metal2 s 149150 0 149206 800 6 wbs_dat_i[26]
port 567 nsew signal input
rlabel metal2 s 154210 0 154266 800 6 wbs_dat_i[27]
port 568 nsew signal input
rlabel metal2 s 159178 0 159234 800 6 wbs_dat_i[28]
port 569 nsew signal input
rlabel metal2 s 164146 0 164202 800 6 wbs_dat_i[29]
port 570 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 wbs_dat_i[2]
port 571 nsew signal input
rlabel metal2 s 169206 0 169262 800 6 wbs_dat_i[30]
port 572 nsew signal input
rlabel metal2 s 174174 0 174230 800 6 wbs_dat_i[31]
port 573 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 wbs_dat_i[3]
port 574 nsew signal input
rlabel metal2 s 39118 0 39174 800 6 wbs_dat_i[4]
port 575 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 wbs_dat_i[5]
port 576 nsew signal input
rlabel metal2 s 49146 0 49202 800 6 wbs_dat_i[6]
port 577 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 wbs_dat_i[7]
port 578 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 wbs_dat_i[8]
port 579 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 wbs_dat_i[9]
port 580 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 wbs_dat_o[0]
port 581 nsew signal output
rlabel metal2 s 70858 0 70914 800 6 wbs_dat_o[10]
port 582 nsew signal output
rlabel metal2 s 75826 0 75882 800 6 wbs_dat_o[11]
port 583 nsew signal output
rlabel metal2 s 80794 0 80850 800 6 wbs_dat_o[12]
port 584 nsew signal output
rlabel metal2 s 85854 0 85910 800 6 wbs_dat_o[13]
port 585 nsew signal output
rlabel metal2 s 90822 0 90878 800 6 wbs_dat_o[14]
port 586 nsew signal output
rlabel metal2 s 95790 0 95846 800 6 wbs_dat_o[15]
port 587 nsew signal output
rlabel metal2 s 100850 0 100906 800 6 wbs_dat_o[16]
port 588 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 wbs_dat_o[17]
port 589 nsew signal output
rlabel metal2 s 110786 0 110842 800 6 wbs_dat_o[18]
port 590 nsew signal output
rlabel metal2 s 115846 0 115902 800 6 wbs_dat_o[19]
port 591 nsew signal output
rlabel metal2 s 20810 0 20866 800 6 wbs_dat_o[1]
port 592 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 wbs_dat_o[20]
port 593 nsew signal output
rlabel metal2 s 125874 0 125930 800 6 wbs_dat_o[21]
port 594 nsew signal output
rlabel metal2 s 130842 0 130898 800 6 wbs_dat_o[22]
port 595 nsew signal output
rlabel metal2 s 135810 0 135866 800 6 wbs_dat_o[23]
port 596 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 wbs_dat_o[24]
port 597 nsew signal output
rlabel metal2 s 145838 0 145894 800 6 wbs_dat_o[25]
port 598 nsew signal output
rlabel metal2 s 150806 0 150862 800 6 wbs_dat_o[26]
port 599 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 wbs_dat_o[27]
port 600 nsew signal output
rlabel metal2 s 160834 0 160890 800 6 wbs_dat_o[28]
port 601 nsew signal output
rlabel metal2 s 165802 0 165858 800 6 wbs_dat_o[29]
port 602 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 wbs_dat_o[2]
port 603 nsew signal output
rlabel metal2 s 170862 0 170918 800 6 wbs_dat_o[30]
port 604 nsew signal output
rlabel metal2 s 175830 0 175886 800 6 wbs_dat_o[31]
port 605 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 wbs_dat_o[3]
port 606 nsew signal output
rlabel metal2 s 40774 0 40830 800 6 wbs_dat_o[4]
port 607 nsew signal output
rlabel metal2 s 45834 0 45890 800 6 wbs_dat_o[5]
port 608 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 wbs_dat_o[6]
port 609 nsew signal output
rlabel metal2 s 55770 0 55826 800 6 wbs_dat_o[7]
port 610 nsew signal output
rlabel metal2 s 60830 0 60886 800 6 wbs_dat_o[8]
port 611 nsew signal output
rlabel metal2 s 65798 0 65854 800 6 wbs_dat_o[9]
port 612 nsew signal output
rlabel metal2 s 15842 0 15898 800 6 wbs_sel_i[0]
port 613 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 wbs_sel_i[1]
port 614 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 wbs_sel_i[2]
port 615 nsew signal input
rlabel metal2 s 35806 0 35862 800 6 wbs_sel_i[3]
port 616 nsew signal input
rlabel metal2 s 7470 0 7526 800 6 wbs_stb_i
port 617 nsew signal input
rlabel metal2 s 9126 0 9182 800 6 wbs_we_i
port 618 nsew signal input
rlabel metal4 s 157808 2128 158128 117552 6 vccd1
port 619 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 117552 6 vccd1
port 620 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 117552 6 vccd1
port 621 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 117552 6 vccd1
port 622 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 117552 6 vccd1
port 623 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 117552 6 vccd1
port 624 nsew power bidirectional
rlabel metal4 s 173168 2128 173488 117552 6 vssd1
port 625 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 117552 6 vssd1
port 626 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 117552 6 vssd1
port 627 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 117552 6 vssd1
port 628 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 117552 6 vssd1
port 629 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 117552 6 vssd1
port 630 nsew ground bidirectional
rlabel metal4 s 158468 2176 158788 117504 6 vccd2
port 631 nsew power bidirectional
rlabel metal4 s 127748 2176 128068 117504 6 vccd2
port 632 nsew power bidirectional
rlabel metal4 s 97028 2176 97348 117504 6 vccd2
port 633 nsew power bidirectional
rlabel metal4 s 66308 2176 66628 117504 6 vccd2
port 634 nsew power bidirectional
rlabel metal4 s 35588 2176 35908 117504 6 vccd2
port 635 nsew power bidirectional
rlabel metal4 s 4868 2176 5188 117504 6 vccd2
port 636 nsew power bidirectional
rlabel metal4 s 173828 2176 174148 117504 6 vssd2
port 637 nsew ground bidirectional
rlabel metal4 s 143108 2176 143428 117504 6 vssd2
port 638 nsew ground bidirectional
rlabel metal4 s 112388 2176 112708 117504 6 vssd2
port 639 nsew ground bidirectional
rlabel metal4 s 81668 2176 81988 117504 6 vssd2
port 640 nsew ground bidirectional
rlabel metal4 s 50948 2176 51268 117504 6 vssd2
port 641 nsew ground bidirectional
rlabel metal4 s 20228 2176 20548 117504 6 vssd2
port 642 nsew ground bidirectional
rlabel metal4 s 159128 2176 159448 117504 6 vdda1
port 643 nsew power bidirectional
rlabel metal4 s 128408 2176 128728 117504 6 vdda1
port 644 nsew power bidirectional
rlabel metal4 s 97688 2176 98008 117504 6 vdda1
port 645 nsew power bidirectional
rlabel metal4 s 66968 2176 67288 117504 6 vdda1
port 646 nsew power bidirectional
rlabel metal4 s 36248 2176 36568 117504 6 vdda1
port 647 nsew power bidirectional
rlabel metal4 s 5528 2176 5848 117504 6 vdda1
port 648 nsew power bidirectional
rlabel metal4 s 174488 2176 174808 117504 6 vssa1
port 649 nsew ground bidirectional
rlabel metal4 s 143768 2176 144088 117504 6 vssa1
port 650 nsew ground bidirectional
rlabel metal4 s 113048 2176 113368 117504 6 vssa1
port 651 nsew ground bidirectional
rlabel metal4 s 82328 2176 82648 117504 6 vssa1
port 652 nsew ground bidirectional
rlabel metal4 s 51608 2176 51928 117504 6 vssa1
port 653 nsew ground bidirectional
rlabel metal4 s 20888 2176 21208 117504 6 vssa1
port 654 nsew ground bidirectional
rlabel metal4 s 159788 2176 160108 117504 6 vdda2
port 655 nsew power bidirectional
rlabel metal4 s 129068 2176 129388 117504 6 vdda2
port 656 nsew power bidirectional
rlabel metal4 s 98348 2176 98668 117504 6 vdda2
port 657 nsew power bidirectional
rlabel metal4 s 67628 2176 67948 117504 6 vdda2
port 658 nsew power bidirectional
rlabel metal4 s 36908 2176 37228 117504 6 vdda2
port 659 nsew power bidirectional
rlabel metal4 s 6188 2176 6508 117504 6 vdda2
port 660 nsew power bidirectional
rlabel metal4 s 175148 2176 175468 117504 6 vssa2
port 661 nsew ground bidirectional
rlabel metal4 s 144428 2176 144748 117504 6 vssa2
port 662 nsew ground bidirectional
rlabel metal4 s 113708 2176 114028 117504 6 vssa2
port 663 nsew ground bidirectional
rlabel metal4 s 82988 2176 83308 117504 6 vssa2
port 664 nsew ground bidirectional
rlabel metal4 s 52268 2176 52588 117504 6 vssa2
port 665 nsew ground bidirectional
rlabel metal4 s 21548 2176 21868 117504 6 vssa2
port 666 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 180000 120000
string LEFview TRUE
string GDS_FILE /project/openlane/vco_adc_wrapper/runs/vco_adc_wrapper/results/magic/vco_adc_wrapper.gds
string GDS_END 17821656
string GDS_START 973706
<< end >>

